-------------------------------------------------------
--! @file exp_pkg.vhd
--! @brief Package for the exponential
--! @details 
--! @author Guido Baccelli
--! @version 1.
--! @date 23/08/2019
--! @bug NONE
--! @todo NONE
--! @copyright  GNU Public License [GPL-3.0].
-------------------------------------------------------
---------------- Copyright (c) notice -----------------------------------------
--
-- The VHDL code, the logic and concepts described in this file constitute
-- the intellectual property of the authors listed below, who are affiliated
-- to KTH(Kungliga Tekniska Högskolan), School of ICT, Kista.
-- Any unauthorised use, copy or distribution is strictly prohibited.
-- Any authorised use, copy or distribution should carry this copyright notice
-- unaltered.
-------------------------------------------------------------------------------
-- Title      : Exponential package
-- Project    : SiLago
-------------------------------------------------------------------------------
-- File       : exp_pkg.vhd
-- Author     : Guido Baccelli
-- Company    : KTH
-- Created    : 23/08/2019
-- Last update: 2020-03-15
-- Platform   : SiLago
-- Standard   : VHDL'08
-- Supervisor : Dimitrios Stathis
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Contact    : Dimitrios Stathis <stathis@kth.se>
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author                  Description
-- 23/08/2019  1.0      Guido Baccelli          Create
-- 2020-03-15  1.1      Dimitrios Stathis       Preparation for Git
-------------------------------------------------------------------------------

--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#
--                                                                         #
--This file is part of SiLago.                                             #
--                                                                         #
--    SiLago platform source code is distributed freely: you can           #
--    redistribute it and/or modify it under the terms of the GNU          #
--    General Public License as published by the Free Software Foundation, #
--    either version 3 of the License, or (at your option) any             #
--    later version.                                                       #
--                                                                         #
--    SiLago is distributed in the hope that it will be useful,            #
--    but WITHOUT ANY WARRANTY; without even the implied warranty of       #
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the        #
--    GNU General Public License for more details.                         #
--                                                                         #
--    You should have received a copy of the GNU General Public License    #
--    along with SiLago.  If not, see <https://www.gnu.org/licenses/>.     #
--                                                                         #
--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#

--! Standard ieee library
LIBRARY ieee;
--! Default working library
LIBRARY work;
--! Standard logic package
USE ieee.std_logic_1164.ALL;
--! Standard numeric package for signed and unsigned
USE ieee.numeric_std.ALL;

--! Package file with Exponential tail behavior model for Q4.11 fixed-point format (Generate with the help of matlab).

--! The only content is the 'exp_fp11' function that emulates behavior of Exponential tail calculation inside 'ann_unit'
PACKAGE exp_pkg IS

    FUNCTION exp_fp11(
        x : INTEGER
    ) RETURN INTEGER;

END PACKAGE exp_pkg;

--! @brief Contains body of function 'exp_fp11'
--! @details The function 'exp_fp11' (and the testbench) interpret input and output data words
--! as integer values instead of fixed-point values. This makes the model easier to describe.
--! The function describes the Exponential tail by assigning the corresponding output to each possible
--! input value representable on Q4.11.
PACKAGE BODY exp_pkg IS
    FUNCTION exp_fp11(
        x : INTEGER)
        RETURN INTEGER IS
        VARIABLE exp_f : INTEGER;
    BEGIN
        IF x =- 32768 THEN
            exp_f := 0;
        ELSIF x =- 32767 THEN
            exp_f := 0;
        ELSIF x =- 32766 THEN
            exp_f := 0;
        ELSIF x =- 32765 THEN
            exp_f := 0;
        ELSIF x =- 32764 THEN
            exp_f := 0;
        ELSIF x =- 32763 THEN
            exp_f := 0;
        ELSIF x =- 32762 THEN
            exp_f := 0;
        ELSIF x =- 32761 THEN
            exp_f := 0;
        ELSIF x =- 32760 THEN
            exp_f := 0;
        ELSIF x =- 32759 THEN
            exp_f := 0;
        ELSIF x =- 32758 THEN
            exp_f := 0;
        ELSIF x =- 32757 THEN
            exp_f := 0;
        ELSIF x =- 32756 THEN
            exp_f := 0;
        ELSIF x =- 32755 THEN
            exp_f := 0;
        ELSIF x =- 32754 THEN
            exp_f := 0;
        ELSIF x =- 32753 THEN
            exp_f := 0;
        ELSIF x =- 32752 THEN
            exp_f := 0;
        ELSIF x =- 32751 THEN
            exp_f := 0;
        ELSIF x =- 32750 THEN
            exp_f := 0;
        ELSIF x =- 32749 THEN
            exp_f := 0;
        ELSIF x =- 32748 THEN
            exp_f := 0;
        ELSIF x =- 32747 THEN
            exp_f := 0;
        ELSIF x =- 32746 THEN
            exp_f := 0;
        ELSIF x =- 32745 THEN
            exp_f := 0;
        ELSIF x =- 32744 THEN
            exp_f := 0;
        ELSIF x =- 32743 THEN
            exp_f := 0;
        ELSIF x =- 32742 THEN
            exp_f := 0;
        ELSIF x =- 32741 THEN
            exp_f := 0;
        ELSIF x =- 32740 THEN
            exp_f := 0;
        ELSIF x =- 32739 THEN
            exp_f := 0;
        ELSIF x =- 32738 THEN
            exp_f := 0;
        ELSIF x =- 32737 THEN
            exp_f := 0;
        ELSIF x =- 32736 THEN
            exp_f := 0;
        ELSIF x =- 32735 THEN
            exp_f := 0;
        ELSIF x =- 32734 THEN
            exp_f := 0;
        ELSIF x =- 32733 THEN
            exp_f := 0;
        ELSIF x =- 32732 THEN
            exp_f := 0;
        ELSIF x =- 32731 THEN
            exp_f := 0;
        ELSIF x =- 32730 THEN
            exp_f := 0;
        ELSIF x =- 32729 THEN
            exp_f := 0;
        ELSIF x =- 32728 THEN
            exp_f := 0;
        ELSIF x =- 32727 THEN
            exp_f := 0;
        ELSIF x =- 32726 THEN
            exp_f := 0;
        ELSIF x =- 32725 THEN
            exp_f := 0;
        ELSIF x =- 32724 THEN
            exp_f := 0;
        ELSIF x =- 32723 THEN
            exp_f := 0;
        ELSIF x =- 32722 THEN
            exp_f := 0;
        ELSIF x =- 32721 THEN
            exp_f := 0;
        ELSIF x =- 32720 THEN
            exp_f := 0;
        ELSIF x =- 32719 THEN
            exp_f := 0;
        ELSIF x =- 32718 THEN
            exp_f := 0;
        ELSIF x =- 32717 THEN
            exp_f := 0;
        ELSIF x =- 32716 THEN
            exp_f := 0;
        ELSIF x =- 32715 THEN
            exp_f := 0;
        ELSIF x =- 32714 THEN
            exp_f := 0;
        ELSIF x =- 32713 THEN
            exp_f := 0;
        ELSIF x =- 32712 THEN
            exp_f := 0;
        ELSIF x =- 32711 THEN
            exp_f := 0;
        ELSIF x =- 32710 THEN
            exp_f := 0;
        ELSIF x =- 32709 THEN
            exp_f := 0;
        ELSIF x =- 32708 THEN
            exp_f := 0;
        ELSIF x =- 32707 THEN
            exp_f := 0;
        ELSIF x =- 32706 THEN
            exp_f := 0;
        ELSIF x =- 32705 THEN
            exp_f := 0;
        ELSIF x =- 32704 THEN
            exp_f := 0;
        ELSIF x =- 32703 THEN
            exp_f := 0;
        ELSIF x =- 32702 THEN
            exp_f := 0;
        ELSIF x =- 32701 THEN
            exp_f := 0;
        ELSIF x =- 32700 THEN
            exp_f := 0;
        ELSIF x =- 32699 THEN
            exp_f := 0;
        ELSIF x =- 32698 THEN
            exp_f := 0;
        ELSIF x =- 32697 THEN
            exp_f := 0;
        ELSIF x =- 32696 THEN
            exp_f := 0;
        ELSIF x =- 32695 THEN
            exp_f := 0;
        ELSIF x =- 32694 THEN
            exp_f := 0;
        ELSIF x =- 32693 THEN
            exp_f := 0;
        ELSIF x =- 32692 THEN
            exp_f := 0;
        ELSIF x =- 32691 THEN
            exp_f := 0;
        ELSIF x =- 32690 THEN
            exp_f := 0;
        ELSIF x =- 32689 THEN
            exp_f := 0;
        ELSIF x =- 32688 THEN
            exp_f := 0;
        ELSIF x =- 32687 THEN
            exp_f := 0;
        ELSIF x =- 32686 THEN
            exp_f := 0;
        ELSIF x =- 32685 THEN
            exp_f := 0;
        ELSIF x =- 32684 THEN
            exp_f := 0;
        ELSIF x =- 32683 THEN
            exp_f := 0;
        ELSIF x =- 32682 THEN
            exp_f := 0;
        ELSIF x =- 32681 THEN
            exp_f := 0;
        ELSIF x =- 32680 THEN
            exp_f := 0;
        ELSIF x =- 32679 THEN
            exp_f := 0;
        ELSIF x =- 32678 THEN
            exp_f := 0;
        ELSIF x =- 32677 THEN
            exp_f := 0;
        ELSIF x =- 32676 THEN
            exp_f := 0;
        ELSIF x =- 32675 THEN
            exp_f := 0;
        ELSIF x =- 32674 THEN
            exp_f := 0;
        ELSIF x =- 32673 THEN
            exp_f := 0;
        ELSIF x =- 32672 THEN
            exp_f := 0;
        ELSIF x =- 32671 THEN
            exp_f := 0;
        ELSIF x =- 32670 THEN
            exp_f := 0;
        ELSIF x =- 32669 THEN
            exp_f := 0;
        ELSIF x =- 32668 THEN
            exp_f := 0;
        ELSIF x =- 32667 THEN
            exp_f := 0;
        ELSIF x =- 32666 THEN
            exp_f := 0;
        ELSIF x =- 32665 THEN
            exp_f := 0;
        ELSIF x =- 32664 THEN
            exp_f := 0;
        ELSIF x =- 32663 THEN
            exp_f := 0;
        ELSIF x =- 32662 THEN
            exp_f := 0;
        ELSIF x =- 32661 THEN
            exp_f := 0;
        ELSIF x =- 32660 THEN
            exp_f := 0;
        ELSIF x =- 32659 THEN
            exp_f := 0;
        ELSIF x =- 32658 THEN
            exp_f := 0;
        ELSIF x =- 32657 THEN
            exp_f := 0;
        ELSIF x =- 32656 THEN
            exp_f := 0;
        ELSIF x =- 32655 THEN
            exp_f := 0;
        ELSIF x =- 32654 THEN
            exp_f := 0;
        ELSIF x =- 32653 THEN
            exp_f := 0;
        ELSIF x =- 32652 THEN
            exp_f := 0;
        ELSIF x =- 32651 THEN
            exp_f := 0;
        ELSIF x =- 32650 THEN
            exp_f := 0;
        ELSIF x =- 32649 THEN
            exp_f := 0;
        ELSIF x =- 32648 THEN
            exp_f := 0;
        ELSIF x =- 32647 THEN
            exp_f := 0;
        ELSIF x =- 32646 THEN
            exp_f := 0;
        ELSIF x =- 32645 THEN
            exp_f := 0;
        ELSIF x =- 32644 THEN
            exp_f := 0;
        ELSIF x =- 32643 THEN
            exp_f := 0;
        ELSIF x =- 32642 THEN
            exp_f := 0;
        ELSIF x =- 32641 THEN
            exp_f := 0;
        ELSIF x =- 32640 THEN
            exp_f := 0;
        ELSIF x =- 32639 THEN
            exp_f := 0;
        ELSIF x =- 32638 THEN
            exp_f := 0;
        ELSIF x =- 32637 THEN
            exp_f := 0;
        ELSIF x =- 32636 THEN
            exp_f := 0;
        ELSIF x =- 32635 THEN
            exp_f := 0;
        ELSIF x =- 32634 THEN
            exp_f := 0;
        ELSIF x =- 32633 THEN
            exp_f := 0;
        ELSIF x =- 32632 THEN
            exp_f := 0;
        ELSIF x =- 32631 THEN
            exp_f := 0;
        ELSIF x =- 32630 THEN
            exp_f := 0;
        ELSIF x =- 32629 THEN
            exp_f := 0;
        ELSIF x =- 32628 THEN
            exp_f := 0;
        ELSIF x =- 32627 THEN
            exp_f := 0;
        ELSIF x =- 32626 THEN
            exp_f := 0;
        ELSIF x =- 32625 THEN
            exp_f := 0;
        ELSIF x =- 32624 THEN
            exp_f := 0;
        ELSIF x =- 32623 THEN
            exp_f := 0;
        ELSIF x =- 32622 THEN
            exp_f := 0;
        ELSIF x =- 32621 THEN
            exp_f := 0;
        ELSIF x =- 32620 THEN
            exp_f := 0;
        ELSIF x =- 32619 THEN
            exp_f := 0;
        ELSIF x =- 32618 THEN
            exp_f := 0;
        ELSIF x =- 32617 THEN
            exp_f := 0;
        ELSIF x =- 32616 THEN
            exp_f := 0;
        ELSIF x =- 32615 THEN
            exp_f := 0;
        ELSIF x =- 32614 THEN
            exp_f := 0;
        ELSIF x =- 32613 THEN
            exp_f := 0;
        ELSIF x =- 32612 THEN
            exp_f := 0;
        ELSIF x =- 32611 THEN
            exp_f := 0;
        ELSIF x =- 32610 THEN
            exp_f := 0;
        ELSIF x =- 32609 THEN
            exp_f := 0;
        ELSIF x =- 32608 THEN
            exp_f := 0;
        ELSIF x =- 32607 THEN
            exp_f := 0;
        ELSIF x =- 32606 THEN
            exp_f := 0;
        ELSIF x =- 32605 THEN
            exp_f := 0;
        ELSIF x =- 32604 THEN
            exp_f := 0;
        ELSIF x =- 32603 THEN
            exp_f := 0;
        ELSIF x =- 32602 THEN
            exp_f := 0;
        ELSIF x =- 32601 THEN
            exp_f := 0;
        ELSIF x =- 32600 THEN
            exp_f := 0;
        ELSIF x =- 32599 THEN
            exp_f := 0;
        ELSIF x =- 32598 THEN
            exp_f := 0;
        ELSIF x =- 32597 THEN
            exp_f := 0;
        ELSIF x =- 32596 THEN
            exp_f := 0;
        ELSIF x =- 32595 THEN
            exp_f := 0;
        ELSIF x =- 32594 THEN
            exp_f := 0;
        ELSIF x =- 32593 THEN
            exp_f := 0;
        ELSIF x =- 32592 THEN
            exp_f := 0;
        ELSIF x =- 32591 THEN
            exp_f := 0;
        ELSIF x =- 32590 THEN
            exp_f := 0;
        ELSIF x =- 32589 THEN
            exp_f := 0;
        ELSIF x =- 32588 THEN
            exp_f := 0;
        ELSIF x =- 32587 THEN
            exp_f := 0;
        ELSIF x =- 32586 THEN
            exp_f := 0;
        ELSIF x =- 32585 THEN
            exp_f := 0;
        ELSIF x =- 32584 THEN
            exp_f := 0;
        ELSIF x =- 32583 THEN
            exp_f := 0;
        ELSIF x =- 32582 THEN
            exp_f := 0;
        ELSIF x =- 32581 THEN
            exp_f := 0;
        ELSIF x =- 32580 THEN
            exp_f := 0;
        ELSIF x =- 32579 THEN
            exp_f := 0;
        ELSIF x =- 32578 THEN
            exp_f := 0;
        ELSIF x =- 32577 THEN
            exp_f := 0;
        ELSIF x =- 32576 THEN
            exp_f := 0;
        ELSIF x =- 32575 THEN
            exp_f := 0;
        ELSIF x =- 32574 THEN
            exp_f := 0;
        ELSIF x =- 32573 THEN
            exp_f := 0;
        ELSIF x =- 32572 THEN
            exp_f := 0;
        ELSIF x =- 32571 THEN
            exp_f := 0;
        ELSIF x =- 32570 THEN
            exp_f := 0;
        ELSIF x =- 32569 THEN
            exp_f := 0;
        ELSIF x =- 32568 THEN
            exp_f := 0;
        ELSIF x =- 32567 THEN
            exp_f := 0;
        ELSIF x =- 32566 THEN
            exp_f := 0;
        ELSIF x =- 32565 THEN
            exp_f := 0;
        ELSIF x =- 32564 THEN
            exp_f := 0;
        ELSIF x =- 32563 THEN
            exp_f := 0;
        ELSIF x =- 32562 THEN
            exp_f := 0;
        ELSIF x =- 32561 THEN
            exp_f := 0;
        ELSIF x =- 32560 THEN
            exp_f := 0;
        ELSIF x =- 32559 THEN
            exp_f := 0;
        ELSIF x =- 32558 THEN
            exp_f := 0;
        ELSIF x =- 32557 THEN
            exp_f := 0;
        ELSIF x =- 32556 THEN
            exp_f := 0;
        ELSIF x =- 32555 THEN
            exp_f := 0;
        ELSIF x =- 32554 THEN
            exp_f := 0;
        ELSIF x =- 32553 THEN
            exp_f := 0;
        ELSIF x =- 32552 THEN
            exp_f := 0;
        ELSIF x =- 32551 THEN
            exp_f := 0;
        ELSIF x =- 32550 THEN
            exp_f := 0;
        ELSIF x =- 32549 THEN
            exp_f := 0;
        ELSIF x =- 32548 THEN
            exp_f := 0;
        ELSIF x =- 32547 THEN
            exp_f := 0;
        ELSIF x =- 32546 THEN
            exp_f := 0;
        ELSIF x =- 32545 THEN
            exp_f := 0;
        ELSIF x =- 32544 THEN
            exp_f := 0;
        ELSIF x =- 32543 THEN
            exp_f := 0;
        ELSIF x =- 32542 THEN
            exp_f := 0;
        ELSIF x =- 32541 THEN
            exp_f := 0;
        ELSIF x =- 32540 THEN
            exp_f := 0;
        ELSIF x =- 32539 THEN
            exp_f := 0;
        ELSIF x =- 32538 THEN
            exp_f := 0;
        ELSIF x =- 32537 THEN
            exp_f := 0;
        ELSIF x =- 32536 THEN
            exp_f := 0;
        ELSIF x =- 32535 THEN
            exp_f := 0;
        ELSIF x =- 32534 THEN
            exp_f := 0;
        ELSIF x =- 32533 THEN
            exp_f := 0;
        ELSIF x =- 32532 THEN
            exp_f := 0;
        ELSIF x =- 32531 THEN
            exp_f := 0;
        ELSIF x =- 32530 THEN
            exp_f := 0;
        ELSIF x =- 32529 THEN
            exp_f := 0;
        ELSIF x =- 32528 THEN
            exp_f := 0;
        ELSIF x =- 32527 THEN
            exp_f := 0;
        ELSIF x =- 32526 THEN
            exp_f := 0;
        ELSIF x =- 32525 THEN
            exp_f := 0;
        ELSIF x =- 32524 THEN
            exp_f := 0;
        ELSIF x =- 32523 THEN
            exp_f := 0;
        ELSIF x =- 32522 THEN
            exp_f := 0;
        ELSIF x =- 32521 THEN
            exp_f := 0;
        ELSIF x =- 32520 THEN
            exp_f := 0;
        ELSIF x =- 32519 THEN
            exp_f := 0;
        ELSIF x =- 32518 THEN
            exp_f := 0;
        ELSIF x =- 32517 THEN
            exp_f := 0;
        ELSIF x =- 32516 THEN
            exp_f := 0;
        ELSIF x =- 32515 THEN
            exp_f := 0;
        ELSIF x =- 32514 THEN
            exp_f := 0;
        ELSIF x =- 32513 THEN
            exp_f := 0;
        ELSIF x =- 32512 THEN
            exp_f := 0;
        ELSIF x =- 32511 THEN
            exp_f := 0;
        ELSIF x =- 32510 THEN
            exp_f := 0;
        ELSIF x =- 32509 THEN
            exp_f := 0;
        ELSIF x =- 32508 THEN
            exp_f := 0;
        ELSIF x =- 32507 THEN
            exp_f := 0;
        ELSIF x =- 32506 THEN
            exp_f := 0;
        ELSIF x =- 32505 THEN
            exp_f := 0;
        ELSIF x =- 32504 THEN
            exp_f := 0;
        ELSIF x =- 32503 THEN
            exp_f := 0;
        ELSIF x =- 32502 THEN
            exp_f := 0;
        ELSIF x =- 32501 THEN
            exp_f := 0;
        ELSIF x =- 32500 THEN
            exp_f := 0;
        ELSIF x =- 32499 THEN
            exp_f := 0;
        ELSIF x =- 32498 THEN
            exp_f := 0;
        ELSIF x =- 32497 THEN
            exp_f := 0;
        ELSIF x =- 32496 THEN
            exp_f := 0;
        ELSIF x =- 32495 THEN
            exp_f := 0;
        ELSIF x =- 32494 THEN
            exp_f := 0;
        ELSIF x =- 32493 THEN
            exp_f := 0;
        ELSIF x =- 32492 THEN
            exp_f := 0;
        ELSIF x =- 32491 THEN
            exp_f := 0;
        ELSIF x =- 32490 THEN
            exp_f := 0;
        ELSIF x =- 32489 THEN
            exp_f := 0;
        ELSIF x =- 32488 THEN
            exp_f := 0;
        ELSIF x =- 32487 THEN
            exp_f := 0;
        ELSIF x =- 32486 THEN
            exp_f := 0;
        ELSIF x =- 32485 THEN
            exp_f := 0;
        ELSIF x =- 32484 THEN
            exp_f := 0;
        ELSIF x =- 32483 THEN
            exp_f := 0;
        ELSIF x =- 32482 THEN
            exp_f := 0;
        ELSIF x =- 32481 THEN
            exp_f := 0;
        ELSIF x =- 32480 THEN
            exp_f := 0;
        ELSIF x =- 32479 THEN
            exp_f := 0;
        ELSIF x =- 32478 THEN
            exp_f := 0;
        ELSIF x =- 32477 THEN
            exp_f := 0;
        ELSIF x =- 32476 THEN
            exp_f := 0;
        ELSIF x =- 32475 THEN
            exp_f := 0;
        ELSIF x =- 32474 THEN
            exp_f := 0;
        ELSIF x =- 32473 THEN
            exp_f := 0;
        ELSIF x =- 32472 THEN
            exp_f := 0;
        ELSIF x =- 32471 THEN
            exp_f := 0;
        ELSIF x =- 32470 THEN
            exp_f := 0;
        ELSIF x =- 32469 THEN
            exp_f := 0;
        ELSIF x =- 32468 THEN
            exp_f := 0;
        ELSIF x =- 32467 THEN
            exp_f := 0;
        ELSIF x =- 32466 THEN
            exp_f := 0;
        ELSIF x =- 32465 THEN
            exp_f := 0;
        ELSIF x =- 32464 THEN
            exp_f := 0;
        ELSIF x =- 32463 THEN
            exp_f := 0;
        ELSIF x =- 32462 THEN
            exp_f := 0;
        ELSIF x =- 32461 THEN
            exp_f := 0;
        ELSIF x =- 32460 THEN
            exp_f := 0;
        ELSIF x =- 32459 THEN
            exp_f := 0;
        ELSIF x =- 32458 THEN
            exp_f := 0;
        ELSIF x =- 32457 THEN
            exp_f := 0;
        ELSIF x =- 32456 THEN
            exp_f := 0;
        ELSIF x =- 32455 THEN
            exp_f := 0;
        ELSIF x =- 32454 THEN
            exp_f := 0;
        ELSIF x =- 32453 THEN
            exp_f := 0;
        ELSIF x =- 32452 THEN
            exp_f := 0;
        ELSIF x =- 32451 THEN
            exp_f := 0;
        ELSIF x =- 32450 THEN
            exp_f := 0;
        ELSIF x =- 32449 THEN
            exp_f := 0;
        ELSIF x =- 32448 THEN
            exp_f := 0;
        ELSIF x =- 32447 THEN
            exp_f := 0;
        ELSIF x =- 32446 THEN
            exp_f := 0;
        ELSIF x =- 32445 THEN
            exp_f := 0;
        ELSIF x =- 32444 THEN
            exp_f := 0;
        ELSIF x =- 32443 THEN
            exp_f := 0;
        ELSIF x =- 32442 THEN
            exp_f := 0;
        ELSIF x =- 32441 THEN
            exp_f := 0;
        ELSIF x =- 32440 THEN
            exp_f := 0;
        ELSIF x =- 32439 THEN
            exp_f := 0;
        ELSIF x =- 32438 THEN
            exp_f := 0;
        ELSIF x =- 32437 THEN
            exp_f := 0;
        ELSIF x =- 32436 THEN
            exp_f := 0;
        ELSIF x =- 32435 THEN
            exp_f := 0;
        ELSIF x =- 32434 THEN
            exp_f := 0;
        ELSIF x =- 32433 THEN
            exp_f := 0;
        ELSIF x =- 32432 THEN
            exp_f := 0;
        ELSIF x =- 32431 THEN
            exp_f := 0;
        ELSIF x =- 32430 THEN
            exp_f := 0;
        ELSIF x =- 32429 THEN
            exp_f := 0;
        ELSIF x =- 32428 THEN
            exp_f := 0;
        ELSIF x =- 32427 THEN
            exp_f := 0;
        ELSIF x =- 32426 THEN
            exp_f := 0;
        ELSIF x =- 32425 THEN
            exp_f := 0;
        ELSIF x =- 32424 THEN
            exp_f := 0;
        ELSIF x =- 32423 THEN
            exp_f := 0;
        ELSIF x =- 32422 THEN
            exp_f := 0;
        ELSIF x =- 32421 THEN
            exp_f := 0;
        ELSIF x =- 32420 THEN
            exp_f := 0;
        ELSIF x =- 32419 THEN
            exp_f := 0;
        ELSIF x =- 32418 THEN
            exp_f := 0;
        ELSIF x =- 32417 THEN
            exp_f := 0;
        ELSIF x =- 32416 THEN
            exp_f := 0;
        ELSIF x =- 32415 THEN
            exp_f := 0;
        ELSIF x =- 32414 THEN
            exp_f := 0;
        ELSIF x =- 32413 THEN
            exp_f := 0;
        ELSIF x =- 32412 THEN
            exp_f := 0;
        ELSIF x =- 32411 THEN
            exp_f := 0;
        ELSIF x =- 32410 THEN
            exp_f := 0;
        ELSIF x =- 32409 THEN
            exp_f := 0;
        ELSIF x =- 32408 THEN
            exp_f := 0;
        ELSIF x =- 32407 THEN
            exp_f := 0;
        ELSIF x =- 32406 THEN
            exp_f := 0;
        ELSIF x =- 32405 THEN
            exp_f := 0;
        ELSIF x =- 32404 THEN
            exp_f := 0;
        ELSIF x =- 32403 THEN
            exp_f := 0;
        ELSIF x =- 32402 THEN
            exp_f := 0;
        ELSIF x =- 32401 THEN
            exp_f := 0;
        ELSIF x =- 32400 THEN
            exp_f := 0;
        ELSIF x =- 32399 THEN
            exp_f := 0;
        ELSIF x =- 32398 THEN
            exp_f := 0;
        ELSIF x =- 32397 THEN
            exp_f := 0;
        ELSIF x =- 32396 THEN
            exp_f := 0;
        ELSIF x =- 32395 THEN
            exp_f := 0;
        ELSIF x =- 32394 THEN
            exp_f := 0;
        ELSIF x =- 32393 THEN
            exp_f := 0;
        ELSIF x =- 32392 THEN
            exp_f := 0;
        ELSIF x =- 32391 THEN
            exp_f := 0;
        ELSIF x =- 32390 THEN
            exp_f := 0;
        ELSIF x =- 32389 THEN
            exp_f := 0;
        ELSIF x =- 32388 THEN
            exp_f := 0;
        ELSIF x =- 32387 THEN
            exp_f := 0;
        ELSIF x =- 32386 THEN
            exp_f := 0;
        ELSIF x =- 32385 THEN
            exp_f := 0;
        ELSIF x =- 32384 THEN
            exp_f := 0;
        ELSIF x =- 32383 THEN
            exp_f := 0;
        ELSIF x =- 32382 THEN
            exp_f := 0;
        ELSIF x =- 32381 THEN
            exp_f := 0;
        ELSIF x =- 32380 THEN
            exp_f := 0;
        ELSIF x =- 32379 THEN
            exp_f := 0;
        ELSIF x =- 32378 THEN
            exp_f := 0;
        ELSIF x =- 32377 THEN
            exp_f := 0;
        ELSIF x =- 32376 THEN
            exp_f := 0;
        ELSIF x =- 32375 THEN
            exp_f := 0;
        ELSIF x =- 32374 THEN
            exp_f := 0;
        ELSIF x =- 32373 THEN
            exp_f := 0;
        ELSIF x =- 32372 THEN
            exp_f := 0;
        ELSIF x =- 32371 THEN
            exp_f := 0;
        ELSIF x =- 32370 THEN
            exp_f := 0;
        ELSIF x =- 32369 THEN
            exp_f := 0;
        ELSIF x =- 32368 THEN
            exp_f := 0;
        ELSIF x =- 32367 THEN
            exp_f := 0;
        ELSIF x =- 32366 THEN
            exp_f := 0;
        ELSIF x =- 32365 THEN
            exp_f := 0;
        ELSIF x =- 32364 THEN
            exp_f := 0;
        ELSIF x =- 32363 THEN
            exp_f := 0;
        ELSIF x =- 32362 THEN
            exp_f := 0;
        ELSIF x =- 32361 THEN
            exp_f := 0;
        ELSIF x =- 32360 THEN
            exp_f := 0;
        ELSIF x =- 32359 THEN
            exp_f := 0;
        ELSIF x =- 32358 THEN
            exp_f := 0;
        ELSIF x =- 32357 THEN
            exp_f := 0;
        ELSIF x =- 32356 THEN
            exp_f := 0;
        ELSIF x =- 32355 THEN
            exp_f := 0;
        ELSIF x =- 32354 THEN
            exp_f := 0;
        ELSIF x =- 32353 THEN
            exp_f := 0;
        ELSIF x =- 32352 THEN
            exp_f := 0;
        ELSIF x =- 32351 THEN
            exp_f := 0;
        ELSIF x =- 32350 THEN
            exp_f := 0;
        ELSIF x =- 32349 THEN
            exp_f := 0;
        ELSIF x =- 32348 THEN
            exp_f := 0;
        ELSIF x =- 32347 THEN
            exp_f := 0;
        ELSIF x =- 32346 THEN
            exp_f := 0;
        ELSIF x =- 32345 THEN
            exp_f := 0;
        ELSIF x =- 32344 THEN
            exp_f := 0;
        ELSIF x =- 32343 THEN
            exp_f := 0;
        ELSIF x =- 32342 THEN
            exp_f := 0;
        ELSIF x =- 32341 THEN
            exp_f := 0;
        ELSIF x =- 32340 THEN
            exp_f := 0;
        ELSIF x =- 32339 THEN
            exp_f := 0;
        ELSIF x =- 32338 THEN
            exp_f := 0;
        ELSIF x =- 32337 THEN
            exp_f := 0;
        ELSIF x =- 32336 THEN
            exp_f := 0;
        ELSIF x =- 32335 THEN
            exp_f := 0;
        ELSIF x =- 32334 THEN
            exp_f := 0;
        ELSIF x =- 32333 THEN
            exp_f := 0;
        ELSIF x =- 32332 THEN
            exp_f := 0;
        ELSIF x =- 32331 THEN
            exp_f := 0;
        ELSIF x =- 32330 THEN
            exp_f := 0;
        ELSIF x =- 32329 THEN
            exp_f := 0;
        ELSIF x =- 32328 THEN
            exp_f := 0;
        ELSIF x =- 32327 THEN
            exp_f := 0;
        ELSIF x =- 32326 THEN
            exp_f := 0;
        ELSIF x =- 32325 THEN
            exp_f := 0;
        ELSIF x =- 32324 THEN
            exp_f := 0;
        ELSIF x =- 32323 THEN
            exp_f := 0;
        ELSIF x =- 32322 THEN
            exp_f := 0;
        ELSIF x =- 32321 THEN
            exp_f := 0;
        ELSIF x =- 32320 THEN
            exp_f := 0;
        ELSIF x =- 32319 THEN
            exp_f := 0;
        ELSIF x =- 32318 THEN
            exp_f := 0;
        ELSIF x =- 32317 THEN
            exp_f := 0;
        ELSIF x =- 32316 THEN
            exp_f := 0;
        ELSIF x =- 32315 THEN
            exp_f := 0;
        ELSIF x =- 32314 THEN
            exp_f := 0;
        ELSIF x =- 32313 THEN
            exp_f := 0;
        ELSIF x =- 32312 THEN
            exp_f := 0;
        ELSIF x =- 32311 THEN
            exp_f := 0;
        ELSIF x =- 32310 THEN
            exp_f := 0;
        ELSIF x =- 32309 THEN
            exp_f := 0;
        ELSIF x =- 32308 THEN
            exp_f := 0;
        ELSIF x =- 32307 THEN
            exp_f := 0;
        ELSIF x =- 32306 THEN
            exp_f := 0;
        ELSIF x =- 32305 THEN
            exp_f := 0;
        ELSIF x =- 32304 THEN
            exp_f := 0;
        ELSIF x =- 32303 THEN
            exp_f := 0;
        ELSIF x =- 32302 THEN
            exp_f := 0;
        ELSIF x =- 32301 THEN
            exp_f := 0;
        ELSIF x =- 32300 THEN
            exp_f := 0;
        ELSIF x =- 32299 THEN
            exp_f := 0;
        ELSIF x =- 32298 THEN
            exp_f := 0;
        ELSIF x =- 32297 THEN
            exp_f := 0;
        ELSIF x =- 32296 THEN
            exp_f := 0;
        ELSIF x =- 32295 THEN
            exp_f := 0;
        ELSIF x =- 32294 THEN
            exp_f := 0;
        ELSIF x =- 32293 THEN
            exp_f := 0;
        ELSIF x =- 32292 THEN
            exp_f := 0;
        ELSIF x =- 32291 THEN
            exp_f := 0;
        ELSIF x =- 32290 THEN
            exp_f := 0;
        ELSIF x =- 32289 THEN
            exp_f := 0;
        ELSIF x =- 32288 THEN
            exp_f := 0;
        ELSIF x =- 32287 THEN
            exp_f := 0;
        ELSIF x =- 32286 THEN
            exp_f := 0;
        ELSIF x =- 32285 THEN
            exp_f := 0;
        ELSIF x =- 32284 THEN
            exp_f := 0;
        ELSIF x =- 32283 THEN
            exp_f := 0;
        ELSIF x =- 32282 THEN
            exp_f := 0;
        ELSIF x =- 32281 THEN
            exp_f := 0;
        ELSIF x =- 32280 THEN
            exp_f := 0;
        ELSIF x =- 32279 THEN
            exp_f := 0;
        ELSIF x =- 32278 THEN
            exp_f := 0;
        ELSIF x =- 32277 THEN
            exp_f := 0;
        ELSIF x =- 32276 THEN
            exp_f := 0;
        ELSIF x =- 32275 THEN
            exp_f := 0;
        ELSIF x =- 32274 THEN
            exp_f := 0;
        ELSIF x =- 32273 THEN
            exp_f := 0;
        ELSIF x =- 32272 THEN
            exp_f := 0;
        ELSIF x =- 32271 THEN
            exp_f := 0;
        ELSIF x =- 32270 THEN
            exp_f := 0;
        ELSIF x =- 32269 THEN
            exp_f := 0;
        ELSIF x =- 32268 THEN
            exp_f := 0;
        ELSIF x =- 32267 THEN
            exp_f := 0;
        ELSIF x =- 32266 THEN
            exp_f := 0;
        ELSIF x =- 32265 THEN
            exp_f := 0;
        ELSIF x =- 32264 THEN
            exp_f := 0;
        ELSIF x =- 32263 THEN
            exp_f := 0;
        ELSIF x =- 32262 THEN
            exp_f := 0;
        ELSIF x =- 32261 THEN
            exp_f := 0;
        ELSIF x =- 32260 THEN
            exp_f := 0;
        ELSIF x =- 32259 THEN
            exp_f := 0;
        ELSIF x =- 32258 THEN
            exp_f := 0;
        ELSIF x =- 32257 THEN
            exp_f := 0;
        ELSIF x =- 32256 THEN
            exp_f := 0;
        ELSIF x =- 32255 THEN
            exp_f := 0;
        ELSIF x =- 32254 THEN
            exp_f := 0;
        ELSIF x =- 32253 THEN
            exp_f := 0;
        ELSIF x =- 32252 THEN
            exp_f := 0;
        ELSIF x =- 32251 THEN
            exp_f := 0;
        ELSIF x =- 32250 THEN
            exp_f := 0;
        ELSIF x =- 32249 THEN
            exp_f := 0;
        ELSIF x =- 32248 THEN
            exp_f := 0;
        ELSIF x =- 32247 THEN
            exp_f := 0;
        ELSIF x =- 32246 THEN
            exp_f := 0;
        ELSIF x =- 32245 THEN
            exp_f := 0;
        ELSIF x =- 32244 THEN
            exp_f := 0;
        ELSIF x =- 32243 THEN
            exp_f := 0;
        ELSIF x =- 32242 THEN
            exp_f := 0;
        ELSIF x =- 32241 THEN
            exp_f := 0;
        ELSIF x =- 32240 THEN
            exp_f := 0;
        ELSIF x =- 32239 THEN
            exp_f := 0;
        ELSIF x =- 32238 THEN
            exp_f := 0;
        ELSIF x =- 32237 THEN
            exp_f := 0;
        ELSIF x =- 32236 THEN
            exp_f := 0;
        ELSIF x =- 32235 THEN
            exp_f := 0;
        ELSIF x =- 32234 THEN
            exp_f := 0;
        ELSIF x =- 32233 THEN
            exp_f := 0;
        ELSIF x =- 32232 THEN
            exp_f := 0;
        ELSIF x =- 32231 THEN
            exp_f := 0;
        ELSIF x =- 32230 THEN
            exp_f := 0;
        ELSIF x =- 32229 THEN
            exp_f := 0;
        ELSIF x =- 32228 THEN
            exp_f := 0;
        ELSIF x =- 32227 THEN
            exp_f := 0;
        ELSIF x =- 32226 THEN
            exp_f := 0;
        ELSIF x =- 32225 THEN
            exp_f := 0;
        ELSIF x =- 32224 THEN
            exp_f := 0;
        ELSIF x =- 32223 THEN
            exp_f := 0;
        ELSIF x =- 32222 THEN
            exp_f := 0;
        ELSIF x =- 32221 THEN
            exp_f := 0;
        ELSIF x =- 32220 THEN
            exp_f := 0;
        ELSIF x =- 32219 THEN
            exp_f := 0;
        ELSIF x =- 32218 THEN
            exp_f := 0;
        ELSIF x =- 32217 THEN
            exp_f := 0;
        ELSIF x =- 32216 THEN
            exp_f := 0;
        ELSIF x =- 32215 THEN
            exp_f := 0;
        ELSIF x =- 32214 THEN
            exp_f := 0;
        ELSIF x =- 32213 THEN
            exp_f := 0;
        ELSIF x =- 32212 THEN
            exp_f := 0;
        ELSIF x =- 32211 THEN
            exp_f := 0;
        ELSIF x =- 32210 THEN
            exp_f := 0;
        ELSIF x =- 32209 THEN
            exp_f := 0;
        ELSIF x =- 32208 THEN
            exp_f := 0;
        ELSIF x =- 32207 THEN
            exp_f := 0;
        ELSIF x =- 32206 THEN
            exp_f := 0;
        ELSIF x =- 32205 THEN
            exp_f := 0;
        ELSIF x =- 32204 THEN
            exp_f := 0;
        ELSIF x =- 32203 THEN
            exp_f := 0;
        ELSIF x =- 32202 THEN
            exp_f := 0;
        ELSIF x =- 32201 THEN
            exp_f := 0;
        ELSIF x =- 32200 THEN
            exp_f := 0;
        ELSIF x =- 32199 THEN
            exp_f := 0;
        ELSIF x =- 32198 THEN
            exp_f := 0;
        ELSIF x =- 32197 THEN
            exp_f := 0;
        ELSIF x =- 32196 THEN
            exp_f := 0;
        ELSIF x =- 32195 THEN
            exp_f := 0;
        ELSIF x =- 32194 THEN
            exp_f := 0;
        ELSIF x =- 32193 THEN
            exp_f := 0;
        ELSIF x =- 32192 THEN
            exp_f := 0;
        ELSIF x =- 32191 THEN
            exp_f := 0;
        ELSIF x =- 32190 THEN
            exp_f := 0;
        ELSIF x =- 32189 THEN
            exp_f := 0;
        ELSIF x =- 32188 THEN
            exp_f := 0;
        ELSIF x =- 32187 THEN
            exp_f := 0;
        ELSIF x =- 32186 THEN
            exp_f := 0;
        ELSIF x =- 32185 THEN
            exp_f := 0;
        ELSIF x =- 32184 THEN
            exp_f := 0;
        ELSIF x =- 32183 THEN
            exp_f := 0;
        ELSIF x =- 32182 THEN
            exp_f := 0;
        ELSIF x =- 32181 THEN
            exp_f := 0;
        ELSIF x =- 32180 THEN
            exp_f := 0;
        ELSIF x =- 32179 THEN
            exp_f := 0;
        ELSIF x =- 32178 THEN
            exp_f := 0;
        ELSIF x =- 32177 THEN
            exp_f := 0;
        ELSIF x =- 32176 THEN
            exp_f := 0;
        ELSIF x =- 32175 THEN
            exp_f := 0;
        ELSIF x =- 32174 THEN
            exp_f := 0;
        ELSIF x =- 32173 THEN
            exp_f := 0;
        ELSIF x =- 32172 THEN
            exp_f := 0;
        ELSIF x =- 32171 THEN
            exp_f := 0;
        ELSIF x =- 32170 THEN
            exp_f := 0;
        ELSIF x =- 32169 THEN
            exp_f := 0;
        ELSIF x =- 32168 THEN
            exp_f := 0;
        ELSIF x =- 32167 THEN
            exp_f := 0;
        ELSIF x =- 32166 THEN
            exp_f := 0;
        ELSIF x =- 32165 THEN
            exp_f := 0;
        ELSIF x =- 32164 THEN
            exp_f := 0;
        ELSIF x =- 32163 THEN
            exp_f := 0;
        ELSIF x =- 32162 THEN
            exp_f := 0;
        ELSIF x =- 32161 THEN
            exp_f := 0;
        ELSIF x =- 32160 THEN
            exp_f := 0;
        ELSIF x =- 32159 THEN
            exp_f := 0;
        ELSIF x =- 32158 THEN
            exp_f := 0;
        ELSIF x =- 32157 THEN
            exp_f := 0;
        ELSIF x =- 32156 THEN
            exp_f := 0;
        ELSIF x =- 32155 THEN
            exp_f := 0;
        ELSIF x =- 32154 THEN
            exp_f := 0;
        ELSIF x =- 32153 THEN
            exp_f := 0;
        ELSIF x =- 32152 THEN
            exp_f := 0;
        ELSIF x =- 32151 THEN
            exp_f := 0;
        ELSIF x =- 32150 THEN
            exp_f := 0;
        ELSIF x =- 32149 THEN
            exp_f := 0;
        ELSIF x =- 32148 THEN
            exp_f := 0;
        ELSIF x =- 32147 THEN
            exp_f := 0;
        ELSIF x =- 32146 THEN
            exp_f := 0;
        ELSIF x =- 32145 THEN
            exp_f := 0;
        ELSIF x =- 32144 THEN
            exp_f := 0;
        ELSIF x =- 32143 THEN
            exp_f := 0;
        ELSIF x =- 32142 THEN
            exp_f := 0;
        ELSIF x =- 32141 THEN
            exp_f := 0;
        ELSIF x =- 32140 THEN
            exp_f := 0;
        ELSIF x =- 32139 THEN
            exp_f := 0;
        ELSIF x =- 32138 THEN
            exp_f := 0;
        ELSIF x =- 32137 THEN
            exp_f := 0;
        ELSIF x =- 32136 THEN
            exp_f := 0;
        ELSIF x =- 32135 THEN
            exp_f := 0;
        ELSIF x =- 32134 THEN
            exp_f := 0;
        ELSIF x =- 32133 THEN
            exp_f := 0;
        ELSIF x =- 32132 THEN
            exp_f := 0;
        ELSIF x =- 32131 THEN
            exp_f := 0;
        ELSIF x =- 32130 THEN
            exp_f := 0;
        ELSIF x =- 32129 THEN
            exp_f := 0;
        ELSIF x =- 32128 THEN
            exp_f := 0;
        ELSIF x =- 32127 THEN
            exp_f := 0;
        ELSIF x =- 32126 THEN
            exp_f := 0;
        ELSIF x =- 32125 THEN
            exp_f := 0;
        ELSIF x =- 32124 THEN
            exp_f := 0;
        ELSIF x =- 32123 THEN
            exp_f := 0;
        ELSIF x =- 32122 THEN
            exp_f := 0;
        ELSIF x =- 32121 THEN
            exp_f := 0;
        ELSIF x =- 32120 THEN
            exp_f := 0;
        ELSIF x =- 32119 THEN
            exp_f := 0;
        ELSIF x =- 32118 THEN
            exp_f := 0;
        ELSIF x =- 32117 THEN
            exp_f := 0;
        ELSIF x =- 32116 THEN
            exp_f := 0;
        ELSIF x =- 32115 THEN
            exp_f := 0;
        ELSIF x =- 32114 THEN
            exp_f := 0;
        ELSIF x =- 32113 THEN
            exp_f := 0;
        ELSIF x =- 32112 THEN
            exp_f := 0;
        ELSIF x =- 32111 THEN
            exp_f := 0;
        ELSIF x =- 32110 THEN
            exp_f := 0;
        ELSIF x =- 32109 THEN
            exp_f := 0;
        ELSIF x =- 32108 THEN
            exp_f := 0;
        ELSIF x =- 32107 THEN
            exp_f := 0;
        ELSIF x =- 32106 THEN
            exp_f := 0;
        ELSIF x =- 32105 THEN
            exp_f := 0;
        ELSIF x =- 32104 THEN
            exp_f := 0;
        ELSIF x =- 32103 THEN
            exp_f := 0;
        ELSIF x =- 32102 THEN
            exp_f := 0;
        ELSIF x =- 32101 THEN
            exp_f := 0;
        ELSIF x =- 32100 THEN
            exp_f := 0;
        ELSIF x =- 32099 THEN
            exp_f := 0;
        ELSIF x =- 32098 THEN
            exp_f := 0;
        ELSIF x =- 32097 THEN
            exp_f := 0;
        ELSIF x =- 32096 THEN
            exp_f := 0;
        ELSIF x =- 32095 THEN
            exp_f := 0;
        ELSIF x =- 32094 THEN
            exp_f := 0;
        ELSIF x =- 32093 THEN
            exp_f := 0;
        ELSIF x =- 32092 THEN
            exp_f := 0;
        ELSIF x =- 32091 THEN
            exp_f := 0;
        ELSIF x =- 32090 THEN
            exp_f := 0;
        ELSIF x =- 32089 THEN
            exp_f := 0;
        ELSIF x =- 32088 THEN
            exp_f := 0;
        ELSIF x =- 32087 THEN
            exp_f := 0;
        ELSIF x =- 32086 THEN
            exp_f := 0;
        ELSIF x =- 32085 THEN
            exp_f := 0;
        ELSIF x =- 32084 THEN
            exp_f := 0;
        ELSIF x =- 32083 THEN
            exp_f := 0;
        ELSIF x =- 32082 THEN
            exp_f := 0;
        ELSIF x =- 32081 THEN
            exp_f := 0;
        ELSIF x =- 32080 THEN
            exp_f := 0;
        ELSIF x =- 32079 THEN
            exp_f := 0;
        ELSIF x =- 32078 THEN
            exp_f := 0;
        ELSIF x =- 32077 THEN
            exp_f := 0;
        ELSIF x =- 32076 THEN
            exp_f := 0;
        ELSIF x =- 32075 THEN
            exp_f := 0;
        ELSIF x =- 32074 THEN
            exp_f := 0;
        ELSIF x =- 32073 THEN
            exp_f := 0;
        ELSIF x =- 32072 THEN
            exp_f := 0;
        ELSIF x =- 32071 THEN
            exp_f := 0;
        ELSIF x =- 32070 THEN
            exp_f := 0;
        ELSIF x =- 32069 THEN
            exp_f := 0;
        ELSIF x =- 32068 THEN
            exp_f := 0;
        ELSIF x =- 32067 THEN
            exp_f := 0;
        ELSIF x =- 32066 THEN
            exp_f := 0;
        ELSIF x =- 32065 THEN
            exp_f := 0;
        ELSIF x =- 32064 THEN
            exp_f := 0;
        ELSIF x =- 32063 THEN
            exp_f := 0;
        ELSIF x =- 32062 THEN
            exp_f := 0;
        ELSIF x =- 32061 THEN
            exp_f := 0;
        ELSIF x =- 32060 THEN
            exp_f := 0;
        ELSIF x =- 32059 THEN
            exp_f := 0;
        ELSIF x =- 32058 THEN
            exp_f := 0;
        ELSIF x =- 32057 THEN
            exp_f := 0;
        ELSIF x =- 32056 THEN
            exp_f := 0;
        ELSIF x =- 32055 THEN
            exp_f := 0;
        ELSIF x =- 32054 THEN
            exp_f := 0;
        ELSIF x =- 32053 THEN
            exp_f := 0;
        ELSIF x =- 32052 THEN
            exp_f := 0;
        ELSIF x =- 32051 THEN
            exp_f := 0;
        ELSIF x =- 32050 THEN
            exp_f := 0;
        ELSIF x =- 32049 THEN
            exp_f := 0;
        ELSIF x =- 32048 THEN
            exp_f := 0;
        ELSIF x =- 32047 THEN
            exp_f := 0;
        ELSIF x =- 32046 THEN
            exp_f := 0;
        ELSIF x =- 32045 THEN
            exp_f := 0;
        ELSIF x =- 32044 THEN
            exp_f := 0;
        ELSIF x =- 32043 THEN
            exp_f := 0;
        ELSIF x =- 32042 THEN
            exp_f := 0;
        ELSIF x =- 32041 THEN
            exp_f := 0;
        ELSIF x =- 32040 THEN
            exp_f := 0;
        ELSIF x =- 32039 THEN
            exp_f := 0;
        ELSIF x =- 32038 THEN
            exp_f := 0;
        ELSIF x =- 32037 THEN
            exp_f := 0;
        ELSIF x =- 32036 THEN
            exp_f := 0;
        ELSIF x =- 32035 THEN
            exp_f := 0;
        ELSIF x =- 32034 THEN
            exp_f := 0;
        ELSIF x =- 32033 THEN
            exp_f := 0;
        ELSIF x =- 32032 THEN
            exp_f := 0;
        ELSIF x =- 32031 THEN
            exp_f := 0;
        ELSIF x =- 32030 THEN
            exp_f := 0;
        ELSIF x =- 32029 THEN
            exp_f := 0;
        ELSIF x =- 32028 THEN
            exp_f := 0;
        ELSIF x =- 32027 THEN
            exp_f := 0;
        ELSIF x =- 32026 THEN
            exp_f := 0;
        ELSIF x =- 32025 THEN
            exp_f := 0;
        ELSIF x =- 32024 THEN
            exp_f := 0;
        ELSIF x =- 32023 THEN
            exp_f := 0;
        ELSIF x =- 32022 THEN
            exp_f := 0;
        ELSIF x =- 32021 THEN
            exp_f := 0;
        ELSIF x =- 32020 THEN
            exp_f := 0;
        ELSIF x =- 32019 THEN
            exp_f := 0;
        ELSIF x =- 32018 THEN
            exp_f := 0;
        ELSIF x =- 32017 THEN
            exp_f := 0;
        ELSIF x =- 32016 THEN
            exp_f := 0;
        ELSIF x =- 32015 THEN
            exp_f := 0;
        ELSIF x =- 32014 THEN
            exp_f := 0;
        ELSIF x =- 32013 THEN
            exp_f := 0;
        ELSIF x =- 32012 THEN
            exp_f := 0;
        ELSIF x =- 32011 THEN
            exp_f := 0;
        ELSIF x =- 32010 THEN
            exp_f := 0;
        ELSIF x =- 32009 THEN
            exp_f := 0;
        ELSIF x =- 32008 THEN
            exp_f := 0;
        ELSIF x =- 32007 THEN
            exp_f := 0;
        ELSIF x =- 32006 THEN
            exp_f := 0;
        ELSIF x =- 32005 THEN
            exp_f := 0;
        ELSIF x =- 32004 THEN
            exp_f := 0;
        ELSIF x =- 32003 THEN
            exp_f := 0;
        ELSIF x =- 32002 THEN
            exp_f := 0;
        ELSIF x =- 32001 THEN
            exp_f := 0;
        ELSIF x =- 32000 THEN
            exp_f := 0;
        ELSIF x =- 31999 THEN
            exp_f := 0;
        ELSIF x =- 31998 THEN
            exp_f := 0;
        ELSIF x =- 31997 THEN
            exp_f := 0;
        ELSIF x =- 31996 THEN
            exp_f := 0;
        ELSIF x =- 31995 THEN
            exp_f := 0;
        ELSIF x =- 31994 THEN
            exp_f := 0;
        ELSIF x =- 31993 THEN
            exp_f := 0;
        ELSIF x =- 31992 THEN
            exp_f := 0;
        ELSIF x =- 31991 THEN
            exp_f := 0;
        ELSIF x =- 31990 THEN
            exp_f := 0;
        ELSIF x =- 31989 THEN
            exp_f := 0;
        ELSIF x =- 31988 THEN
            exp_f := 0;
        ELSIF x =- 31987 THEN
            exp_f := 0;
        ELSIF x =- 31986 THEN
            exp_f := 0;
        ELSIF x =- 31985 THEN
            exp_f := 0;
        ELSIF x =- 31984 THEN
            exp_f := 0;
        ELSIF x =- 31983 THEN
            exp_f := 0;
        ELSIF x =- 31982 THEN
            exp_f := 0;
        ELSIF x =- 31981 THEN
            exp_f := 0;
        ELSIF x =- 31980 THEN
            exp_f := 0;
        ELSIF x =- 31979 THEN
            exp_f := 0;
        ELSIF x =- 31978 THEN
            exp_f := 0;
        ELSIF x =- 31977 THEN
            exp_f := 0;
        ELSIF x =- 31976 THEN
            exp_f := 0;
        ELSIF x =- 31975 THEN
            exp_f := 0;
        ELSIF x =- 31974 THEN
            exp_f := 0;
        ELSIF x =- 31973 THEN
            exp_f := 0;
        ELSIF x =- 31972 THEN
            exp_f := 0;
        ELSIF x =- 31971 THEN
            exp_f := 0;
        ELSIF x =- 31970 THEN
            exp_f := 0;
        ELSIF x =- 31969 THEN
            exp_f := 0;
        ELSIF x =- 31968 THEN
            exp_f := 0;
        ELSIF x =- 31967 THEN
            exp_f := 0;
        ELSIF x =- 31966 THEN
            exp_f := 0;
        ELSIF x =- 31965 THEN
            exp_f := 0;
        ELSIF x =- 31964 THEN
            exp_f := 0;
        ELSIF x =- 31963 THEN
            exp_f := 0;
        ELSIF x =- 31962 THEN
            exp_f := 0;
        ELSIF x =- 31961 THEN
            exp_f := 0;
        ELSIF x =- 31960 THEN
            exp_f := 0;
        ELSIF x =- 31959 THEN
            exp_f := 0;
        ELSIF x =- 31958 THEN
            exp_f := 0;
        ELSIF x =- 31957 THEN
            exp_f := 0;
        ELSIF x =- 31956 THEN
            exp_f := 0;
        ELSIF x =- 31955 THEN
            exp_f := 0;
        ELSIF x =- 31954 THEN
            exp_f := 0;
        ELSIF x =- 31953 THEN
            exp_f := 0;
        ELSIF x =- 31952 THEN
            exp_f := 0;
        ELSIF x =- 31951 THEN
            exp_f := 0;
        ELSIF x =- 31950 THEN
            exp_f := 0;
        ELSIF x =- 31949 THEN
            exp_f := 0;
        ELSIF x =- 31948 THEN
            exp_f := 0;
        ELSIF x =- 31947 THEN
            exp_f := 0;
        ELSIF x =- 31946 THEN
            exp_f := 0;
        ELSIF x =- 31945 THEN
            exp_f := 0;
        ELSIF x =- 31944 THEN
            exp_f := 0;
        ELSIF x =- 31943 THEN
            exp_f := 0;
        ELSIF x =- 31942 THEN
            exp_f := 0;
        ELSIF x =- 31941 THEN
            exp_f := 0;
        ELSIF x =- 31940 THEN
            exp_f := 0;
        ELSIF x =- 31939 THEN
            exp_f := 0;
        ELSIF x =- 31938 THEN
            exp_f := 0;
        ELSIF x =- 31937 THEN
            exp_f := 0;
        ELSIF x =- 31936 THEN
            exp_f := 0;
        ELSIF x =- 31935 THEN
            exp_f := 0;
        ELSIF x =- 31934 THEN
            exp_f := 0;
        ELSIF x =- 31933 THEN
            exp_f := 0;
        ELSIF x =- 31932 THEN
            exp_f := 0;
        ELSIF x =- 31931 THEN
            exp_f := 0;
        ELSIF x =- 31930 THEN
            exp_f := 0;
        ELSIF x =- 31929 THEN
            exp_f := 0;
        ELSIF x =- 31928 THEN
            exp_f := 0;
        ELSIF x =- 31927 THEN
            exp_f := 0;
        ELSIF x =- 31926 THEN
            exp_f := 0;
        ELSIF x =- 31925 THEN
            exp_f := 0;
        ELSIF x =- 31924 THEN
            exp_f := 0;
        ELSIF x =- 31923 THEN
            exp_f := 0;
        ELSIF x =- 31922 THEN
            exp_f := 0;
        ELSIF x =- 31921 THEN
            exp_f := 0;
        ELSIF x =- 31920 THEN
            exp_f := 0;
        ELSIF x =- 31919 THEN
            exp_f := 0;
        ELSIF x =- 31918 THEN
            exp_f := 0;
        ELSIF x =- 31917 THEN
            exp_f := 0;
        ELSIF x =- 31916 THEN
            exp_f := 0;
        ELSIF x =- 31915 THEN
            exp_f := 0;
        ELSIF x =- 31914 THEN
            exp_f := 0;
        ELSIF x =- 31913 THEN
            exp_f := 0;
        ELSIF x =- 31912 THEN
            exp_f := 0;
        ELSIF x =- 31911 THEN
            exp_f := 0;
        ELSIF x =- 31910 THEN
            exp_f := 0;
        ELSIF x =- 31909 THEN
            exp_f := 0;
        ELSIF x =- 31908 THEN
            exp_f := 0;
        ELSIF x =- 31907 THEN
            exp_f := 0;
        ELSIF x =- 31906 THEN
            exp_f := 0;
        ELSIF x =- 31905 THEN
            exp_f := 0;
        ELSIF x =- 31904 THEN
            exp_f := 0;
        ELSIF x =- 31903 THEN
            exp_f := 0;
        ELSIF x =- 31902 THEN
            exp_f := 0;
        ELSIF x =- 31901 THEN
            exp_f := 0;
        ELSIF x =- 31900 THEN
            exp_f := 0;
        ELSIF x =- 31899 THEN
            exp_f := 0;
        ELSIF x =- 31898 THEN
            exp_f := 0;
        ELSIF x =- 31897 THEN
            exp_f := 0;
        ELSIF x =- 31896 THEN
            exp_f := 0;
        ELSIF x =- 31895 THEN
            exp_f := 0;
        ELSIF x =- 31894 THEN
            exp_f := 0;
        ELSIF x =- 31893 THEN
            exp_f := 0;
        ELSIF x =- 31892 THEN
            exp_f := 0;
        ELSIF x =- 31891 THEN
            exp_f := 0;
        ELSIF x =- 31890 THEN
            exp_f := 0;
        ELSIF x =- 31889 THEN
            exp_f := 0;
        ELSIF x =- 31888 THEN
            exp_f := 0;
        ELSIF x =- 31887 THEN
            exp_f := 0;
        ELSIF x =- 31886 THEN
            exp_f := 0;
        ELSIF x =- 31885 THEN
            exp_f := 0;
        ELSIF x =- 31884 THEN
            exp_f := 0;
        ELSIF x =- 31883 THEN
            exp_f := 0;
        ELSIF x =- 31882 THEN
            exp_f := 0;
        ELSIF x =- 31881 THEN
            exp_f := 0;
        ELSIF x =- 31880 THEN
            exp_f := 0;
        ELSIF x =- 31879 THEN
            exp_f := 0;
        ELSIF x =- 31878 THEN
            exp_f := 0;
        ELSIF x =- 31877 THEN
            exp_f := 0;
        ELSIF x =- 31876 THEN
            exp_f := 0;
        ELSIF x =- 31875 THEN
            exp_f := 0;
        ELSIF x =- 31874 THEN
            exp_f := 0;
        ELSIF x =- 31873 THEN
            exp_f := 0;
        ELSIF x =- 31872 THEN
            exp_f := 0;
        ELSIF x =- 31871 THEN
            exp_f := 0;
        ELSIF x =- 31870 THEN
            exp_f := 0;
        ELSIF x =- 31869 THEN
            exp_f := 0;
        ELSIF x =- 31868 THEN
            exp_f := 0;
        ELSIF x =- 31867 THEN
            exp_f := 0;
        ELSIF x =- 31866 THEN
            exp_f := 0;
        ELSIF x =- 31865 THEN
            exp_f := 0;
        ELSIF x =- 31864 THEN
            exp_f := 0;
        ELSIF x =- 31863 THEN
            exp_f := 0;
        ELSIF x =- 31862 THEN
            exp_f := 0;
        ELSIF x =- 31861 THEN
            exp_f := 0;
        ELSIF x =- 31860 THEN
            exp_f := 0;
        ELSIF x =- 31859 THEN
            exp_f := 0;
        ELSIF x =- 31858 THEN
            exp_f := 0;
        ELSIF x =- 31857 THEN
            exp_f := 0;
        ELSIF x =- 31856 THEN
            exp_f := 0;
        ELSIF x =- 31855 THEN
            exp_f := 0;
        ELSIF x =- 31854 THEN
            exp_f := 0;
        ELSIF x =- 31853 THEN
            exp_f := 0;
        ELSIF x =- 31852 THEN
            exp_f := 0;
        ELSIF x =- 31851 THEN
            exp_f := 0;
        ELSIF x =- 31850 THEN
            exp_f := 0;
        ELSIF x =- 31849 THEN
            exp_f := 0;
        ELSIF x =- 31848 THEN
            exp_f := 0;
        ELSIF x =- 31847 THEN
            exp_f := 0;
        ELSIF x =- 31846 THEN
            exp_f := 0;
        ELSIF x =- 31845 THEN
            exp_f := 0;
        ELSIF x =- 31844 THEN
            exp_f := 0;
        ELSIF x =- 31843 THEN
            exp_f := 0;
        ELSIF x =- 31842 THEN
            exp_f := 0;
        ELSIF x =- 31841 THEN
            exp_f := 0;
        ELSIF x =- 31840 THEN
            exp_f := 0;
        ELSIF x =- 31839 THEN
            exp_f := 0;
        ELSIF x =- 31838 THEN
            exp_f := 0;
        ELSIF x =- 31837 THEN
            exp_f := 0;
        ELSIF x =- 31836 THEN
            exp_f := 0;
        ELSIF x =- 31835 THEN
            exp_f := 0;
        ELSIF x =- 31834 THEN
            exp_f := 0;
        ELSIF x =- 31833 THEN
            exp_f := 0;
        ELSIF x =- 31832 THEN
            exp_f := 0;
        ELSIF x =- 31831 THEN
            exp_f := 0;
        ELSIF x =- 31830 THEN
            exp_f := 0;
        ELSIF x =- 31829 THEN
            exp_f := 0;
        ELSIF x =- 31828 THEN
            exp_f := 0;
        ELSIF x =- 31827 THEN
            exp_f := 0;
        ELSIF x =- 31826 THEN
            exp_f := 0;
        ELSIF x =- 31825 THEN
            exp_f := 0;
        ELSIF x =- 31824 THEN
            exp_f := 0;
        ELSIF x =- 31823 THEN
            exp_f := 0;
        ELSIF x =- 31822 THEN
            exp_f := 0;
        ELSIF x =- 31821 THEN
            exp_f := 0;
        ELSIF x =- 31820 THEN
            exp_f := 0;
        ELSIF x =- 31819 THEN
            exp_f := 0;
        ELSIF x =- 31818 THEN
            exp_f := 0;
        ELSIF x =- 31817 THEN
            exp_f := 0;
        ELSIF x =- 31816 THEN
            exp_f := 0;
        ELSIF x =- 31815 THEN
            exp_f := 0;
        ELSIF x =- 31814 THEN
            exp_f := 0;
        ELSIF x =- 31813 THEN
            exp_f := 0;
        ELSIF x =- 31812 THEN
            exp_f := 0;
        ELSIF x =- 31811 THEN
            exp_f := 0;
        ELSIF x =- 31810 THEN
            exp_f := 0;
        ELSIF x =- 31809 THEN
            exp_f := 0;
        ELSIF x =- 31808 THEN
            exp_f := 0;
        ELSIF x =- 31807 THEN
            exp_f := 0;
        ELSIF x =- 31806 THEN
            exp_f := 0;
        ELSIF x =- 31805 THEN
            exp_f := 0;
        ELSIF x =- 31804 THEN
            exp_f := 0;
        ELSIF x =- 31803 THEN
            exp_f := 0;
        ELSIF x =- 31802 THEN
            exp_f := 0;
        ELSIF x =- 31801 THEN
            exp_f := 0;
        ELSIF x =- 31800 THEN
            exp_f := 0;
        ELSIF x =- 31799 THEN
            exp_f := 0;
        ELSIF x =- 31798 THEN
            exp_f := 0;
        ELSIF x =- 31797 THEN
            exp_f := 0;
        ELSIF x =- 31796 THEN
            exp_f := 0;
        ELSIF x =- 31795 THEN
            exp_f := 0;
        ELSIF x =- 31794 THEN
            exp_f := 0;
        ELSIF x =- 31793 THEN
            exp_f := 0;
        ELSIF x =- 31792 THEN
            exp_f := 0;
        ELSIF x =- 31791 THEN
            exp_f := 0;
        ELSIF x =- 31790 THEN
            exp_f := 0;
        ELSIF x =- 31789 THEN
            exp_f := 0;
        ELSIF x =- 31788 THEN
            exp_f := 0;
        ELSIF x =- 31787 THEN
            exp_f := 0;
        ELSIF x =- 31786 THEN
            exp_f := 0;
        ELSIF x =- 31785 THEN
            exp_f := 0;
        ELSIF x =- 31784 THEN
            exp_f := 0;
        ELSIF x =- 31783 THEN
            exp_f := 0;
        ELSIF x =- 31782 THEN
            exp_f := 0;
        ELSIF x =- 31781 THEN
            exp_f := 0;
        ELSIF x =- 31780 THEN
            exp_f := 0;
        ELSIF x =- 31779 THEN
            exp_f := 0;
        ELSIF x =- 31778 THEN
            exp_f := 0;
        ELSIF x =- 31777 THEN
            exp_f := 0;
        ELSIF x =- 31776 THEN
            exp_f := 0;
        ELSIF x =- 31775 THEN
            exp_f := 0;
        ELSIF x =- 31774 THEN
            exp_f := 0;
        ELSIF x =- 31773 THEN
            exp_f := 0;
        ELSIF x =- 31772 THEN
            exp_f := 0;
        ELSIF x =- 31771 THEN
            exp_f := 0;
        ELSIF x =- 31770 THEN
            exp_f := 0;
        ELSIF x =- 31769 THEN
            exp_f := 0;
        ELSIF x =- 31768 THEN
            exp_f := 0;
        ELSIF x =- 31767 THEN
            exp_f := 0;
        ELSIF x =- 31766 THEN
            exp_f := 0;
        ELSIF x =- 31765 THEN
            exp_f := 0;
        ELSIF x =- 31764 THEN
            exp_f := 0;
        ELSIF x =- 31763 THEN
            exp_f := 0;
        ELSIF x =- 31762 THEN
            exp_f := 0;
        ELSIF x =- 31761 THEN
            exp_f := 0;
        ELSIF x =- 31760 THEN
            exp_f := 0;
        ELSIF x =- 31759 THEN
            exp_f := 0;
        ELSIF x =- 31758 THEN
            exp_f := 0;
        ELSIF x =- 31757 THEN
            exp_f := 0;
        ELSIF x =- 31756 THEN
            exp_f := 0;
        ELSIF x =- 31755 THEN
            exp_f := 0;
        ELSIF x =- 31754 THEN
            exp_f := 0;
        ELSIF x =- 31753 THEN
            exp_f := 0;
        ELSIF x =- 31752 THEN
            exp_f := 0;
        ELSIF x =- 31751 THEN
            exp_f := 0;
        ELSIF x =- 31750 THEN
            exp_f := 0;
        ELSIF x =- 31749 THEN
            exp_f := 0;
        ELSIF x =- 31748 THEN
            exp_f := 0;
        ELSIF x =- 31747 THEN
            exp_f := 0;
        ELSIF x =- 31746 THEN
            exp_f := 0;
        ELSIF x =- 31745 THEN
            exp_f := 0;
        ELSIF x =- 31744 THEN
            exp_f := 0;
        ELSIF x =- 31743 THEN
            exp_f := 0;
        ELSIF x =- 31742 THEN
            exp_f := 0;
        ELSIF x =- 31741 THEN
            exp_f := 0;
        ELSIF x =- 31740 THEN
            exp_f := 0;
        ELSIF x =- 31739 THEN
            exp_f := 0;
        ELSIF x =- 31738 THEN
            exp_f := 0;
        ELSIF x =- 31737 THEN
            exp_f := 0;
        ELSIF x =- 31736 THEN
            exp_f := 0;
        ELSIF x =- 31735 THEN
            exp_f := 0;
        ELSIF x =- 31734 THEN
            exp_f := 0;
        ELSIF x =- 31733 THEN
            exp_f := 0;
        ELSIF x =- 31732 THEN
            exp_f := 0;
        ELSIF x =- 31731 THEN
            exp_f := 0;
        ELSIF x =- 31730 THEN
            exp_f := 0;
        ELSIF x =- 31729 THEN
            exp_f := 0;
        ELSIF x =- 31728 THEN
            exp_f := 0;
        ELSIF x =- 31727 THEN
            exp_f := 0;
        ELSIF x =- 31726 THEN
            exp_f := 0;
        ELSIF x =- 31725 THEN
            exp_f := 0;
        ELSIF x =- 31724 THEN
            exp_f := 0;
        ELSIF x =- 31723 THEN
            exp_f := 0;
        ELSIF x =- 31722 THEN
            exp_f := 0;
        ELSIF x =- 31721 THEN
            exp_f := 0;
        ELSIF x =- 31720 THEN
            exp_f := 0;
        ELSIF x =- 31719 THEN
            exp_f := 0;
        ELSIF x =- 31718 THEN
            exp_f := 0;
        ELSIF x =- 31717 THEN
            exp_f := 0;
        ELSIF x =- 31716 THEN
            exp_f := 0;
        ELSIF x =- 31715 THEN
            exp_f := 0;
        ELSIF x =- 31714 THEN
            exp_f := 0;
        ELSIF x =- 31713 THEN
            exp_f := 0;
        ELSIF x =- 31712 THEN
            exp_f := 0;
        ELSIF x =- 31711 THEN
            exp_f := 0;
        ELSIF x =- 31710 THEN
            exp_f := 0;
        ELSIF x =- 31709 THEN
            exp_f := 0;
        ELSIF x =- 31708 THEN
            exp_f := 0;
        ELSIF x =- 31707 THEN
            exp_f := 0;
        ELSIF x =- 31706 THEN
            exp_f := 0;
        ELSIF x =- 31705 THEN
            exp_f := 0;
        ELSIF x =- 31704 THEN
            exp_f := 0;
        ELSIF x =- 31703 THEN
            exp_f := 0;
        ELSIF x =- 31702 THEN
            exp_f := 0;
        ELSIF x =- 31701 THEN
            exp_f := 0;
        ELSIF x =- 31700 THEN
            exp_f := 0;
        ELSIF x =- 31699 THEN
            exp_f := 0;
        ELSIF x =- 31698 THEN
            exp_f := 0;
        ELSIF x =- 31697 THEN
            exp_f := 0;
        ELSIF x =- 31696 THEN
            exp_f := 0;
        ELSIF x =- 31695 THEN
            exp_f := 0;
        ELSIF x =- 31694 THEN
            exp_f := 0;
        ELSIF x =- 31693 THEN
            exp_f := 0;
        ELSIF x =- 31692 THEN
            exp_f := 0;
        ELSIF x =- 31691 THEN
            exp_f := 0;
        ELSIF x =- 31690 THEN
            exp_f := 0;
        ELSIF x =- 31689 THEN
            exp_f := 0;
        ELSIF x =- 31688 THEN
            exp_f := 0;
        ELSIF x =- 31687 THEN
            exp_f := 0;
        ELSIF x =- 31686 THEN
            exp_f := 0;
        ELSIF x =- 31685 THEN
            exp_f := 0;
        ELSIF x =- 31684 THEN
            exp_f := 0;
        ELSIF x =- 31683 THEN
            exp_f := 0;
        ELSIF x =- 31682 THEN
            exp_f := 0;
        ELSIF x =- 31681 THEN
            exp_f := 0;
        ELSIF x =- 31680 THEN
            exp_f := 0;
        ELSIF x =- 31679 THEN
            exp_f := 0;
        ELSIF x =- 31678 THEN
            exp_f := 0;
        ELSIF x =- 31677 THEN
            exp_f := 0;
        ELSIF x =- 31676 THEN
            exp_f := 0;
        ELSIF x =- 31675 THEN
            exp_f := 0;
        ELSIF x =- 31674 THEN
            exp_f := 0;
        ELSIF x =- 31673 THEN
            exp_f := 0;
        ELSIF x =- 31672 THEN
            exp_f := 0;
        ELSIF x =- 31671 THEN
            exp_f := 0;
        ELSIF x =- 31670 THEN
            exp_f := 0;
        ELSIF x =- 31669 THEN
            exp_f := 0;
        ELSIF x =- 31668 THEN
            exp_f := 0;
        ELSIF x =- 31667 THEN
            exp_f := 0;
        ELSIF x =- 31666 THEN
            exp_f := 0;
        ELSIF x =- 31665 THEN
            exp_f := 0;
        ELSIF x =- 31664 THEN
            exp_f := 0;
        ELSIF x =- 31663 THEN
            exp_f := 0;
        ELSIF x =- 31662 THEN
            exp_f := 0;
        ELSIF x =- 31661 THEN
            exp_f := 0;
        ELSIF x =- 31660 THEN
            exp_f := 0;
        ELSIF x =- 31659 THEN
            exp_f := 0;
        ELSIF x =- 31658 THEN
            exp_f := 0;
        ELSIF x =- 31657 THEN
            exp_f := 0;
        ELSIF x =- 31656 THEN
            exp_f := 0;
        ELSIF x =- 31655 THEN
            exp_f := 0;
        ELSIF x =- 31654 THEN
            exp_f := 0;
        ELSIF x =- 31653 THEN
            exp_f := 0;
        ELSIF x =- 31652 THEN
            exp_f := 0;
        ELSIF x =- 31651 THEN
            exp_f := 0;
        ELSIF x =- 31650 THEN
            exp_f := 0;
        ELSIF x =- 31649 THEN
            exp_f := 0;
        ELSIF x =- 31648 THEN
            exp_f := 0;
        ELSIF x =- 31647 THEN
            exp_f := 0;
        ELSIF x =- 31646 THEN
            exp_f := 0;
        ELSIF x =- 31645 THEN
            exp_f := 0;
        ELSIF x =- 31644 THEN
            exp_f := 0;
        ELSIF x =- 31643 THEN
            exp_f := 0;
        ELSIF x =- 31642 THEN
            exp_f := 0;
        ELSIF x =- 31641 THEN
            exp_f := 0;
        ELSIF x =- 31640 THEN
            exp_f := 0;
        ELSIF x =- 31639 THEN
            exp_f := 0;
        ELSIF x =- 31638 THEN
            exp_f := 0;
        ELSIF x =- 31637 THEN
            exp_f := 0;
        ELSIF x =- 31636 THEN
            exp_f := 0;
        ELSIF x =- 31635 THEN
            exp_f := 0;
        ELSIF x =- 31634 THEN
            exp_f := 0;
        ELSIF x =- 31633 THEN
            exp_f := 0;
        ELSIF x =- 31632 THEN
            exp_f := 0;
        ELSIF x =- 31631 THEN
            exp_f := 0;
        ELSIF x =- 31630 THEN
            exp_f := 0;
        ELSIF x =- 31629 THEN
            exp_f := 0;
        ELSIF x =- 31628 THEN
            exp_f := 0;
        ELSIF x =- 31627 THEN
            exp_f := 0;
        ELSIF x =- 31626 THEN
            exp_f := 0;
        ELSIF x =- 31625 THEN
            exp_f := 0;
        ELSIF x =- 31624 THEN
            exp_f := 0;
        ELSIF x =- 31623 THEN
            exp_f := 0;
        ELSIF x =- 31622 THEN
            exp_f := 0;
        ELSIF x =- 31621 THEN
            exp_f := 0;
        ELSIF x =- 31620 THEN
            exp_f := 0;
        ELSIF x =- 31619 THEN
            exp_f := 0;
        ELSIF x =- 31618 THEN
            exp_f := 0;
        ELSIF x =- 31617 THEN
            exp_f := 0;
        ELSIF x =- 31616 THEN
            exp_f := 0;
        ELSIF x =- 31615 THEN
            exp_f := 0;
        ELSIF x =- 31614 THEN
            exp_f := 0;
        ELSIF x =- 31613 THEN
            exp_f := 0;
        ELSIF x =- 31612 THEN
            exp_f := 0;
        ELSIF x =- 31611 THEN
            exp_f := 0;
        ELSIF x =- 31610 THEN
            exp_f := 0;
        ELSIF x =- 31609 THEN
            exp_f := 0;
        ELSIF x =- 31608 THEN
            exp_f := 0;
        ELSIF x =- 31607 THEN
            exp_f := 0;
        ELSIF x =- 31606 THEN
            exp_f := 0;
        ELSIF x =- 31605 THEN
            exp_f := 0;
        ELSIF x =- 31604 THEN
            exp_f := 0;
        ELSIF x =- 31603 THEN
            exp_f := 0;
        ELSIF x =- 31602 THEN
            exp_f := 0;
        ELSIF x =- 31601 THEN
            exp_f := 0;
        ELSIF x =- 31600 THEN
            exp_f := 0;
        ELSIF x =- 31599 THEN
            exp_f := 0;
        ELSIF x =- 31598 THEN
            exp_f := 0;
        ELSIF x =- 31597 THEN
            exp_f := 0;
        ELSIF x =- 31596 THEN
            exp_f := 0;
        ELSIF x =- 31595 THEN
            exp_f := 0;
        ELSIF x =- 31594 THEN
            exp_f := 0;
        ELSIF x =- 31593 THEN
            exp_f := 0;
        ELSIF x =- 31592 THEN
            exp_f := 0;
        ELSIF x =- 31591 THEN
            exp_f := 0;
        ELSIF x =- 31590 THEN
            exp_f := 0;
        ELSIF x =- 31589 THEN
            exp_f := 0;
        ELSIF x =- 31588 THEN
            exp_f := 0;
        ELSIF x =- 31587 THEN
            exp_f := 0;
        ELSIF x =- 31586 THEN
            exp_f := 0;
        ELSIF x =- 31585 THEN
            exp_f := 0;
        ELSIF x =- 31584 THEN
            exp_f := 0;
        ELSIF x =- 31583 THEN
            exp_f := 0;
        ELSIF x =- 31582 THEN
            exp_f := 0;
        ELSIF x =- 31581 THEN
            exp_f := 0;
        ELSIF x =- 31580 THEN
            exp_f := 0;
        ELSIF x =- 31579 THEN
            exp_f := 0;
        ELSIF x =- 31578 THEN
            exp_f := 0;
        ELSIF x =- 31577 THEN
            exp_f := 0;
        ELSIF x =- 31576 THEN
            exp_f := 0;
        ELSIF x =- 31575 THEN
            exp_f := 0;
        ELSIF x =- 31574 THEN
            exp_f := 0;
        ELSIF x =- 31573 THEN
            exp_f := 0;
        ELSIF x =- 31572 THEN
            exp_f := 0;
        ELSIF x =- 31571 THEN
            exp_f := 0;
        ELSIF x =- 31570 THEN
            exp_f := 0;
        ELSIF x =- 31569 THEN
            exp_f := 0;
        ELSIF x =- 31568 THEN
            exp_f := 0;
        ELSIF x =- 31567 THEN
            exp_f := 0;
        ELSIF x =- 31566 THEN
            exp_f := 0;
        ELSIF x =- 31565 THEN
            exp_f := 0;
        ELSIF x =- 31564 THEN
            exp_f := 0;
        ELSIF x =- 31563 THEN
            exp_f := 0;
        ELSIF x =- 31562 THEN
            exp_f := 0;
        ELSIF x =- 31561 THEN
            exp_f := 0;
        ELSIF x =- 31560 THEN
            exp_f := 0;
        ELSIF x =- 31559 THEN
            exp_f := 0;
        ELSIF x =- 31558 THEN
            exp_f := 0;
        ELSIF x =- 31557 THEN
            exp_f := 0;
        ELSIF x =- 31556 THEN
            exp_f := 0;
        ELSIF x =- 31555 THEN
            exp_f := 0;
        ELSIF x =- 31554 THEN
            exp_f := 0;
        ELSIF x =- 31553 THEN
            exp_f := 0;
        ELSIF x =- 31552 THEN
            exp_f := 0;
        ELSIF x =- 31551 THEN
            exp_f := 0;
        ELSIF x =- 31550 THEN
            exp_f := 0;
        ELSIF x =- 31549 THEN
            exp_f := 0;
        ELSIF x =- 31548 THEN
            exp_f := 0;
        ELSIF x =- 31547 THEN
            exp_f := 0;
        ELSIF x =- 31546 THEN
            exp_f := 0;
        ELSIF x =- 31545 THEN
            exp_f := 0;
        ELSIF x =- 31544 THEN
            exp_f := 0;
        ELSIF x =- 31543 THEN
            exp_f := 0;
        ELSIF x =- 31542 THEN
            exp_f := 0;
        ELSIF x =- 31541 THEN
            exp_f := 0;
        ELSIF x =- 31540 THEN
            exp_f := 0;
        ELSIF x =- 31539 THEN
            exp_f := 0;
        ELSIF x =- 31538 THEN
            exp_f := 0;
        ELSIF x =- 31537 THEN
            exp_f := 0;
        ELSIF x =- 31536 THEN
            exp_f := 0;
        ELSIF x =- 31535 THEN
            exp_f := 0;
        ELSIF x =- 31534 THEN
            exp_f := 0;
        ELSIF x =- 31533 THEN
            exp_f := 0;
        ELSIF x =- 31532 THEN
            exp_f := 0;
        ELSIF x =- 31531 THEN
            exp_f := 0;
        ELSIF x =- 31530 THEN
            exp_f := 0;
        ELSIF x =- 31529 THEN
            exp_f := 0;
        ELSIF x =- 31528 THEN
            exp_f := 0;
        ELSIF x =- 31527 THEN
            exp_f := 0;
        ELSIF x =- 31526 THEN
            exp_f := 0;
        ELSIF x =- 31525 THEN
            exp_f := 0;
        ELSIF x =- 31524 THEN
            exp_f := 0;
        ELSIF x =- 31523 THEN
            exp_f := 0;
        ELSIF x =- 31522 THEN
            exp_f := 0;
        ELSIF x =- 31521 THEN
            exp_f := 0;
        ELSIF x =- 31520 THEN
            exp_f := 0;
        ELSIF x =- 31519 THEN
            exp_f := 0;
        ELSIF x =- 31518 THEN
            exp_f := 0;
        ELSIF x =- 31517 THEN
            exp_f := 0;
        ELSIF x =- 31516 THEN
            exp_f := 0;
        ELSIF x =- 31515 THEN
            exp_f := 0;
        ELSIF x =- 31514 THEN
            exp_f := 0;
        ELSIF x =- 31513 THEN
            exp_f := 0;
        ELSIF x =- 31512 THEN
            exp_f := 0;
        ELSIF x =- 31511 THEN
            exp_f := 0;
        ELSIF x =- 31510 THEN
            exp_f := 0;
        ELSIF x =- 31509 THEN
            exp_f := 0;
        ELSIF x =- 31508 THEN
            exp_f := 0;
        ELSIF x =- 31507 THEN
            exp_f := 0;
        ELSIF x =- 31506 THEN
            exp_f := 0;
        ELSIF x =- 31505 THEN
            exp_f := 0;
        ELSIF x =- 31504 THEN
            exp_f := 0;
        ELSIF x =- 31503 THEN
            exp_f := 0;
        ELSIF x =- 31502 THEN
            exp_f := 0;
        ELSIF x =- 31501 THEN
            exp_f := 0;
        ELSIF x =- 31500 THEN
            exp_f := 0;
        ELSIF x =- 31499 THEN
            exp_f := 0;
        ELSIF x =- 31498 THEN
            exp_f := 0;
        ELSIF x =- 31497 THEN
            exp_f := 0;
        ELSIF x =- 31496 THEN
            exp_f := 0;
        ELSIF x =- 31495 THEN
            exp_f := 0;
        ELSIF x =- 31494 THEN
            exp_f := 0;
        ELSIF x =- 31493 THEN
            exp_f := 0;
        ELSIF x =- 31492 THEN
            exp_f := 0;
        ELSIF x =- 31491 THEN
            exp_f := 0;
        ELSIF x =- 31490 THEN
            exp_f := 0;
        ELSIF x =- 31489 THEN
            exp_f := 0;
        ELSIF x =- 31488 THEN
            exp_f := 0;
        ELSIF x =- 31487 THEN
            exp_f := 0;
        ELSIF x =- 31486 THEN
            exp_f := 0;
        ELSIF x =- 31485 THEN
            exp_f := 0;
        ELSIF x =- 31484 THEN
            exp_f := 0;
        ELSIF x =- 31483 THEN
            exp_f := 0;
        ELSIF x =- 31482 THEN
            exp_f := 0;
        ELSIF x =- 31481 THEN
            exp_f := 0;
        ELSIF x =- 31480 THEN
            exp_f := 0;
        ELSIF x =- 31479 THEN
            exp_f := 0;
        ELSIF x =- 31478 THEN
            exp_f := 0;
        ELSIF x =- 31477 THEN
            exp_f := 0;
        ELSIF x =- 31476 THEN
            exp_f := 0;
        ELSIF x =- 31475 THEN
            exp_f := 0;
        ELSIF x =- 31474 THEN
            exp_f := 0;
        ELSIF x =- 31473 THEN
            exp_f := 0;
        ELSIF x =- 31472 THEN
            exp_f := 0;
        ELSIF x =- 31471 THEN
            exp_f := 0;
        ELSIF x =- 31470 THEN
            exp_f := 0;
        ELSIF x =- 31469 THEN
            exp_f := 0;
        ELSIF x =- 31468 THEN
            exp_f := 0;
        ELSIF x =- 31467 THEN
            exp_f := 0;
        ELSIF x =- 31466 THEN
            exp_f := 0;
        ELSIF x =- 31465 THEN
            exp_f := 0;
        ELSIF x =- 31464 THEN
            exp_f := 0;
        ELSIF x =- 31463 THEN
            exp_f := 0;
        ELSIF x =- 31462 THEN
            exp_f := 0;
        ELSIF x =- 31461 THEN
            exp_f := 0;
        ELSIF x =- 31460 THEN
            exp_f := 0;
        ELSIF x =- 31459 THEN
            exp_f := 0;
        ELSIF x =- 31458 THEN
            exp_f := 0;
        ELSIF x =- 31457 THEN
            exp_f := 0;
        ELSIF x =- 31456 THEN
            exp_f := 0;
        ELSIF x =- 31455 THEN
            exp_f := 0;
        ELSIF x =- 31454 THEN
            exp_f := 0;
        ELSIF x =- 31453 THEN
            exp_f := 0;
        ELSIF x =- 31452 THEN
            exp_f := 0;
        ELSIF x =- 31451 THEN
            exp_f := 0;
        ELSIF x =- 31450 THEN
            exp_f := 0;
        ELSIF x =- 31449 THEN
            exp_f := 0;
        ELSIF x =- 31448 THEN
            exp_f := 0;
        ELSIF x =- 31447 THEN
            exp_f := 0;
        ELSIF x =- 31446 THEN
            exp_f := 0;
        ELSIF x =- 31445 THEN
            exp_f := 0;
        ELSIF x =- 31444 THEN
            exp_f := 0;
        ELSIF x =- 31443 THEN
            exp_f := 0;
        ELSIF x =- 31442 THEN
            exp_f := 0;
        ELSIF x =- 31441 THEN
            exp_f := 0;
        ELSIF x =- 31440 THEN
            exp_f := 0;
        ELSIF x =- 31439 THEN
            exp_f := 0;
        ELSIF x =- 31438 THEN
            exp_f := 0;
        ELSIF x =- 31437 THEN
            exp_f := 0;
        ELSIF x =- 31436 THEN
            exp_f := 0;
        ELSIF x =- 31435 THEN
            exp_f := 0;
        ELSIF x =- 31434 THEN
            exp_f := 0;
        ELSIF x =- 31433 THEN
            exp_f := 0;
        ELSIF x =- 31432 THEN
            exp_f := 0;
        ELSIF x =- 31431 THEN
            exp_f := 0;
        ELSIF x =- 31430 THEN
            exp_f := 0;
        ELSIF x =- 31429 THEN
            exp_f := 0;
        ELSIF x =- 31428 THEN
            exp_f := 0;
        ELSIF x =- 31427 THEN
            exp_f := 0;
        ELSIF x =- 31426 THEN
            exp_f := 0;
        ELSIF x =- 31425 THEN
            exp_f := 0;
        ELSIF x =- 31424 THEN
            exp_f := 0;
        ELSIF x =- 31423 THEN
            exp_f := 0;
        ELSIF x =- 31422 THEN
            exp_f := 0;
        ELSIF x =- 31421 THEN
            exp_f := 0;
        ELSIF x =- 31420 THEN
            exp_f := 0;
        ELSIF x =- 31419 THEN
            exp_f := 0;
        ELSIF x =- 31418 THEN
            exp_f := 0;
        ELSIF x =- 31417 THEN
            exp_f := 0;
        ELSIF x =- 31416 THEN
            exp_f := 0;
        ELSIF x =- 31415 THEN
            exp_f := 0;
        ELSIF x =- 31414 THEN
            exp_f := 0;
        ELSIF x =- 31413 THEN
            exp_f := 0;
        ELSIF x =- 31412 THEN
            exp_f := 0;
        ELSIF x =- 31411 THEN
            exp_f := 0;
        ELSIF x =- 31410 THEN
            exp_f := 0;
        ELSIF x =- 31409 THEN
            exp_f := 0;
        ELSIF x =- 31408 THEN
            exp_f := 0;
        ELSIF x =- 31407 THEN
            exp_f := 0;
        ELSIF x =- 31406 THEN
            exp_f := 0;
        ELSIF x =- 31405 THEN
            exp_f := 0;
        ELSIF x =- 31404 THEN
            exp_f := 0;
        ELSIF x =- 31403 THEN
            exp_f := 0;
        ELSIF x =- 31402 THEN
            exp_f := 0;
        ELSIF x =- 31401 THEN
            exp_f := 0;
        ELSIF x =- 31400 THEN
            exp_f := 0;
        ELSIF x =- 31399 THEN
            exp_f := 0;
        ELSIF x =- 31398 THEN
            exp_f := 0;
        ELSIF x =- 31397 THEN
            exp_f := 0;
        ELSIF x =- 31396 THEN
            exp_f := 0;
        ELSIF x =- 31395 THEN
            exp_f := 0;
        ELSIF x =- 31394 THEN
            exp_f := 0;
        ELSIF x =- 31393 THEN
            exp_f := 0;
        ELSIF x =- 31392 THEN
            exp_f := 0;
        ELSIF x =- 31391 THEN
            exp_f := 0;
        ELSIF x =- 31390 THEN
            exp_f := 0;
        ELSIF x =- 31389 THEN
            exp_f := 0;
        ELSIF x =- 31388 THEN
            exp_f := 0;
        ELSIF x =- 31387 THEN
            exp_f := 0;
        ELSIF x =- 31386 THEN
            exp_f := 0;
        ELSIF x =- 31385 THEN
            exp_f := 0;
        ELSIF x =- 31384 THEN
            exp_f := 0;
        ELSIF x =- 31383 THEN
            exp_f := 0;
        ELSIF x =- 31382 THEN
            exp_f := 0;
        ELSIF x =- 31381 THEN
            exp_f := 0;
        ELSIF x =- 31380 THEN
            exp_f := 0;
        ELSIF x =- 31379 THEN
            exp_f := 0;
        ELSIF x =- 31378 THEN
            exp_f := 0;
        ELSIF x =- 31377 THEN
            exp_f := 0;
        ELSIF x =- 31376 THEN
            exp_f := 0;
        ELSIF x =- 31375 THEN
            exp_f := 0;
        ELSIF x =- 31374 THEN
            exp_f := 0;
        ELSIF x =- 31373 THEN
            exp_f := 0;
        ELSIF x =- 31372 THEN
            exp_f := 0;
        ELSIF x =- 31371 THEN
            exp_f := 0;
        ELSIF x =- 31370 THEN
            exp_f := 0;
        ELSIF x =- 31369 THEN
            exp_f := 0;
        ELSIF x =- 31368 THEN
            exp_f := 0;
        ELSIF x =- 31367 THEN
            exp_f := 0;
        ELSIF x =- 31366 THEN
            exp_f := 0;
        ELSIF x =- 31365 THEN
            exp_f := 0;
        ELSIF x =- 31364 THEN
            exp_f := 0;
        ELSIF x =- 31363 THEN
            exp_f := 0;
        ELSIF x =- 31362 THEN
            exp_f := 0;
        ELSIF x =- 31361 THEN
            exp_f := 0;
        ELSIF x =- 31360 THEN
            exp_f := 0;
        ELSIF x =- 31359 THEN
            exp_f := 0;
        ELSIF x =- 31358 THEN
            exp_f := 0;
        ELSIF x =- 31357 THEN
            exp_f := 0;
        ELSIF x =- 31356 THEN
            exp_f := 0;
        ELSIF x =- 31355 THEN
            exp_f := 0;
        ELSIF x =- 31354 THEN
            exp_f := 0;
        ELSIF x =- 31353 THEN
            exp_f := 0;
        ELSIF x =- 31352 THEN
            exp_f := 0;
        ELSIF x =- 31351 THEN
            exp_f := 0;
        ELSIF x =- 31350 THEN
            exp_f := 0;
        ELSIF x =- 31349 THEN
            exp_f := 0;
        ELSIF x =- 31348 THEN
            exp_f := 0;
        ELSIF x =- 31347 THEN
            exp_f := 0;
        ELSIF x =- 31346 THEN
            exp_f := 0;
        ELSIF x =- 31345 THEN
            exp_f := 0;
        ELSIF x =- 31344 THEN
            exp_f := 0;
        ELSIF x =- 31343 THEN
            exp_f := 0;
        ELSIF x =- 31342 THEN
            exp_f := 0;
        ELSIF x =- 31341 THEN
            exp_f := 0;
        ELSIF x =- 31340 THEN
            exp_f := 0;
        ELSIF x =- 31339 THEN
            exp_f := 0;
        ELSIF x =- 31338 THEN
            exp_f := 0;
        ELSIF x =- 31337 THEN
            exp_f := 0;
        ELSIF x =- 31336 THEN
            exp_f := 0;
        ELSIF x =- 31335 THEN
            exp_f := 0;
        ELSIF x =- 31334 THEN
            exp_f := 0;
        ELSIF x =- 31333 THEN
            exp_f := 0;
        ELSIF x =- 31332 THEN
            exp_f := 0;
        ELSIF x =- 31331 THEN
            exp_f := 0;
        ELSIF x =- 31330 THEN
            exp_f := 0;
        ELSIF x =- 31329 THEN
            exp_f := 0;
        ELSIF x =- 31328 THEN
            exp_f := 0;
        ELSIF x =- 31327 THEN
            exp_f := 0;
        ELSIF x =- 31326 THEN
            exp_f := 0;
        ELSIF x =- 31325 THEN
            exp_f := 0;
        ELSIF x =- 31324 THEN
            exp_f := 0;
        ELSIF x =- 31323 THEN
            exp_f := 0;
        ELSIF x =- 31322 THEN
            exp_f := 0;
        ELSIF x =- 31321 THEN
            exp_f := 0;
        ELSIF x =- 31320 THEN
            exp_f := 0;
        ELSIF x =- 31319 THEN
            exp_f := 0;
        ELSIF x =- 31318 THEN
            exp_f := 0;
        ELSIF x =- 31317 THEN
            exp_f := 0;
        ELSIF x =- 31316 THEN
            exp_f := 0;
        ELSIF x =- 31315 THEN
            exp_f := 0;
        ELSIF x =- 31314 THEN
            exp_f := 0;
        ELSIF x =- 31313 THEN
            exp_f := 0;
        ELSIF x =- 31312 THEN
            exp_f := 0;
        ELSIF x =- 31311 THEN
            exp_f := 0;
        ELSIF x =- 31310 THEN
            exp_f := 0;
        ELSIF x =- 31309 THEN
            exp_f := 0;
        ELSIF x =- 31308 THEN
            exp_f := 0;
        ELSIF x =- 31307 THEN
            exp_f := 0;
        ELSIF x =- 31306 THEN
            exp_f := 0;
        ELSIF x =- 31305 THEN
            exp_f := 0;
        ELSIF x =- 31304 THEN
            exp_f := 0;
        ELSIF x =- 31303 THEN
            exp_f := 0;
        ELSIF x =- 31302 THEN
            exp_f := 0;
        ELSIF x =- 31301 THEN
            exp_f := 0;
        ELSIF x =- 31300 THEN
            exp_f := 0;
        ELSIF x =- 31299 THEN
            exp_f := 0;
        ELSIF x =- 31298 THEN
            exp_f := 0;
        ELSIF x =- 31297 THEN
            exp_f := 0;
        ELSIF x =- 31296 THEN
            exp_f := 0;
        ELSIF x =- 31295 THEN
            exp_f := 0;
        ELSIF x =- 31294 THEN
            exp_f := 0;
        ELSIF x =- 31293 THEN
            exp_f := 0;
        ELSIF x =- 31292 THEN
            exp_f := 0;
        ELSIF x =- 31291 THEN
            exp_f := 0;
        ELSIF x =- 31290 THEN
            exp_f := 0;
        ELSIF x =- 31289 THEN
            exp_f := 0;
        ELSIF x =- 31288 THEN
            exp_f := 0;
        ELSIF x =- 31287 THEN
            exp_f := 0;
        ELSIF x =- 31286 THEN
            exp_f := 0;
        ELSIF x =- 31285 THEN
            exp_f := 0;
        ELSIF x =- 31284 THEN
            exp_f := 0;
        ELSIF x =- 31283 THEN
            exp_f := 0;
        ELSIF x =- 31282 THEN
            exp_f := 0;
        ELSIF x =- 31281 THEN
            exp_f := 0;
        ELSIF x =- 31280 THEN
            exp_f := 0;
        ELSIF x =- 31279 THEN
            exp_f := 0;
        ELSIF x =- 31278 THEN
            exp_f := 0;
        ELSIF x =- 31277 THEN
            exp_f := 0;
        ELSIF x =- 31276 THEN
            exp_f := 0;
        ELSIF x =- 31275 THEN
            exp_f := 0;
        ELSIF x =- 31274 THEN
            exp_f := 0;
        ELSIF x =- 31273 THEN
            exp_f := 0;
        ELSIF x =- 31272 THEN
            exp_f := 0;
        ELSIF x =- 31271 THEN
            exp_f := 0;
        ELSIF x =- 31270 THEN
            exp_f := 0;
        ELSIF x =- 31269 THEN
            exp_f := 0;
        ELSIF x =- 31268 THEN
            exp_f := 0;
        ELSIF x =- 31267 THEN
            exp_f := 0;
        ELSIF x =- 31266 THEN
            exp_f := 0;
        ELSIF x =- 31265 THEN
            exp_f := 0;
        ELSIF x =- 31264 THEN
            exp_f := 0;
        ELSIF x =- 31263 THEN
            exp_f := 0;
        ELSIF x =- 31262 THEN
            exp_f := 0;
        ELSIF x =- 31261 THEN
            exp_f := 0;
        ELSIF x =- 31260 THEN
            exp_f := 0;
        ELSIF x =- 31259 THEN
            exp_f := 0;
        ELSIF x =- 31258 THEN
            exp_f := 0;
        ELSIF x =- 31257 THEN
            exp_f := 0;
        ELSIF x =- 31256 THEN
            exp_f := 0;
        ELSIF x =- 31255 THEN
            exp_f := 0;
        ELSIF x =- 31254 THEN
            exp_f := 0;
        ELSIF x =- 31253 THEN
            exp_f := 0;
        ELSIF x =- 31252 THEN
            exp_f := 0;
        ELSIF x =- 31251 THEN
            exp_f := 0;
        ELSIF x =- 31250 THEN
            exp_f := 0;
        ELSIF x =- 31249 THEN
            exp_f := 0;
        ELSIF x =- 31248 THEN
            exp_f := 0;
        ELSIF x =- 31247 THEN
            exp_f := 0;
        ELSIF x =- 31246 THEN
            exp_f := 0;
        ELSIF x =- 31245 THEN
            exp_f := 0;
        ELSIF x =- 31244 THEN
            exp_f := 0;
        ELSIF x =- 31243 THEN
            exp_f := 0;
        ELSIF x =- 31242 THEN
            exp_f := 0;
        ELSIF x =- 31241 THEN
            exp_f := 0;
        ELSIF x =- 31240 THEN
            exp_f := 0;
        ELSIF x =- 31239 THEN
            exp_f := 0;
        ELSIF x =- 31238 THEN
            exp_f := 0;
        ELSIF x =- 31237 THEN
            exp_f := 0;
        ELSIF x =- 31236 THEN
            exp_f := 0;
        ELSIF x =- 31235 THEN
            exp_f := 0;
        ELSIF x =- 31234 THEN
            exp_f := 0;
        ELSIF x =- 31233 THEN
            exp_f := 0;
        ELSIF x =- 31232 THEN
            exp_f := 0;
        ELSIF x =- 31231 THEN
            exp_f := 0;
        ELSIF x =- 31230 THEN
            exp_f := 0;
        ELSIF x =- 31229 THEN
            exp_f := 0;
        ELSIF x =- 31228 THEN
            exp_f := 0;
        ELSIF x =- 31227 THEN
            exp_f := 0;
        ELSIF x =- 31226 THEN
            exp_f := 0;
        ELSIF x =- 31225 THEN
            exp_f := 0;
        ELSIF x =- 31224 THEN
            exp_f := 0;
        ELSIF x =- 31223 THEN
            exp_f := 0;
        ELSIF x =- 31222 THEN
            exp_f := 0;
        ELSIF x =- 31221 THEN
            exp_f := 0;
        ELSIF x =- 31220 THEN
            exp_f := 0;
        ELSIF x =- 31219 THEN
            exp_f := 0;
        ELSIF x =- 31218 THEN
            exp_f := 0;
        ELSIF x =- 31217 THEN
            exp_f := 0;
        ELSIF x =- 31216 THEN
            exp_f := 0;
        ELSIF x =- 31215 THEN
            exp_f := 0;
        ELSIF x =- 31214 THEN
            exp_f := 0;
        ELSIF x =- 31213 THEN
            exp_f := 0;
        ELSIF x =- 31212 THEN
            exp_f := 0;
        ELSIF x =- 31211 THEN
            exp_f := 0;
        ELSIF x =- 31210 THEN
            exp_f := 0;
        ELSIF x =- 31209 THEN
            exp_f := 0;
        ELSIF x =- 31208 THEN
            exp_f := 0;
        ELSIF x =- 31207 THEN
            exp_f := 0;
        ELSIF x =- 31206 THEN
            exp_f := 0;
        ELSIF x =- 31205 THEN
            exp_f := 0;
        ELSIF x =- 31204 THEN
            exp_f := 0;
        ELSIF x =- 31203 THEN
            exp_f := 0;
        ELSIF x =- 31202 THEN
            exp_f := 0;
        ELSIF x =- 31201 THEN
            exp_f := 0;
        ELSIF x =- 31200 THEN
            exp_f := 0;
        ELSIF x =- 31199 THEN
            exp_f := 0;
        ELSIF x =- 31198 THEN
            exp_f := 0;
        ELSIF x =- 31197 THEN
            exp_f := 0;
        ELSIF x =- 31196 THEN
            exp_f := 0;
        ELSIF x =- 31195 THEN
            exp_f := 0;
        ELSIF x =- 31194 THEN
            exp_f := 0;
        ELSIF x =- 31193 THEN
            exp_f := 0;
        ELSIF x =- 31192 THEN
            exp_f := 0;
        ELSIF x =- 31191 THEN
            exp_f := 0;
        ELSIF x =- 31190 THEN
            exp_f := 0;
        ELSIF x =- 31189 THEN
            exp_f := 0;
        ELSIF x =- 31188 THEN
            exp_f := 0;
        ELSIF x =- 31187 THEN
            exp_f := 0;
        ELSIF x =- 31186 THEN
            exp_f := 0;
        ELSIF x =- 31185 THEN
            exp_f := 0;
        ELSIF x =- 31184 THEN
            exp_f := 0;
        ELSIF x =- 31183 THEN
            exp_f := 0;
        ELSIF x =- 31182 THEN
            exp_f := 0;
        ELSIF x =- 31181 THEN
            exp_f := 0;
        ELSIF x =- 31180 THEN
            exp_f := 0;
        ELSIF x =- 31179 THEN
            exp_f := 0;
        ELSIF x =- 31178 THEN
            exp_f := 0;
        ELSIF x =- 31177 THEN
            exp_f := 0;
        ELSIF x =- 31176 THEN
            exp_f := 0;
        ELSIF x =- 31175 THEN
            exp_f := 0;
        ELSIF x =- 31174 THEN
            exp_f := 0;
        ELSIF x =- 31173 THEN
            exp_f := 0;
        ELSIF x =- 31172 THEN
            exp_f := 0;
        ELSIF x =- 31171 THEN
            exp_f := 0;
        ELSIF x =- 31170 THEN
            exp_f := 0;
        ELSIF x =- 31169 THEN
            exp_f := 0;
        ELSIF x =- 31168 THEN
            exp_f := 0;
        ELSIF x =- 31167 THEN
            exp_f := 0;
        ELSIF x =- 31166 THEN
            exp_f := 0;
        ELSIF x =- 31165 THEN
            exp_f := 0;
        ELSIF x =- 31164 THEN
            exp_f := 0;
        ELSIF x =- 31163 THEN
            exp_f := 0;
        ELSIF x =- 31162 THEN
            exp_f := 0;
        ELSIF x =- 31161 THEN
            exp_f := 0;
        ELSIF x =- 31160 THEN
            exp_f := 0;
        ELSIF x =- 31159 THEN
            exp_f := 0;
        ELSIF x =- 31158 THEN
            exp_f := 0;
        ELSIF x =- 31157 THEN
            exp_f := 0;
        ELSIF x =- 31156 THEN
            exp_f := 0;
        ELSIF x =- 31155 THEN
            exp_f := 0;
        ELSIF x =- 31154 THEN
            exp_f := 0;
        ELSIF x =- 31153 THEN
            exp_f := 0;
        ELSIF x =- 31152 THEN
            exp_f := 0;
        ELSIF x =- 31151 THEN
            exp_f := 0;
        ELSIF x =- 31150 THEN
            exp_f := 0;
        ELSIF x =- 31149 THEN
            exp_f := 0;
        ELSIF x =- 31148 THEN
            exp_f := 0;
        ELSIF x =- 31147 THEN
            exp_f := 0;
        ELSIF x =- 31146 THEN
            exp_f := 0;
        ELSIF x =- 31145 THEN
            exp_f := 0;
        ELSIF x =- 31144 THEN
            exp_f := 0;
        ELSIF x =- 31143 THEN
            exp_f := 0;
        ELSIF x =- 31142 THEN
            exp_f := 0;
        ELSIF x =- 31141 THEN
            exp_f := 0;
        ELSIF x =- 31140 THEN
            exp_f := 0;
        ELSIF x =- 31139 THEN
            exp_f := 0;
        ELSIF x =- 31138 THEN
            exp_f := 0;
        ELSIF x =- 31137 THEN
            exp_f := 0;
        ELSIF x =- 31136 THEN
            exp_f := 0;
        ELSIF x =- 31135 THEN
            exp_f := 0;
        ELSIF x =- 31134 THEN
            exp_f := 0;
        ELSIF x =- 31133 THEN
            exp_f := 0;
        ELSIF x =- 31132 THEN
            exp_f := 0;
        ELSIF x =- 31131 THEN
            exp_f := 0;
        ELSIF x =- 31130 THEN
            exp_f := 0;
        ELSIF x =- 31129 THEN
            exp_f := 0;
        ELSIF x =- 31128 THEN
            exp_f := 0;
        ELSIF x =- 31127 THEN
            exp_f := 0;
        ELSIF x =- 31126 THEN
            exp_f := 0;
        ELSIF x =- 31125 THEN
            exp_f := 0;
        ELSIF x =- 31124 THEN
            exp_f := 0;
        ELSIF x =- 31123 THEN
            exp_f := 0;
        ELSIF x =- 31122 THEN
            exp_f := 0;
        ELSIF x =- 31121 THEN
            exp_f := 0;
        ELSIF x =- 31120 THEN
            exp_f := 0;
        ELSIF x =- 31119 THEN
            exp_f := 0;
        ELSIF x =- 31118 THEN
            exp_f := 0;
        ELSIF x =- 31117 THEN
            exp_f := 0;
        ELSIF x =- 31116 THEN
            exp_f := 0;
        ELSIF x =- 31115 THEN
            exp_f := 0;
        ELSIF x =- 31114 THEN
            exp_f := 0;
        ELSIF x =- 31113 THEN
            exp_f := 0;
        ELSIF x =- 31112 THEN
            exp_f := 0;
        ELSIF x =- 31111 THEN
            exp_f := 0;
        ELSIF x =- 31110 THEN
            exp_f := 0;
        ELSIF x =- 31109 THEN
            exp_f := 0;
        ELSIF x =- 31108 THEN
            exp_f := 0;
        ELSIF x =- 31107 THEN
            exp_f := 0;
        ELSIF x =- 31106 THEN
            exp_f := 0;
        ELSIF x =- 31105 THEN
            exp_f := 0;
        ELSIF x =- 31104 THEN
            exp_f := 0;
        ELSIF x =- 31103 THEN
            exp_f := 0;
        ELSIF x =- 31102 THEN
            exp_f := 0;
        ELSIF x =- 31101 THEN
            exp_f := 0;
        ELSIF x =- 31100 THEN
            exp_f := 0;
        ELSIF x =- 31099 THEN
            exp_f := 0;
        ELSIF x =- 31098 THEN
            exp_f := 0;
        ELSIF x =- 31097 THEN
            exp_f := 0;
        ELSIF x =- 31096 THEN
            exp_f := 0;
        ELSIF x =- 31095 THEN
            exp_f := 0;
        ELSIF x =- 31094 THEN
            exp_f := 0;
        ELSIF x =- 31093 THEN
            exp_f := 0;
        ELSIF x =- 31092 THEN
            exp_f := 0;
        ELSIF x =- 31091 THEN
            exp_f := 0;
        ELSIF x =- 31090 THEN
            exp_f := 0;
        ELSIF x =- 31089 THEN
            exp_f := 0;
        ELSIF x =- 31088 THEN
            exp_f := 0;
        ELSIF x =- 31087 THEN
            exp_f := 0;
        ELSIF x =- 31086 THEN
            exp_f := 0;
        ELSIF x =- 31085 THEN
            exp_f := 0;
        ELSIF x =- 31084 THEN
            exp_f := 0;
        ELSIF x =- 31083 THEN
            exp_f := 0;
        ELSIF x =- 31082 THEN
            exp_f := 0;
        ELSIF x =- 31081 THEN
            exp_f := 0;
        ELSIF x =- 31080 THEN
            exp_f := 0;
        ELSIF x =- 31079 THEN
            exp_f := 0;
        ELSIF x =- 31078 THEN
            exp_f := 0;
        ELSIF x =- 31077 THEN
            exp_f := 0;
        ELSIF x =- 31076 THEN
            exp_f := 0;
        ELSIF x =- 31075 THEN
            exp_f := 0;
        ELSIF x =- 31074 THEN
            exp_f := 0;
        ELSIF x =- 31073 THEN
            exp_f := 0;
        ELSIF x =- 31072 THEN
            exp_f := 0;
        ELSIF x =- 31071 THEN
            exp_f := 0;
        ELSIF x =- 31070 THEN
            exp_f := 0;
        ELSIF x =- 31069 THEN
            exp_f := 0;
        ELSIF x =- 31068 THEN
            exp_f := 0;
        ELSIF x =- 31067 THEN
            exp_f := 0;
        ELSIF x =- 31066 THEN
            exp_f := 0;
        ELSIF x =- 31065 THEN
            exp_f := 0;
        ELSIF x =- 31064 THEN
            exp_f := 0;
        ELSIF x =- 31063 THEN
            exp_f := 0;
        ELSIF x =- 31062 THEN
            exp_f := 0;
        ELSIF x =- 31061 THEN
            exp_f := 0;
        ELSIF x =- 31060 THEN
            exp_f := 0;
        ELSIF x =- 31059 THEN
            exp_f := 0;
        ELSIF x =- 31058 THEN
            exp_f := 0;
        ELSIF x =- 31057 THEN
            exp_f := 0;
        ELSIF x =- 31056 THEN
            exp_f := 0;
        ELSIF x =- 31055 THEN
            exp_f := 0;
        ELSIF x =- 31054 THEN
            exp_f := 0;
        ELSIF x =- 31053 THEN
            exp_f := 0;
        ELSIF x =- 31052 THEN
            exp_f := 0;
        ELSIF x =- 31051 THEN
            exp_f := 0;
        ELSIF x =- 31050 THEN
            exp_f := 0;
        ELSIF x =- 31049 THEN
            exp_f := 0;
        ELSIF x =- 31048 THEN
            exp_f := 0;
        ELSIF x =- 31047 THEN
            exp_f := 0;
        ELSIF x =- 31046 THEN
            exp_f := 0;
        ELSIF x =- 31045 THEN
            exp_f := 0;
        ELSIF x =- 31044 THEN
            exp_f := 0;
        ELSIF x =- 31043 THEN
            exp_f := 0;
        ELSIF x =- 31042 THEN
            exp_f := 0;
        ELSIF x =- 31041 THEN
            exp_f := 0;
        ELSIF x =- 31040 THEN
            exp_f := 0;
        ELSIF x =- 31039 THEN
            exp_f := 0;
        ELSIF x =- 31038 THEN
            exp_f := 0;
        ELSIF x =- 31037 THEN
            exp_f := 0;
        ELSIF x =- 31036 THEN
            exp_f := 0;
        ELSIF x =- 31035 THEN
            exp_f := 0;
        ELSIF x =- 31034 THEN
            exp_f := 0;
        ELSIF x =- 31033 THEN
            exp_f := 0;
        ELSIF x =- 31032 THEN
            exp_f := 0;
        ELSIF x =- 31031 THEN
            exp_f := 0;
        ELSIF x =- 31030 THEN
            exp_f := 0;
        ELSIF x =- 31029 THEN
            exp_f := 0;
        ELSIF x =- 31028 THEN
            exp_f := 0;
        ELSIF x =- 31027 THEN
            exp_f := 0;
        ELSIF x =- 31026 THEN
            exp_f := 0;
        ELSIF x =- 31025 THEN
            exp_f := 0;
        ELSIF x =- 31024 THEN
            exp_f := 0;
        ELSIF x =- 31023 THEN
            exp_f := 0;
        ELSIF x =- 31022 THEN
            exp_f := 0;
        ELSIF x =- 31021 THEN
            exp_f := 0;
        ELSIF x =- 31020 THEN
            exp_f := 0;
        ELSIF x =- 31019 THEN
            exp_f := 0;
        ELSIF x =- 31018 THEN
            exp_f := 0;
        ELSIF x =- 31017 THEN
            exp_f := 0;
        ELSIF x =- 31016 THEN
            exp_f := 0;
        ELSIF x =- 31015 THEN
            exp_f := 0;
        ELSIF x =- 31014 THEN
            exp_f := 0;
        ELSIF x =- 31013 THEN
            exp_f := 0;
        ELSIF x =- 31012 THEN
            exp_f := 0;
        ELSIF x =- 31011 THEN
            exp_f := 0;
        ELSIF x =- 31010 THEN
            exp_f := 0;
        ELSIF x =- 31009 THEN
            exp_f := 0;
        ELSIF x =- 31008 THEN
            exp_f := 0;
        ELSIF x =- 31007 THEN
            exp_f := 0;
        ELSIF x =- 31006 THEN
            exp_f := 0;
        ELSIF x =- 31005 THEN
            exp_f := 0;
        ELSIF x =- 31004 THEN
            exp_f := 0;
        ELSIF x =- 31003 THEN
            exp_f := 0;
        ELSIF x =- 31002 THEN
            exp_f := 0;
        ELSIF x =- 31001 THEN
            exp_f := 0;
        ELSIF x =- 31000 THEN
            exp_f := 0;
        ELSIF x =- 30999 THEN
            exp_f := 0;
        ELSIF x =- 30998 THEN
            exp_f := 0;
        ELSIF x =- 30997 THEN
            exp_f := 0;
        ELSIF x =- 30996 THEN
            exp_f := 0;
        ELSIF x =- 30995 THEN
            exp_f := 0;
        ELSIF x =- 30994 THEN
            exp_f := 0;
        ELSIF x =- 30993 THEN
            exp_f := 0;
        ELSIF x =- 30992 THEN
            exp_f := 0;
        ELSIF x =- 30991 THEN
            exp_f := 0;
        ELSIF x =- 30990 THEN
            exp_f := 0;
        ELSIF x =- 30989 THEN
            exp_f := 0;
        ELSIF x =- 30988 THEN
            exp_f := 0;
        ELSIF x =- 30987 THEN
            exp_f := 0;
        ELSIF x =- 30986 THEN
            exp_f := 0;
        ELSIF x =- 30985 THEN
            exp_f := 0;
        ELSIF x =- 30984 THEN
            exp_f := 0;
        ELSIF x =- 30983 THEN
            exp_f := 0;
        ELSIF x =- 30982 THEN
            exp_f := 0;
        ELSIF x =- 30981 THEN
            exp_f := 0;
        ELSIF x =- 30980 THEN
            exp_f := 0;
        ELSIF x =- 30979 THEN
            exp_f := 0;
        ELSIF x =- 30978 THEN
            exp_f := 0;
        ELSIF x =- 30977 THEN
            exp_f := 0;
        ELSIF x =- 30976 THEN
            exp_f := 0;
        ELSIF x =- 30975 THEN
            exp_f := 0;
        ELSIF x =- 30974 THEN
            exp_f := 0;
        ELSIF x =- 30973 THEN
            exp_f := 0;
        ELSIF x =- 30972 THEN
            exp_f := 0;
        ELSIF x =- 30971 THEN
            exp_f := 0;
        ELSIF x =- 30970 THEN
            exp_f := 0;
        ELSIF x =- 30969 THEN
            exp_f := 0;
        ELSIF x =- 30968 THEN
            exp_f := 0;
        ELSIF x =- 30967 THEN
            exp_f := 0;
        ELSIF x =- 30966 THEN
            exp_f := 0;
        ELSIF x =- 30965 THEN
            exp_f := 0;
        ELSIF x =- 30964 THEN
            exp_f := 0;
        ELSIF x =- 30963 THEN
            exp_f := 0;
        ELSIF x =- 30962 THEN
            exp_f := 0;
        ELSIF x =- 30961 THEN
            exp_f := 0;
        ELSIF x =- 30960 THEN
            exp_f := 0;
        ELSIF x =- 30959 THEN
            exp_f := 0;
        ELSIF x =- 30958 THEN
            exp_f := 0;
        ELSIF x =- 30957 THEN
            exp_f := 0;
        ELSIF x =- 30956 THEN
            exp_f := 0;
        ELSIF x =- 30955 THEN
            exp_f := 0;
        ELSIF x =- 30954 THEN
            exp_f := 0;
        ELSIF x =- 30953 THEN
            exp_f := 0;
        ELSIF x =- 30952 THEN
            exp_f := 0;
        ELSIF x =- 30951 THEN
            exp_f := 0;
        ELSIF x =- 30950 THEN
            exp_f := 0;
        ELSIF x =- 30949 THEN
            exp_f := 0;
        ELSIF x =- 30948 THEN
            exp_f := 0;
        ELSIF x =- 30947 THEN
            exp_f := 0;
        ELSIF x =- 30946 THEN
            exp_f := 0;
        ELSIF x =- 30945 THEN
            exp_f := 0;
        ELSIF x =- 30944 THEN
            exp_f := 0;
        ELSIF x =- 30943 THEN
            exp_f := 0;
        ELSIF x =- 30942 THEN
            exp_f := 0;
        ELSIF x =- 30941 THEN
            exp_f := 0;
        ELSIF x =- 30940 THEN
            exp_f := 0;
        ELSIF x =- 30939 THEN
            exp_f := 0;
        ELSIF x =- 30938 THEN
            exp_f := 0;
        ELSIF x =- 30937 THEN
            exp_f := 0;
        ELSIF x =- 30936 THEN
            exp_f := 0;
        ELSIF x =- 30935 THEN
            exp_f := 0;
        ELSIF x =- 30934 THEN
            exp_f := 0;
        ELSIF x =- 30933 THEN
            exp_f := 0;
        ELSIF x =- 30932 THEN
            exp_f := 0;
        ELSIF x =- 30931 THEN
            exp_f := 0;
        ELSIF x =- 30930 THEN
            exp_f := 0;
        ELSIF x =- 30929 THEN
            exp_f := 0;
        ELSIF x =- 30928 THEN
            exp_f := 0;
        ELSIF x =- 30927 THEN
            exp_f := 0;
        ELSIF x =- 30926 THEN
            exp_f := 0;
        ELSIF x =- 30925 THEN
            exp_f := 0;
        ELSIF x =- 30924 THEN
            exp_f := 0;
        ELSIF x =- 30923 THEN
            exp_f := 0;
        ELSIF x =- 30922 THEN
            exp_f := 0;
        ELSIF x =- 30921 THEN
            exp_f := 0;
        ELSIF x =- 30920 THEN
            exp_f := 0;
        ELSIF x =- 30919 THEN
            exp_f := 0;
        ELSIF x =- 30918 THEN
            exp_f := 0;
        ELSIF x =- 30917 THEN
            exp_f := 0;
        ELSIF x =- 30916 THEN
            exp_f := 0;
        ELSIF x =- 30915 THEN
            exp_f := 0;
        ELSIF x =- 30914 THEN
            exp_f := 0;
        ELSIF x =- 30913 THEN
            exp_f := 0;
        ELSIF x =- 30912 THEN
            exp_f := 0;
        ELSIF x =- 30911 THEN
            exp_f := 0;
        ELSIF x =- 30910 THEN
            exp_f := 0;
        ELSIF x =- 30909 THEN
            exp_f := 0;
        ELSIF x =- 30908 THEN
            exp_f := 0;
        ELSIF x =- 30907 THEN
            exp_f := 0;
        ELSIF x =- 30906 THEN
            exp_f := 0;
        ELSIF x =- 30905 THEN
            exp_f := 0;
        ELSIF x =- 30904 THEN
            exp_f := 0;
        ELSIF x =- 30903 THEN
            exp_f := 0;
        ELSIF x =- 30902 THEN
            exp_f := 0;
        ELSIF x =- 30901 THEN
            exp_f := 0;
        ELSIF x =- 30900 THEN
            exp_f := 0;
        ELSIF x =- 30899 THEN
            exp_f := 0;
        ELSIF x =- 30898 THEN
            exp_f := 0;
        ELSIF x =- 30897 THEN
            exp_f := 0;
        ELSIF x =- 30896 THEN
            exp_f := 0;
        ELSIF x =- 30895 THEN
            exp_f := 0;
        ELSIF x =- 30894 THEN
            exp_f := 0;
        ELSIF x =- 30893 THEN
            exp_f := 0;
        ELSIF x =- 30892 THEN
            exp_f := 0;
        ELSIF x =- 30891 THEN
            exp_f := 0;
        ELSIF x =- 30890 THEN
            exp_f := 0;
        ELSIF x =- 30889 THEN
            exp_f := 0;
        ELSIF x =- 30888 THEN
            exp_f := 0;
        ELSIF x =- 30887 THEN
            exp_f := 0;
        ELSIF x =- 30886 THEN
            exp_f := 0;
        ELSIF x =- 30885 THEN
            exp_f := 0;
        ELSIF x =- 30884 THEN
            exp_f := 0;
        ELSIF x =- 30883 THEN
            exp_f := 0;
        ELSIF x =- 30882 THEN
            exp_f := 0;
        ELSIF x =- 30881 THEN
            exp_f := 0;
        ELSIF x =- 30880 THEN
            exp_f := 0;
        ELSIF x =- 30879 THEN
            exp_f := 0;
        ELSIF x =- 30878 THEN
            exp_f := 0;
        ELSIF x =- 30877 THEN
            exp_f := 0;
        ELSIF x =- 30876 THEN
            exp_f := 0;
        ELSIF x =- 30875 THEN
            exp_f := 0;
        ELSIF x =- 30874 THEN
            exp_f := 0;
        ELSIF x =- 30873 THEN
            exp_f := 0;
        ELSIF x =- 30872 THEN
            exp_f := 0;
        ELSIF x =- 30871 THEN
            exp_f := 0;
        ELSIF x =- 30870 THEN
            exp_f := 0;
        ELSIF x =- 30869 THEN
            exp_f := 0;
        ELSIF x =- 30868 THEN
            exp_f := 0;
        ELSIF x =- 30867 THEN
            exp_f := 0;
        ELSIF x =- 30866 THEN
            exp_f := 0;
        ELSIF x =- 30865 THEN
            exp_f := 0;
        ELSIF x =- 30864 THEN
            exp_f := 0;
        ELSIF x =- 30863 THEN
            exp_f := 0;
        ELSIF x =- 30862 THEN
            exp_f := 0;
        ELSIF x =- 30861 THEN
            exp_f := 0;
        ELSIF x =- 30860 THEN
            exp_f := 0;
        ELSIF x =- 30859 THEN
            exp_f := 0;
        ELSIF x =- 30858 THEN
            exp_f := 0;
        ELSIF x =- 30857 THEN
            exp_f := 0;
        ELSIF x =- 30856 THEN
            exp_f := 0;
        ELSIF x =- 30855 THEN
            exp_f := 0;
        ELSIF x =- 30854 THEN
            exp_f := 0;
        ELSIF x =- 30853 THEN
            exp_f := 0;
        ELSIF x =- 30852 THEN
            exp_f := 0;
        ELSIF x =- 30851 THEN
            exp_f := 0;
        ELSIF x =- 30850 THEN
            exp_f := 0;
        ELSIF x =- 30849 THEN
            exp_f := 0;
        ELSIF x =- 30848 THEN
            exp_f := 0;
        ELSIF x =- 30847 THEN
            exp_f := 0;
        ELSIF x =- 30846 THEN
            exp_f := 0;
        ELSIF x =- 30845 THEN
            exp_f := 0;
        ELSIF x =- 30844 THEN
            exp_f := 0;
        ELSIF x =- 30843 THEN
            exp_f := 0;
        ELSIF x =- 30842 THEN
            exp_f := 0;
        ELSIF x =- 30841 THEN
            exp_f := 0;
        ELSIF x =- 30840 THEN
            exp_f := 0;
        ELSIF x =- 30839 THEN
            exp_f := 0;
        ELSIF x =- 30838 THEN
            exp_f := 0;
        ELSIF x =- 30837 THEN
            exp_f := 0;
        ELSIF x =- 30836 THEN
            exp_f := 0;
        ELSIF x =- 30835 THEN
            exp_f := 0;
        ELSIF x =- 30834 THEN
            exp_f := 0;
        ELSIF x =- 30833 THEN
            exp_f := 0;
        ELSIF x =- 30832 THEN
            exp_f := 0;
        ELSIF x =- 30831 THEN
            exp_f := 0;
        ELSIF x =- 30830 THEN
            exp_f := 0;
        ELSIF x =- 30829 THEN
            exp_f := 0;
        ELSIF x =- 30828 THEN
            exp_f := 0;
        ELSIF x =- 30827 THEN
            exp_f := 0;
        ELSIF x =- 30826 THEN
            exp_f := 0;
        ELSIF x =- 30825 THEN
            exp_f := 0;
        ELSIF x =- 30824 THEN
            exp_f := 0;
        ELSIF x =- 30823 THEN
            exp_f := 0;
        ELSIF x =- 30822 THEN
            exp_f := 0;
        ELSIF x =- 30821 THEN
            exp_f := 0;
        ELSIF x =- 30820 THEN
            exp_f := 0;
        ELSIF x =- 30819 THEN
            exp_f := 0;
        ELSIF x =- 30818 THEN
            exp_f := 0;
        ELSIF x =- 30817 THEN
            exp_f := 0;
        ELSIF x =- 30816 THEN
            exp_f := 0;
        ELSIF x =- 30815 THEN
            exp_f := 0;
        ELSIF x =- 30814 THEN
            exp_f := 0;
        ELSIF x =- 30813 THEN
            exp_f := 0;
        ELSIF x =- 30812 THEN
            exp_f := 0;
        ELSIF x =- 30811 THEN
            exp_f := 0;
        ELSIF x =- 30810 THEN
            exp_f := 0;
        ELSIF x =- 30809 THEN
            exp_f := 0;
        ELSIF x =- 30808 THEN
            exp_f := 0;
        ELSIF x =- 30807 THEN
            exp_f := 0;
        ELSIF x =- 30806 THEN
            exp_f := 0;
        ELSIF x =- 30805 THEN
            exp_f := 0;
        ELSIF x =- 30804 THEN
            exp_f := 0;
        ELSIF x =- 30803 THEN
            exp_f := 0;
        ELSIF x =- 30802 THEN
            exp_f := 0;
        ELSIF x =- 30801 THEN
            exp_f := 0;
        ELSIF x =- 30800 THEN
            exp_f := 0;
        ELSIF x =- 30799 THEN
            exp_f := 0;
        ELSIF x =- 30798 THEN
            exp_f := 0;
        ELSIF x =- 30797 THEN
            exp_f := 0;
        ELSIF x =- 30796 THEN
            exp_f := 0;
        ELSIF x =- 30795 THEN
            exp_f := 0;
        ELSIF x =- 30794 THEN
            exp_f := 0;
        ELSIF x =- 30793 THEN
            exp_f := 0;
        ELSIF x =- 30792 THEN
            exp_f := 0;
        ELSIF x =- 30791 THEN
            exp_f := 0;
        ELSIF x =- 30790 THEN
            exp_f := 0;
        ELSIF x =- 30789 THEN
            exp_f := 0;
        ELSIF x =- 30788 THEN
            exp_f := 0;
        ELSIF x =- 30787 THEN
            exp_f := 0;
        ELSIF x =- 30786 THEN
            exp_f := 0;
        ELSIF x =- 30785 THEN
            exp_f := 0;
        ELSIF x =- 30784 THEN
            exp_f := 0;
        ELSIF x =- 30783 THEN
            exp_f := 0;
        ELSIF x =- 30782 THEN
            exp_f := 0;
        ELSIF x =- 30781 THEN
            exp_f := 0;
        ELSIF x =- 30780 THEN
            exp_f := 0;
        ELSIF x =- 30779 THEN
            exp_f := 0;
        ELSIF x =- 30778 THEN
            exp_f := 0;
        ELSIF x =- 30777 THEN
            exp_f := 0;
        ELSIF x =- 30776 THEN
            exp_f := 0;
        ELSIF x =- 30775 THEN
            exp_f := 0;
        ELSIF x =- 30774 THEN
            exp_f := 0;
        ELSIF x =- 30773 THEN
            exp_f := 0;
        ELSIF x =- 30772 THEN
            exp_f := 0;
        ELSIF x =- 30771 THEN
            exp_f := 0;
        ELSIF x =- 30770 THEN
            exp_f := 0;
        ELSIF x =- 30769 THEN
            exp_f := 0;
        ELSIF x =- 30768 THEN
            exp_f := 0;
        ELSIF x =- 30767 THEN
            exp_f := 0;
        ELSIF x =- 30766 THEN
            exp_f := 0;
        ELSIF x =- 30765 THEN
            exp_f := 0;
        ELSIF x =- 30764 THEN
            exp_f := 0;
        ELSIF x =- 30763 THEN
            exp_f := 0;
        ELSIF x =- 30762 THEN
            exp_f := 0;
        ELSIF x =- 30761 THEN
            exp_f := 0;
        ELSIF x =- 30760 THEN
            exp_f := 0;
        ELSIF x =- 30759 THEN
            exp_f := 0;
        ELSIF x =- 30758 THEN
            exp_f := 0;
        ELSIF x =- 30757 THEN
            exp_f := 0;
        ELSIF x =- 30756 THEN
            exp_f := 0;
        ELSIF x =- 30755 THEN
            exp_f := 0;
        ELSIF x =- 30754 THEN
            exp_f := 0;
        ELSIF x =- 30753 THEN
            exp_f := 0;
        ELSIF x =- 30752 THEN
            exp_f := 0;
        ELSIF x =- 30751 THEN
            exp_f := 0;
        ELSIF x =- 30750 THEN
            exp_f := 0;
        ELSIF x =- 30749 THEN
            exp_f := 0;
        ELSIF x =- 30748 THEN
            exp_f := 0;
        ELSIF x =- 30747 THEN
            exp_f := 0;
        ELSIF x =- 30746 THEN
            exp_f := 0;
        ELSIF x =- 30745 THEN
            exp_f := 0;
        ELSIF x =- 30744 THEN
            exp_f := 0;
        ELSIF x =- 30743 THEN
            exp_f := 0;
        ELSIF x =- 30742 THEN
            exp_f := 0;
        ELSIF x =- 30741 THEN
            exp_f := 0;
        ELSIF x =- 30740 THEN
            exp_f := 0;
        ELSIF x =- 30739 THEN
            exp_f := 0;
        ELSIF x =- 30738 THEN
            exp_f := 0;
        ELSIF x =- 30737 THEN
            exp_f := 0;
        ELSIF x =- 30736 THEN
            exp_f := 0;
        ELSIF x =- 30735 THEN
            exp_f := 0;
        ELSIF x =- 30734 THEN
            exp_f := 0;
        ELSIF x =- 30733 THEN
            exp_f := 0;
        ELSIF x =- 30732 THEN
            exp_f := 0;
        ELSIF x =- 30731 THEN
            exp_f := 0;
        ELSIF x =- 30730 THEN
            exp_f := 0;
        ELSIF x =- 30729 THEN
            exp_f := 0;
        ELSIF x =- 30728 THEN
            exp_f := 0;
        ELSIF x =- 30727 THEN
            exp_f := 0;
        ELSIF x =- 30726 THEN
            exp_f := 0;
        ELSIF x =- 30725 THEN
            exp_f := 0;
        ELSIF x =- 30724 THEN
            exp_f := 0;
        ELSIF x =- 30723 THEN
            exp_f := 0;
        ELSIF x =- 30722 THEN
            exp_f := 0;
        ELSIF x =- 30721 THEN
            exp_f := 0;
        ELSIF x =- 30720 THEN
            exp_f := 0;
        ELSIF x =- 30719 THEN
            exp_f := 0;
        ELSIF x =- 30718 THEN
            exp_f := 0;
        ELSIF x =- 30717 THEN
            exp_f := 0;
        ELSIF x =- 30716 THEN
            exp_f := 0;
        ELSIF x =- 30715 THEN
            exp_f := 0;
        ELSIF x =- 30714 THEN
            exp_f := 0;
        ELSIF x =- 30713 THEN
            exp_f := 0;
        ELSIF x =- 30712 THEN
            exp_f := 0;
        ELSIF x =- 30711 THEN
            exp_f := 0;
        ELSIF x =- 30710 THEN
            exp_f := 0;
        ELSIF x =- 30709 THEN
            exp_f := 0;
        ELSIF x =- 30708 THEN
            exp_f := 0;
        ELSIF x =- 30707 THEN
            exp_f := 0;
        ELSIF x =- 30706 THEN
            exp_f := 0;
        ELSIF x =- 30705 THEN
            exp_f := 0;
        ELSIF x =- 30704 THEN
            exp_f := 0;
        ELSIF x =- 30703 THEN
            exp_f := 0;
        ELSIF x =- 30702 THEN
            exp_f := 0;
        ELSIF x =- 30701 THEN
            exp_f := 0;
        ELSIF x =- 30700 THEN
            exp_f := 0;
        ELSIF x =- 30699 THEN
            exp_f := 0;
        ELSIF x =- 30698 THEN
            exp_f := 0;
        ELSIF x =- 30697 THEN
            exp_f := 0;
        ELSIF x =- 30696 THEN
            exp_f := 0;
        ELSIF x =- 30695 THEN
            exp_f := 0;
        ELSIF x =- 30694 THEN
            exp_f := 0;
        ELSIF x =- 30693 THEN
            exp_f := 0;
        ELSIF x =- 30692 THEN
            exp_f := 0;
        ELSIF x =- 30691 THEN
            exp_f := 0;
        ELSIF x =- 30690 THEN
            exp_f := 0;
        ELSIF x =- 30689 THEN
            exp_f := 0;
        ELSIF x =- 30688 THEN
            exp_f := 0;
        ELSIF x =- 30687 THEN
            exp_f := 0;
        ELSIF x =- 30686 THEN
            exp_f := 0;
        ELSIF x =- 30685 THEN
            exp_f := 0;
        ELSIF x =- 30684 THEN
            exp_f := 0;
        ELSIF x =- 30683 THEN
            exp_f := 0;
        ELSIF x =- 30682 THEN
            exp_f := 0;
        ELSIF x =- 30681 THEN
            exp_f := 0;
        ELSIF x =- 30680 THEN
            exp_f := 0;
        ELSIF x =- 30679 THEN
            exp_f := 0;
        ELSIF x =- 30678 THEN
            exp_f := 0;
        ELSIF x =- 30677 THEN
            exp_f := 0;
        ELSIF x =- 30676 THEN
            exp_f := 0;
        ELSIF x =- 30675 THEN
            exp_f := 0;
        ELSIF x =- 30674 THEN
            exp_f := 0;
        ELSIF x =- 30673 THEN
            exp_f := 0;
        ELSIF x =- 30672 THEN
            exp_f := 0;
        ELSIF x =- 30671 THEN
            exp_f := 0;
        ELSIF x =- 30670 THEN
            exp_f := 0;
        ELSIF x =- 30669 THEN
            exp_f := 0;
        ELSIF x =- 30668 THEN
            exp_f := 0;
        ELSIF x =- 30667 THEN
            exp_f := 0;
        ELSIF x =- 30666 THEN
            exp_f := 0;
        ELSIF x =- 30665 THEN
            exp_f := 0;
        ELSIF x =- 30664 THEN
            exp_f := 0;
        ELSIF x =- 30663 THEN
            exp_f := 0;
        ELSIF x =- 30662 THEN
            exp_f := 0;
        ELSIF x =- 30661 THEN
            exp_f := 0;
        ELSIF x =- 30660 THEN
            exp_f := 0;
        ELSIF x =- 30659 THEN
            exp_f := 0;
        ELSIF x =- 30658 THEN
            exp_f := 0;
        ELSIF x =- 30657 THEN
            exp_f := 0;
        ELSIF x =- 30656 THEN
            exp_f := 0;
        ELSIF x =- 30655 THEN
            exp_f := 0;
        ELSIF x =- 30654 THEN
            exp_f := 0;
        ELSIF x =- 30653 THEN
            exp_f := 0;
        ELSIF x =- 30652 THEN
            exp_f := 0;
        ELSIF x =- 30651 THEN
            exp_f := 0;
        ELSIF x =- 30650 THEN
            exp_f := 0;
        ELSIF x =- 30649 THEN
            exp_f := 0;
        ELSIF x =- 30648 THEN
            exp_f := 0;
        ELSIF x =- 30647 THEN
            exp_f := 0;
        ELSIF x =- 30646 THEN
            exp_f := 0;
        ELSIF x =- 30645 THEN
            exp_f := 0;
        ELSIF x =- 30644 THEN
            exp_f := 0;
        ELSIF x =- 30643 THEN
            exp_f := 0;
        ELSIF x =- 30642 THEN
            exp_f := 0;
        ELSIF x =- 30641 THEN
            exp_f := 0;
        ELSIF x =- 30640 THEN
            exp_f := 0;
        ELSIF x =- 30639 THEN
            exp_f := 0;
        ELSIF x =- 30638 THEN
            exp_f := 0;
        ELSIF x =- 30637 THEN
            exp_f := 0;
        ELSIF x =- 30636 THEN
            exp_f := 0;
        ELSIF x =- 30635 THEN
            exp_f := 0;
        ELSIF x =- 30634 THEN
            exp_f := 0;
        ELSIF x =- 30633 THEN
            exp_f := 0;
        ELSIF x =- 30632 THEN
            exp_f := 0;
        ELSIF x =- 30631 THEN
            exp_f := 0;
        ELSIF x =- 30630 THEN
            exp_f := 0;
        ELSIF x =- 30629 THEN
            exp_f := 0;
        ELSIF x =- 30628 THEN
            exp_f := 0;
        ELSIF x =- 30627 THEN
            exp_f := 0;
        ELSIF x =- 30626 THEN
            exp_f := 0;
        ELSIF x =- 30625 THEN
            exp_f := 0;
        ELSIF x =- 30624 THEN
            exp_f := 0;
        ELSIF x =- 30623 THEN
            exp_f := 0;
        ELSIF x =- 30622 THEN
            exp_f := 0;
        ELSIF x =- 30621 THEN
            exp_f := 0;
        ELSIF x =- 30620 THEN
            exp_f := 0;
        ELSIF x =- 30619 THEN
            exp_f := 0;
        ELSIF x =- 30618 THEN
            exp_f := 0;
        ELSIF x =- 30617 THEN
            exp_f := 0;
        ELSIF x =- 30616 THEN
            exp_f := 0;
        ELSIF x =- 30615 THEN
            exp_f := 0;
        ELSIF x =- 30614 THEN
            exp_f := 0;
        ELSIF x =- 30613 THEN
            exp_f := 0;
        ELSIF x =- 30612 THEN
            exp_f := 0;
        ELSIF x =- 30611 THEN
            exp_f := 0;
        ELSIF x =- 30610 THEN
            exp_f := 0;
        ELSIF x =- 30609 THEN
            exp_f := 0;
        ELSIF x =- 30608 THEN
            exp_f := 0;
        ELSIF x =- 30607 THEN
            exp_f := 0;
        ELSIF x =- 30606 THEN
            exp_f := 0;
        ELSIF x =- 30605 THEN
            exp_f := 0;
        ELSIF x =- 30604 THEN
            exp_f := 0;
        ELSIF x =- 30603 THEN
            exp_f := 0;
        ELSIF x =- 30602 THEN
            exp_f := 0;
        ELSIF x =- 30601 THEN
            exp_f := 0;
        ELSIF x =- 30600 THEN
            exp_f := 0;
        ELSIF x =- 30599 THEN
            exp_f := 0;
        ELSIF x =- 30598 THEN
            exp_f := 0;
        ELSIF x =- 30597 THEN
            exp_f := 0;
        ELSIF x =- 30596 THEN
            exp_f := 0;
        ELSIF x =- 30595 THEN
            exp_f := 0;
        ELSIF x =- 30594 THEN
            exp_f := 0;
        ELSIF x =- 30593 THEN
            exp_f := 0;
        ELSIF x =- 30592 THEN
            exp_f := 0;
        ELSIF x =- 30591 THEN
            exp_f := 0;
        ELSIF x =- 30590 THEN
            exp_f := 0;
        ELSIF x =- 30589 THEN
            exp_f := 0;
        ELSIF x =- 30588 THEN
            exp_f := 0;
        ELSIF x =- 30587 THEN
            exp_f := 0;
        ELSIF x =- 30586 THEN
            exp_f := 0;
        ELSIF x =- 30585 THEN
            exp_f := 0;
        ELSIF x =- 30584 THEN
            exp_f := 0;
        ELSIF x =- 30583 THEN
            exp_f := 0;
        ELSIF x =- 30582 THEN
            exp_f := 0;
        ELSIF x =- 30581 THEN
            exp_f := 0;
        ELSIF x =- 30580 THEN
            exp_f := 0;
        ELSIF x =- 30579 THEN
            exp_f := 0;
        ELSIF x =- 30578 THEN
            exp_f := 0;
        ELSIF x =- 30577 THEN
            exp_f := 0;
        ELSIF x =- 30576 THEN
            exp_f := 0;
        ELSIF x =- 30575 THEN
            exp_f := 0;
        ELSIF x =- 30574 THEN
            exp_f := 0;
        ELSIF x =- 30573 THEN
            exp_f := 0;
        ELSIF x =- 30572 THEN
            exp_f := 0;
        ELSIF x =- 30571 THEN
            exp_f := 0;
        ELSIF x =- 30570 THEN
            exp_f := 0;
        ELSIF x =- 30569 THEN
            exp_f := 0;
        ELSIF x =- 30568 THEN
            exp_f := 0;
        ELSIF x =- 30567 THEN
            exp_f := 0;
        ELSIF x =- 30566 THEN
            exp_f := 0;
        ELSIF x =- 30565 THEN
            exp_f := 0;
        ELSIF x =- 30564 THEN
            exp_f := 0;
        ELSIF x =- 30563 THEN
            exp_f := 0;
        ELSIF x =- 30562 THEN
            exp_f := 0;
        ELSIF x =- 30561 THEN
            exp_f := 0;
        ELSIF x =- 30560 THEN
            exp_f := 0;
        ELSIF x =- 30559 THEN
            exp_f := 0;
        ELSIF x =- 30558 THEN
            exp_f := 0;
        ELSIF x =- 30557 THEN
            exp_f := 0;
        ELSIF x =- 30556 THEN
            exp_f := 0;
        ELSIF x =- 30555 THEN
            exp_f := 0;
        ELSIF x =- 30554 THEN
            exp_f := 0;
        ELSIF x =- 30553 THEN
            exp_f := 0;
        ELSIF x =- 30552 THEN
            exp_f := 0;
        ELSIF x =- 30551 THEN
            exp_f := 0;
        ELSIF x =- 30550 THEN
            exp_f := 0;
        ELSIF x =- 30549 THEN
            exp_f := 0;
        ELSIF x =- 30548 THEN
            exp_f := 0;
        ELSIF x =- 30547 THEN
            exp_f := 0;
        ELSIF x =- 30546 THEN
            exp_f := 0;
        ELSIF x =- 30545 THEN
            exp_f := 0;
        ELSIF x =- 30544 THEN
            exp_f := 0;
        ELSIF x =- 30543 THEN
            exp_f := 0;
        ELSIF x =- 30542 THEN
            exp_f := 0;
        ELSIF x =- 30541 THEN
            exp_f := 0;
        ELSIF x =- 30540 THEN
            exp_f := 0;
        ELSIF x =- 30539 THEN
            exp_f := 0;
        ELSIF x =- 30538 THEN
            exp_f := 0;
        ELSIF x =- 30537 THEN
            exp_f := 0;
        ELSIF x =- 30536 THEN
            exp_f := 0;
        ELSIF x =- 30535 THEN
            exp_f := 0;
        ELSIF x =- 30534 THEN
            exp_f := 0;
        ELSIF x =- 30533 THEN
            exp_f := 0;
        ELSIF x =- 30532 THEN
            exp_f := 0;
        ELSIF x =- 30531 THEN
            exp_f := 0;
        ELSIF x =- 30530 THEN
            exp_f := 0;
        ELSIF x =- 30529 THEN
            exp_f := 0;
        ELSIF x =- 30528 THEN
            exp_f := 0;
        ELSIF x =- 30527 THEN
            exp_f := 0;
        ELSIF x =- 30526 THEN
            exp_f := 0;
        ELSIF x =- 30525 THEN
            exp_f := 0;
        ELSIF x =- 30524 THEN
            exp_f := 0;
        ELSIF x =- 30523 THEN
            exp_f := 0;
        ELSIF x =- 30522 THEN
            exp_f := 0;
        ELSIF x =- 30521 THEN
            exp_f := 0;
        ELSIF x =- 30520 THEN
            exp_f := 0;
        ELSIF x =- 30519 THEN
            exp_f := 0;
        ELSIF x =- 30518 THEN
            exp_f := 0;
        ELSIF x =- 30517 THEN
            exp_f := 0;
        ELSIF x =- 30516 THEN
            exp_f := 0;
        ELSIF x =- 30515 THEN
            exp_f := 0;
        ELSIF x =- 30514 THEN
            exp_f := 0;
        ELSIF x =- 30513 THEN
            exp_f := 0;
        ELSIF x =- 30512 THEN
            exp_f := 0;
        ELSIF x =- 30511 THEN
            exp_f := 0;
        ELSIF x =- 30510 THEN
            exp_f := 0;
        ELSIF x =- 30509 THEN
            exp_f := 0;
        ELSIF x =- 30508 THEN
            exp_f := 0;
        ELSIF x =- 30507 THEN
            exp_f := 0;
        ELSIF x =- 30506 THEN
            exp_f := 0;
        ELSIF x =- 30505 THEN
            exp_f := 0;
        ELSIF x =- 30504 THEN
            exp_f := 0;
        ELSIF x =- 30503 THEN
            exp_f := 0;
        ELSIF x =- 30502 THEN
            exp_f := 0;
        ELSIF x =- 30501 THEN
            exp_f := 0;
        ELSIF x =- 30500 THEN
            exp_f := 0;
        ELSIF x =- 30499 THEN
            exp_f := 0;
        ELSIF x =- 30498 THEN
            exp_f := 0;
        ELSIF x =- 30497 THEN
            exp_f := 0;
        ELSIF x =- 30496 THEN
            exp_f := 0;
        ELSIF x =- 30495 THEN
            exp_f := 0;
        ELSIF x =- 30494 THEN
            exp_f := 0;
        ELSIF x =- 30493 THEN
            exp_f := 0;
        ELSIF x =- 30492 THEN
            exp_f := 0;
        ELSIF x =- 30491 THEN
            exp_f := 0;
        ELSIF x =- 30490 THEN
            exp_f := 0;
        ELSIF x =- 30489 THEN
            exp_f := 0;
        ELSIF x =- 30488 THEN
            exp_f := 0;
        ELSIF x =- 30487 THEN
            exp_f := 0;
        ELSIF x =- 30486 THEN
            exp_f := 0;
        ELSIF x =- 30485 THEN
            exp_f := 0;
        ELSIF x =- 30484 THEN
            exp_f := 0;
        ELSIF x =- 30483 THEN
            exp_f := 0;
        ELSIF x =- 30482 THEN
            exp_f := 0;
        ELSIF x =- 30481 THEN
            exp_f := 0;
        ELSIF x =- 30480 THEN
            exp_f := 0;
        ELSIF x =- 30479 THEN
            exp_f := 0;
        ELSIF x =- 30478 THEN
            exp_f := 0;
        ELSIF x =- 30477 THEN
            exp_f := 0;
        ELSIF x =- 30476 THEN
            exp_f := 0;
        ELSIF x =- 30475 THEN
            exp_f := 0;
        ELSIF x =- 30474 THEN
            exp_f := 0;
        ELSIF x =- 30473 THEN
            exp_f := 0;
        ELSIF x =- 30472 THEN
            exp_f := 0;
        ELSIF x =- 30471 THEN
            exp_f := 0;
        ELSIF x =- 30470 THEN
            exp_f := 0;
        ELSIF x =- 30469 THEN
            exp_f := 0;
        ELSIF x =- 30468 THEN
            exp_f := 0;
        ELSIF x =- 30467 THEN
            exp_f := 0;
        ELSIF x =- 30466 THEN
            exp_f := 0;
        ELSIF x =- 30465 THEN
            exp_f := 0;
        ELSIF x =- 30464 THEN
            exp_f := 0;
        ELSIF x =- 30463 THEN
            exp_f := 0;
        ELSIF x =- 30462 THEN
            exp_f := 0;
        ELSIF x =- 30461 THEN
            exp_f := 0;
        ELSIF x =- 30460 THEN
            exp_f := 0;
        ELSIF x =- 30459 THEN
            exp_f := 0;
        ELSIF x =- 30458 THEN
            exp_f := 0;
        ELSIF x =- 30457 THEN
            exp_f := 0;
        ELSIF x =- 30456 THEN
            exp_f := 0;
        ELSIF x =- 30455 THEN
            exp_f := 0;
        ELSIF x =- 30454 THEN
            exp_f := 0;
        ELSIF x =- 30453 THEN
            exp_f := 0;
        ELSIF x =- 30452 THEN
            exp_f := 0;
        ELSIF x =- 30451 THEN
            exp_f := 0;
        ELSIF x =- 30450 THEN
            exp_f := 0;
        ELSIF x =- 30449 THEN
            exp_f := 0;
        ELSIF x =- 30448 THEN
            exp_f := 0;
        ELSIF x =- 30447 THEN
            exp_f := 0;
        ELSIF x =- 30446 THEN
            exp_f := 0;
        ELSIF x =- 30445 THEN
            exp_f := 0;
        ELSIF x =- 30444 THEN
            exp_f := 0;
        ELSIF x =- 30443 THEN
            exp_f := 0;
        ELSIF x =- 30442 THEN
            exp_f := 0;
        ELSIF x =- 30441 THEN
            exp_f := 0;
        ELSIF x =- 30440 THEN
            exp_f := 0;
        ELSIF x =- 30439 THEN
            exp_f := 0;
        ELSIF x =- 30438 THEN
            exp_f := 0;
        ELSIF x =- 30437 THEN
            exp_f := 0;
        ELSIF x =- 30436 THEN
            exp_f := 0;
        ELSIF x =- 30435 THEN
            exp_f := 0;
        ELSIF x =- 30434 THEN
            exp_f := 0;
        ELSIF x =- 30433 THEN
            exp_f := 0;
        ELSIF x =- 30432 THEN
            exp_f := 0;
        ELSIF x =- 30431 THEN
            exp_f := 0;
        ELSIF x =- 30430 THEN
            exp_f := 0;
        ELSIF x =- 30429 THEN
            exp_f := 0;
        ELSIF x =- 30428 THEN
            exp_f := 0;
        ELSIF x =- 30427 THEN
            exp_f := 0;
        ELSIF x =- 30426 THEN
            exp_f := 0;
        ELSIF x =- 30425 THEN
            exp_f := 0;
        ELSIF x =- 30424 THEN
            exp_f := 0;
        ELSIF x =- 30423 THEN
            exp_f := 0;
        ELSIF x =- 30422 THEN
            exp_f := 0;
        ELSIF x =- 30421 THEN
            exp_f := 0;
        ELSIF x =- 30420 THEN
            exp_f := 0;
        ELSIF x =- 30419 THEN
            exp_f := 0;
        ELSIF x =- 30418 THEN
            exp_f := 0;
        ELSIF x =- 30417 THEN
            exp_f := 0;
        ELSIF x =- 30416 THEN
            exp_f := 0;
        ELSIF x =- 30415 THEN
            exp_f := 0;
        ELSIF x =- 30414 THEN
            exp_f := 0;
        ELSIF x =- 30413 THEN
            exp_f := 0;
        ELSIF x =- 30412 THEN
            exp_f := 0;
        ELSIF x =- 30411 THEN
            exp_f := 0;
        ELSIF x =- 30410 THEN
            exp_f := 0;
        ELSIF x =- 30409 THEN
            exp_f := 0;
        ELSIF x =- 30408 THEN
            exp_f := 0;
        ELSIF x =- 30407 THEN
            exp_f := 0;
        ELSIF x =- 30406 THEN
            exp_f := 0;
        ELSIF x =- 30405 THEN
            exp_f := 0;
        ELSIF x =- 30404 THEN
            exp_f := 0;
        ELSIF x =- 30403 THEN
            exp_f := 0;
        ELSIF x =- 30402 THEN
            exp_f := 0;
        ELSIF x =- 30401 THEN
            exp_f := 0;
        ELSIF x =- 30400 THEN
            exp_f := 0;
        ELSIF x =- 30399 THEN
            exp_f := 0;
        ELSIF x =- 30398 THEN
            exp_f := 0;
        ELSIF x =- 30397 THEN
            exp_f := 0;
        ELSIF x =- 30396 THEN
            exp_f := 0;
        ELSIF x =- 30395 THEN
            exp_f := 0;
        ELSIF x =- 30394 THEN
            exp_f := 0;
        ELSIF x =- 30393 THEN
            exp_f := 0;
        ELSIF x =- 30392 THEN
            exp_f := 0;
        ELSIF x =- 30391 THEN
            exp_f := 0;
        ELSIF x =- 30390 THEN
            exp_f := 0;
        ELSIF x =- 30389 THEN
            exp_f := 0;
        ELSIF x =- 30388 THEN
            exp_f := 0;
        ELSIF x =- 30387 THEN
            exp_f := 0;
        ELSIF x =- 30386 THEN
            exp_f := 0;
        ELSIF x =- 30385 THEN
            exp_f := 0;
        ELSIF x =- 30384 THEN
            exp_f := 0;
        ELSIF x =- 30383 THEN
            exp_f := 0;
        ELSIF x =- 30382 THEN
            exp_f := 0;
        ELSIF x =- 30381 THEN
            exp_f := 0;
        ELSIF x =- 30380 THEN
            exp_f := 0;
        ELSIF x =- 30379 THEN
            exp_f := 0;
        ELSIF x =- 30378 THEN
            exp_f := 0;
        ELSIF x =- 30377 THEN
            exp_f := 0;
        ELSIF x =- 30376 THEN
            exp_f := 0;
        ELSIF x =- 30375 THEN
            exp_f := 0;
        ELSIF x =- 30374 THEN
            exp_f := 0;
        ELSIF x =- 30373 THEN
            exp_f := 0;
        ELSIF x =- 30372 THEN
            exp_f := 0;
        ELSIF x =- 30371 THEN
            exp_f := 0;
        ELSIF x =- 30370 THEN
            exp_f := 0;
        ELSIF x =- 30369 THEN
            exp_f := 0;
        ELSIF x =- 30368 THEN
            exp_f := 0;
        ELSIF x =- 30367 THEN
            exp_f := 0;
        ELSIF x =- 30366 THEN
            exp_f := 0;
        ELSIF x =- 30365 THEN
            exp_f := 0;
        ELSIF x =- 30364 THEN
            exp_f := 0;
        ELSIF x =- 30363 THEN
            exp_f := 0;
        ELSIF x =- 30362 THEN
            exp_f := 0;
        ELSIF x =- 30361 THEN
            exp_f := 0;
        ELSIF x =- 30360 THEN
            exp_f := 0;
        ELSIF x =- 30359 THEN
            exp_f := 0;
        ELSIF x =- 30358 THEN
            exp_f := 0;
        ELSIF x =- 30357 THEN
            exp_f := 0;
        ELSIF x =- 30356 THEN
            exp_f := 0;
        ELSIF x =- 30355 THEN
            exp_f := 0;
        ELSIF x =- 30354 THEN
            exp_f := 0;
        ELSIF x =- 30353 THEN
            exp_f := 0;
        ELSIF x =- 30352 THEN
            exp_f := 0;
        ELSIF x =- 30351 THEN
            exp_f := 0;
        ELSIF x =- 30350 THEN
            exp_f := 0;
        ELSIF x =- 30349 THEN
            exp_f := 0;
        ELSIF x =- 30348 THEN
            exp_f := 0;
        ELSIF x =- 30347 THEN
            exp_f := 0;
        ELSIF x =- 30346 THEN
            exp_f := 0;
        ELSIF x =- 30345 THEN
            exp_f := 0;
        ELSIF x =- 30344 THEN
            exp_f := 0;
        ELSIF x =- 30343 THEN
            exp_f := 0;
        ELSIF x =- 30342 THEN
            exp_f := 0;
        ELSIF x =- 30341 THEN
            exp_f := 0;
        ELSIF x =- 30340 THEN
            exp_f := 0;
        ELSIF x =- 30339 THEN
            exp_f := 0;
        ELSIF x =- 30338 THEN
            exp_f := 0;
        ELSIF x =- 30337 THEN
            exp_f := 0;
        ELSIF x =- 30336 THEN
            exp_f := 0;
        ELSIF x =- 30335 THEN
            exp_f := 0;
        ELSIF x =- 30334 THEN
            exp_f := 0;
        ELSIF x =- 30333 THEN
            exp_f := 0;
        ELSIF x =- 30332 THEN
            exp_f := 0;
        ELSIF x =- 30331 THEN
            exp_f := 0;
        ELSIF x =- 30330 THEN
            exp_f := 0;
        ELSIF x =- 30329 THEN
            exp_f := 0;
        ELSIF x =- 30328 THEN
            exp_f := 0;
        ELSIF x =- 30327 THEN
            exp_f := 0;
        ELSIF x =- 30326 THEN
            exp_f := 0;
        ELSIF x =- 30325 THEN
            exp_f := 0;
        ELSIF x =- 30324 THEN
            exp_f := 0;
        ELSIF x =- 30323 THEN
            exp_f := 0;
        ELSIF x =- 30322 THEN
            exp_f := 0;
        ELSIF x =- 30321 THEN
            exp_f := 0;
        ELSIF x =- 30320 THEN
            exp_f := 0;
        ELSIF x =- 30319 THEN
            exp_f := 0;
        ELSIF x =- 30318 THEN
            exp_f := 0;
        ELSIF x =- 30317 THEN
            exp_f := 0;
        ELSIF x =- 30316 THEN
            exp_f := 0;
        ELSIF x =- 30315 THEN
            exp_f := 0;
        ELSIF x =- 30314 THEN
            exp_f := 0;
        ELSIF x =- 30313 THEN
            exp_f := 0;
        ELSIF x =- 30312 THEN
            exp_f := 0;
        ELSIF x =- 30311 THEN
            exp_f := 0;
        ELSIF x =- 30310 THEN
            exp_f := 0;
        ELSIF x =- 30309 THEN
            exp_f := 0;
        ELSIF x =- 30308 THEN
            exp_f := 0;
        ELSIF x =- 30307 THEN
            exp_f := 0;
        ELSIF x =- 30306 THEN
            exp_f := 0;
        ELSIF x =- 30305 THEN
            exp_f := 0;
        ELSIF x =- 30304 THEN
            exp_f := 0;
        ELSIF x =- 30303 THEN
            exp_f := 0;
        ELSIF x =- 30302 THEN
            exp_f := 0;
        ELSIF x =- 30301 THEN
            exp_f := 0;
        ELSIF x =- 30300 THEN
            exp_f := 0;
        ELSIF x =- 30299 THEN
            exp_f := 0;
        ELSIF x =- 30298 THEN
            exp_f := 0;
        ELSIF x =- 30297 THEN
            exp_f := 0;
        ELSIF x =- 30296 THEN
            exp_f := 0;
        ELSIF x =- 30295 THEN
            exp_f := 0;
        ELSIF x =- 30294 THEN
            exp_f := 0;
        ELSIF x =- 30293 THEN
            exp_f := 0;
        ELSIF x =- 30292 THEN
            exp_f := 0;
        ELSIF x =- 30291 THEN
            exp_f := 0;
        ELSIF x =- 30290 THEN
            exp_f := 0;
        ELSIF x =- 30289 THEN
            exp_f := 0;
        ELSIF x =- 30288 THEN
            exp_f := 0;
        ELSIF x =- 30287 THEN
            exp_f := 0;
        ELSIF x =- 30286 THEN
            exp_f := 0;
        ELSIF x =- 30285 THEN
            exp_f := 0;
        ELSIF x =- 30284 THEN
            exp_f := 0;
        ELSIF x =- 30283 THEN
            exp_f := 0;
        ELSIF x =- 30282 THEN
            exp_f := 0;
        ELSIF x =- 30281 THEN
            exp_f := 0;
        ELSIF x =- 30280 THEN
            exp_f := 0;
        ELSIF x =- 30279 THEN
            exp_f := 0;
        ELSIF x =- 30278 THEN
            exp_f := 0;
        ELSIF x =- 30277 THEN
            exp_f := 0;
        ELSIF x =- 30276 THEN
            exp_f := 0;
        ELSIF x =- 30275 THEN
            exp_f := 0;
        ELSIF x =- 30274 THEN
            exp_f := 0;
        ELSIF x =- 30273 THEN
            exp_f := 0;
        ELSIF x =- 30272 THEN
            exp_f := 0;
        ELSIF x =- 30271 THEN
            exp_f := 0;
        ELSIF x =- 30270 THEN
            exp_f := 0;
        ELSIF x =- 30269 THEN
            exp_f := 0;
        ELSIF x =- 30268 THEN
            exp_f := 0;
        ELSIF x =- 30267 THEN
            exp_f := 0;
        ELSIF x =- 30266 THEN
            exp_f := 0;
        ELSIF x =- 30265 THEN
            exp_f := 0;
        ELSIF x =- 30264 THEN
            exp_f := 0;
        ELSIF x =- 30263 THEN
            exp_f := 0;
        ELSIF x =- 30262 THEN
            exp_f := 0;
        ELSIF x =- 30261 THEN
            exp_f := 0;
        ELSIF x =- 30260 THEN
            exp_f := 0;
        ELSIF x =- 30259 THEN
            exp_f := 0;
        ELSIF x =- 30258 THEN
            exp_f := 0;
        ELSIF x =- 30257 THEN
            exp_f := 0;
        ELSIF x =- 30256 THEN
            exp_f := 0;
        ELSIF x =- 30255 THEN
            exp_f := 0;
        ELSIF x =- 30254 THEN
            exp_f := 0;
        ELSIF x =- 30253 THEN
            exp_f := 0;
        ELSIF x =- 30252 THEN
            exp_f := 0;
        ELSIF x =- 30251 THEN
            exp_f := 0;
        ELSIF x =- 30250 THEN
            exp_f := 0;
        ELSIF x =- 30249 THEN
            exp_f := 0;
        ELSIF x =- 30248 THEN
            exp_f := 0;
        ELSIF x =- 30247 THEN
            exp_f := 0;
        ELSIF x =- 30246 THEN
            exp_f := 0;
        ELSIF x =- 30245 THEN
            exp_f := 0;
        ELSIF x =- 30244 THEN
            exp_f := 0;
        ELSIF x =- 30243 THEN
            exp_f := 0;
        ELSIF x =- 30242 THEN
            exp_f := 0;
        ELSIF x =- 30241 THEN
            exp_f := 0;
        ELSIF x =- 30240 THEN
            exp_f := 0;
        ELSIF x =- 30239 THEN
            exp_f := 0;
        ELSIF x =- 30238 THEN
            exp_f := 0;
        ELSIF x =- 30237 THEN
            exp_f := 0;
        ELSIF x =- 30236 THEN
            exp_f := 0;
        ELSIF x =- 30235 THEN
            exp_f := 0;
        ELSIF x =- 30234 THEN
            exp_f := 0;
        ELSIF x =- 30233 THEN
            exp_f := 0;
        ELSIF x =- 30232 THEN
            exp_f := 0;
        ELSIF x =- 30231 THEN
            exp_f := 0;
        ELSIF x =- 30230 THEN
            exp_f := 0;
        ELSIF x =- 30229 THEN
            exp_f := 0;
        ELSIF x =- 30228 THEN
            exp_f := 0;
        ELSIF x =- 30227 THEN
            exp_f := 0;
        ELSIF x =- 30226 THEN
            exp_f := 0;
        ELSIF x =- 30225 THEN
            exp_f := 0;
        ELSIF x =- 30224 THEN
            exp_f := 0;
        ELSIF x =- 30223 THEN
            exp_f := 0;
        ELSIF x =- 30222 THEN
            exp_f := 0;
        ELSIF x =- 30221 THEN
            exp_f := 0;
        ELSIF x =- 30220 THEN
            exp_f := 0;
        ELSIF x =- 30219 THEN
            exp_f := 0;
        ELSIF x =- 30218 THEN
            exp_f := 0;
        ELSIF x =- 30217 THEN
            exp_f := 0;
        ELSIF x =- 30216 THEN
            exp_f := 0;
        ELSIF x =- 30215 THEN
            exp_f := 0;
        ELSIF x =- 30214 THEN
            exp_f := 0;
        ELSIF x =- 30213 THEN
            exp_f := 0;
        ELSIF x =- 30212 THEN
            exp_f := 0;
        ELSIF x =- 30211 THEN
            exp_f := 0;
        ELSIF x =- 30210 THEN
            exp_f := 0;
        ELSIF x =- 30209 THEN
            exp_f := 0;
        ELSIF x =- 30208 THEN
            exp_f := 0;
        ELSIF x =- 30207 THEN
            exp_f := 0;
        ELSIF x =- 30206 THEN
            exp_f := 0;
        ELSIF x =- 30205 THEN
            exp_f := 0;
        ELSIF x =- 30204 THEN
            exp_f := 0;
        ELSIF x =- 30203 THEN
            exp_f := 0;
        ELSIF x =- 30202 THEN
            exp_f := 0;
        ELSIF x =- 30201 THEN
            exp_f := 0;
        ELSIF x =- 30200 THEN
            exp_f := 0;
        ELSIF x =- 30199 THEN
            exp_f := 0;
        ELSIF x =- 30198 THEN
            exp_f := 0;
        ELSIF x =- 30197 THEN
            exp_f := 0;
        ELSIF x =- 30196 THEN
            exp_f := 0;
        ELSIF x =- 30195 THEN
            exp_f := 0;
        ELSIF x =- 30194 THEN
            exp_f := 0;
        ELSIF x =- 30193 THEN
            exp_f := 0;
        ELSIF x =- 30192 THEN
            exp_f := 0;
        ELSIF x =- 30191 THEN
            exp_f := 0;
        ELSIF x =- 30190 THEN
            exp_f := 0;
        ELSIF x =- 30189 THEN
            exp_f := 0;
        ELSIF x =- 30188 THEN
            exp_f := 0;
        ELSIF x =- 30187 THEN
            exp_f := 0;
        ELSIF x =- 30186 THEN
            exp_f := 0;
        ELSIF x =- 30185 THEN
            exp_f := 0;
        ELSIF x =- 30184 THEN
            exp_f := 0;
        ELSIF x =- 30183 THEN
            exp_f := 0;
        ELSIF x =- 30182 THEN
            exp_f := 0;
        ELSIF x =- 30181 THEN
            exp_f := 0;
        ELSIF x =- 30180 THEN
            exp_f := 0;
        ELSIF x =- 30179 THEN
            exp_f := 0;
        ELSIF x =- 30178 THEN
            exp_f := 0;
        ELSIF x =- 30177 THEN
            exp_f := 0;
        ELSIF x =- 30176 THEN
            exp_f := 0;
        ELSIF x =- 30175 THEN
            exp_f := 0;
        ELSIF x =- 30174 THEN
            exp_f := 0;
        ELSIF x =- 30173 THEN
            exp_f := 0;
        ELSIF x =- 30172 THEN
            exp_f := 0;
        ELSIF x =- 30171 THEN
            exp_f := 0;
        ELSIF x =- 30170 THEN
            exp_f := 0;
        ELSIF x =- 30169 THEN
            exp_f := 0;
        ELSIF x =- 30168 THEN
            exp_f := 0;
        ELSIF x =- 30167 THEN
            exp_f := 0;
        ELSIF x =- 30166 THEN
            exp_f := 0;
        ELSIF x =- 30165 THEN
            exp_f := 0;
        ELSIF x =- 30164 THEN
            exp_f := 0;
        ELSIF x =- 30163 THEN
            exp_f := 0;
        ELSIF x =- 30162 THEN
            exp_f := 0;
        ELSIF x =- 30161 THEN
            exp_f := 0;
        ELSIF x =- 30160 THEN
            exp_f := 0;
        ELSIF x =- 30159 THEN
            exp_f := 0;
        ELSIF x =- 30158 THEN
            exp_f := 0;
        ELSIF x =- 30157 THEN
            exp_f := 0;
        ELSIF x =- 30156 THEN
            exp_f := 0;
        ELSIF x =- 30155 THEN
            exp_f := 0;
        ELSIF x =- 30154 THEN
            exp_f := 0;
        ELSIF x =- 30153 THEN
            exp_f := 0;
        ELSIF x =- 30152 THEN
            exp_f := 0;
        ELSIF x =- 30151 THEN
            exp_f := 0;
        ELSIF x =- 30150 THEN
            exp_f := 0;
        ELSIF x =- 30149 THEN
            exp_f := 0;
        ELSIF x =- 30148 THEN
            exp_f := 0;
        ELSIF x =- 30147 THEN
            exp_f := 0;
        ELSIF x =- 30146 THEN
            exp_f := 0;
        ELSIF x =- 30145 THEN
            exp_f := 0;
        ELSIF x =- 30144 THEN
            exp_f := 0;
        ELSIF x =- 30143 THEN
            exp_f := 0;
        ELSIF x =- 30142 THEN
            exp_f := 0;
        ELSIF x =- 30141 THEN
            exp_f := 0;
        ELSIF x =- 30140 THEN
            exp_f := 0;
        ELSIF x =- 30139 THEN
            exp_f := 0;
        ELSIF x =- 30138 THEN
            exp_f := 0;
        ELSIF x =- 30137 THEN
            exp_f := 0;
        ELSIF x =- 30136 THEN
            exp_f := 0;
        ELSIF x =- 30135 THEN
            exp_f := 0;
        ELSIF x =- 30134 THEN
            exp_f := 0;
        ELSIF x =- 30133 THEN
            exp_f := 0;
        ELSIF x =- 30132 THEN
            exp_f := 0;
        ELSIF x =- 30131 THEN
            exp_f := 0;
        ELSIF x =- 30130 THEN
            exp_f := 0;
        ELSIF x =- 30129 THEN
            exp_f := 0;
        ELSIF x =- 30128 THEN
            exp_f := 0;
        ELSIF x =- 30127 THEN
            exp_f := 0;
        ELSIF x =- 30126 THEN
            exp_f := 0;
        ELSIF x =- 30125 THEN
            exp_f := 0;
        ELSIF x =- 30124 THEN
            exp_f := 0;
        ELSIF x =- 30123 THEN
            exp_f := 0;
        ELSIF x =- 30122 THEN
            exp_f := 0;
        ELSIF x =- 30121 THEN
            exp_f := 0;
        ELSIF x =- 30120 THEN
            exp_f := 0;
        ELSIF x =- 30119 THEN
            exp_f := 0;
        ELSIF x =- 30118 THEN
            exp_f := 0;
        ELSIF x =- 30117 THEN
            exp_f := 0;
        ELSIF x =- 30116 THEN
            exp_f := 0;
        ELSIF x =- 30115 THEN
            exp_f := 0;
        ELSIF x =- 30114 THEN
            exp_f := 0;
        ELSIF x =- 30113 THEN
            exp_f := 0;
        ELSIF x =- 30112 THEN
            exp_f := 0;
        ELSIF x =- 30111 THEN
            exp_f := 0;
        ELSIF x =- 30110 THEN
            exp_f := 0;
        ELSIF x =- 30109 THEN
            exp_f := 0;
        ELSIF x =- 30108 THEN
            exp_f := 0;
        ELSIF x =- 30107 THEN
            exp_f := 0;
        ELSIF x =- 30106 THEN
            exp_f := 0;
        ELSIF x =- 30105 THEN
            exp_f := 0;
        ELSIF x =- 30104 THEN
            exp_f := 0;
        ELSIF x =- 30103 THEN
            exp_f := 0;
        ELSIF x =- 30102 THEN
            exp_f := 0;
        ELSIF x =- 30101 THEN
            exp_f := 0;
        ELSIF x =- 30100 THEN
            exp_f := 0;
        ELSIF x =- 30099 THEN
            exp_f := 0;
        ELSIF x =- 30098 THEN
            exp_f := 0;
        ELSIF x =- 30097 THEN
            exp_f := 0;
        ELSIF x =- 30096 THEN
            exp_f := 0;
        ELSIF x =- 30095 THEN
            exp_f := 0;
        ELSIF x =- 30094 THEN
            exp_f := 0;
        ELSIF x =- 30093 THEN
            exp_f := 0;
        ELSIF x =- 30092 THEN
            exp_f := 0;
        ELSIF x =- 30091 THEN
            exp_f := 0;
        ELSIF x =- 30090 THEN
            exp_f := 0;
        ELSIF x =- 30089 THEN
            exp_f := 0;
        ELSIF x =- 30088 THEN
            exp_f := 0;
        ELSIF x =- 30087 THEN
            exp_f := 0;
        ELSIF x =- 30086 THEN
            exp_f := 0;
        ELSIF x =- 30085 THEN
            exp_f := 0;
        ELSIF x =- 30084 THEN
            exp_f := 0;
        ELSIF x =- 30083 THEN
            exp_f := 0;
        ELSIF x =- 30082 THEN
            exp_f := 0;
        ELSIF x =- 30081 THEN
            exp_f := 0;
        ELSIF x =- 30080 THEN
            exp_f := 0;
        ELSIF x =- 30079 THEN
            exp_f := 0;
        ELSIF x =- 30078 THEN
            exp_f := 0;
        ELSIF x =- 30077 THEN
            exp_f := 0;
        ELSIF x =- 30076 THEN
            exp_f := 0;
        ELSIF x =- 30075 THEN
            exp_f := 0;
        ELSIF x =- 30074 THEN
            exp_f := 0;
        ELSIF x =- 30073 THEN
            exp_f := 0;
        ELSIF x =- 30072 THEN
            exp_f := 0;
        ELSIF x =- 30071 THEN
            exp_f := 0;
        ELSIF x =- 30070 THEN
            exp_f := 0;
        ELSIF x =- 30069 THEN
            exp_f := 0;
        ELSIF x =- 30068 THEN
            exp_f := 0;
        ELSIF x =- 30067 THEN
            exp_f := 0;
        ELSIF x =- 30066 THEN
            exp_f := 0;
        ELSIF x =- 30065 THEN
            exp_f := 0;
        ELSIF x =- 30064 THEN
            exp_f := 0;
        ELSIF x =- 30063 THEN
            exp_f := 0;
        ELSIF x =- 30062 THEN
            exp_f := 0;
        ELSIF x =- 30061 THEN
            exp_f := 0;
        ELSIF x =- 30060 THEN
            exp_f := 0;
        ELSIF x =- 30059 THEN
            exp_f := 0;
        ELSIF x =- 30058 THEN
            exp_f := 0;
        ELSIF x =- 30057 THEN
            exp_f := 0;
        ELSIF x =- 30056 THEN
            exp_f := 0;
        ELSIF x =- 30055 THEN
            exp_f := 0;
        ELSIF x =- 30054 THEN
            exp_f := 0;
        ELSIF x =- 30053 THEN
            exp_f := 0;
        ELSIF x =- 30052 THEN
            exp_f := 0;
        ELSIF x =- 30051 THEN
            exp_f := 0;
        ELSIF x =- 30050 THEN
            exp_f := 0;
        ELSIF x =- 30049 THEN
            exp_f := 0;
        ELSIF x =- 30048 THEN
            exp_f := 0;
        ELSIF x =- 30047 THEN
            exp_f := 0;
        ELSIF x =- 30046 THEN
            exp_f := 0;
        ELSIF x =- 30045 THEN
            exp_f := 0;
        ELSIF x =- 30044 THEN
            exp_f := 0;
        ELSIF x =- 30043 THEN
            exp_f := 0;
        ELSIF x =- 30042 THEN
            exp_f := 0;
        ELSIF x =- 30041 THEN
            exp_f := 0;
        ELSIF x =- 30040 THEN
            exp_f := 0;
        ELSIF x =- 30039 THEN
            exp_f := 0;
        ELSIF x =- 30038 THEN
            exp_f := 0;
        ELSIF x =- 30037 THEN
            exp_f := 0;
        ELSIF x =- 30036 THEN
            exp_f := 0;
        ELSIF x =- 30035 THEN
            exp_f := 0;
        ELSIF x =- 30034 THEN
            exp_f := 0;
        ELSIF x =- 30033 THEN
            exp_f := 0;
        ELSIF x =- 30032 THEN
            exp_f := 0;
        ELSIF x =- 30031 THEN
            exp_f := 0;
        ELSIF x =- 30030 THEN
            exp_f := 0;
        ELSIF x =- 30029 THEN
            exp_f := 0;
        ELSIF x =- 30028 THEN
            exp_f := 0;
        ELSIF x =- 30027 THEN
            exp_f := 0;
        ELSIF x =- 30026 THEN
            exp_f := 0;
        ELSIF x =- 30025 THEN
            exp_f := 0;
        ELSIF x =- 30024 THEN
            exp_f := 0;
        ELSIF x =- 30023 THEN
            exp_f := 0;
        ELSIF x =- 30022 THEN
            exp_f := 0;
        ELSIF x =- 30021 THEN
            exp_f := 0;
        ELSIF x =- 30020 THEN
            exp_f := 0;
        ELSIF x =- 30019 THEN
            exp_f := 0;
        ELSIF x =- 30018 THEN
            exp_f := 0;
        ELSIF x =- 30017 THEN
            exp_f := 0;
        ELSIF x =- 30016 THEN
            exp_f := 0;
        ELSIF x =- 30015 THEN
            exp_f := 0;
        ELSIF x =- 30014 THEN
            exp_f := 0;
        ELSIF x =- 30013 THEN
            exp_f := 0;
        ELSIF x =- 30012 THEN
            exp_f := 0;
        ELSIF x =- 30011 THEN
            exp_f := 0;
        ELSIF x =- 30010 THEN
            exp_f := 0;
        ELSIF x =- 30009 THEN
            exp_f := 0;
        ELSIF x =- 30008 THEN
            exp_f := 0;
        ELSIF x =- 30007 THEN
            exp_f := 0;
        ELSIF x =- 30006 THEN
            exp_f := 0;
        ELSIF x =- 30005 THEN
            exp_f := 0;
        ELSIF x =- 30004 THEN
            exp_f := 0;
        ELSIF x =- 30003 THEN
            exp_f := 0;
        ELSIF x =- 30002 THEN
            exp_f := 0;
        ELSIF x =- 30001 THEN
            exp_f := 0;
        ELSIF x =- 30000 THEN
            exp_f := 0;
        ELSIF x =- 29999 THEN
            exp_f := 0;
        ELSIF x =- 29998 THEN
            exp_f := 0;
        ELSIF x =- 29997 THEN
            exp_f := 0;
        ELSIF x =- 29996 THEN
            exp_f := 0;
        ELSIF x =- 29995 THEN
            exp_f := 0;
        ELSIF x =- 29994 THEN
            exp_f := 0;
        ELSIF x =- 29993 THEN
            exp_f := 0;
        ELSIF x =- 29992 THEN
            exp_f := 0;
        ELSIF x =- 29991 THEN
            exp_f := 0;
        ELSIF x =- 29990 THEN
            exp_f := 0;
        ELSIF x =- 29989 THEN
            exp_f := 0;
        ELSIF x =- 29988 THEN
            exp_f := 0;
        ELSIF x =- 29987 THEN
            exp_f := 0;
        ELSIF x =- 29986 THEN
            exp_f := 0;
        ELSIF x =- 29985 THEN
            exp_f := 0;
        ELSIF x =- 29984 THEN
            exp_f := 0;
        ELSIF x =- 29983 THEN
            exp_f := 0;
        ELSIF x =- 29982 THEN
            exp_f := 0;
        ELSIF x =- 29981 THEN
            exp_f := 0;
        ELSIF x =- 29980 THEN
            exp_f := 0;
        ELSIF x =- 29979 THEN
            exp_f := 0;
        ELSIF x =- 29978 THEN
            exp_f := 0;
        ELSIF x =- 29977 THEN
            exp_f := 0;
        ELSIF x =- 29976 THEN
            exp_f := 0;
        ELSIF x =- 29975 THEN
            exp_f := 0;
        ELSIF x =- 29974 THEN
            exp_f := 0;
        ELSIF x =- 29973 THEN
            exp_f := 0;
        ELSIF x =- 29972 THEN
            exp_f := 0;
        ELSIF x =- 29971 THEN
            exp_f := 0;
        ELSIF x =- 29970 THEN
            exp_f := 0;
        ELSIF x =- 29969 THEN
            exp_f := 0;
        ELSIF x =- 29968 THEN
            exp_f := 0;
        ELSIF x =- 29967 THEN
            exp_f := 0;
        ELSIF x =- 29966 THEN
            exp_f := 0;
        ELSIF x =- 29965 THEN
            exp_f := 0;
        ELSIF x =- 29964 THEN
            exp_f := 0;
        ELSIF x =- 29963 THEN
            exp_f := 0;
        ELSIF x =- 29962 THEN
            exp_f := 0;
        ELSIF x =- 29961 THEN
            exp_f := 0;
        ELSIF x =- 29960 THEN
            exp_f := 0;
        ELSIF x =- 29959 THEN
            exp_f := 0;
        ELSIF x =- 29958 THEN
            exp_f := 0;
        ELSIF x =- 29957 THEN
            exp_f := 0;
        ELSIF x =- 29956 THEN
            exp_f := 0;
        ELSIF x =- 29955 THEN
            exp_f := 0;
        ELSIF x =- 29954 THEN
            exp_f := 0;
        ELSIF x =- 29953 THEN
            exp_f := 0;
        ELSIF x =- 29952 THEN
            exp_f := 0;
        ELSIF x =- 29951 THEN
            exp_f := 0;
        ELSIF x =- 29950 THEN
            exp_f := 0;
        ELSIF x =- 29949 THEN
            exp_f := 0;
        ELSIF x =- 29948 THEN
            exp_f := 0;
        ELSIF x =- 29947 THEN
            exp_f := 0;
        ELSIF x =- 29946 THEN
            exp_f := 0;
        ELSIF x =- 29945 THEN
            exp_f := 0;
        ELSIF x =- 29944 THEN
            exp_f := 0;
        ELSIF x =- 29943 THEN
            exp_f := 0;
        ELSIF x =- 29942 THEN
            exp_f := 0;
        ELSIF x =- 29941 THEN
            exp_f := 0;
        ELSIF x =- 29940 THEN
            exp_f := 0;
        ELSIF x =- 29939 THEN
            exp_f := 0;
        ELSIF x =- 29938 THEN
            exp_f := 0;
        ELSIF x =- 29937 THEN
            exp_f := 0;
        ELSIF x =- 29936 THEN
            exp_f := 0;
        ELSIF x =- 29935 THEN
            exp_f := 0;
        ELSIF x =- 29934 THEN
            exp_f := 0;
        ELSIF x =- 29933 THEN
            exp_f := 0;
        ELSIF x =- 29932 THEN
            exp_f := 0;
        ELSIF x =- 29931 THEN
            exp_f := 0;
        ELSIF x =- 29930 THEN
            exp_f := 0;
        ELSIF x =- 29929 THEN
            exp_f := 0;
        ELSIF x =- 29928 THEN
            exp_f := 0;
        ELSIF x =- 29927 THEN
            exp_f := 0;
        ELSIF x =- 29926 THEN
            exp_f := 0;
        ELSIF x =- 29925 THEN
            exp_f := 0;
        ELSIF x =- 29924 THEN
            exp_f := 0;
        ELSIF x =- 29923 THEN
            exp_f := 0;
        ELSIF x =- 29922 THEN
            exp_f := 0;
        ELSIF x =- 29921 THEN
            exp_f := 0;
        ELSIF x =- 29920 THEN
            exp_f := 0;
        ELSIF x =- 29919 THEN
            exp_f := 0;
        ELSIF x =- 29918 THEN
            exp_f := 0;
        ELSIF x =- 29917 THEN
            exp_f := 0;
        ELSIF x =- 29916 THEN
            exp_f := 0;
        ELSIF x =- 29915 THEN
            exp_f := 0;
        ELSIF x =- 29914 THEN
            exp_f := 0;
        ELSIF x =- 29913 THEN
            exp_f := 0;
        ELSIF x =- 29912 THEN
            exp_f := 0;
        ELSIF x =- 29911 THEN
            exp_f := 0;
        ELSIF x =- 29910 THEN
            exp_f := 0;
        ELSIF x =- 29909 THEN
            exp_f := 0;
        ELSIF x =- 29908 THEN
            exp_f := 0;
        ELSIF x =- 29907 THEN
            exp_f := 0;
        ELSIF x =- 29906 THEN
            exp_f := 0;
        ELSIF x =- 29905 THEN
            exp_f := 0;
        ELSIF x =- 29904 THEN
            exp_f := 0;
        ELSIF x =- 29903 THEN
            exp_f := 0;
        ELSIF x =- 29902 THEN
            exp_f := 0;
        ELSIF x =- 29901 THEN
            exp_f := 0;
        ELSIF x =- 29900 THEN
            exp_f := 0;
        ELSIF x =- 29899 THEN
            exp_f := 0;
        ELSIF x =- 29898 THEN
            exp_f := 0;
        ELSIF x =- 29897 THEN
            exp_f := 0;
        ELSIF x =- 29896 THEN
            exp_f := 0;
        ELSIF x =- 29895 THEN
            exp_f := 0;
        ELSIF x =- 29894 THEN
            exp_f := 0;
        ELSIF x =- 29893 THEN
            exp_f := 0;
        ELSIF x =- 29892 THEN
            exp_f := 0;
        ELSIF x =- 29891 THEN
            exp_f := 0;
        ELSIF x =- 29890 THEN
            exp_f := 0;
        ELSIF x =- 29889 THEN
            exp_f := 0;
        ELSIF x =- 29888 THEN
            exp_f := 0;
        ELSIF x =- 29887 THEN
            exp_f := 0;
        ELSIF x =- 29886 THEN
            exp_f := 0;
        ELSIF x =- 29885 THEN
            exp_f := 0;
        ELSIF x =- 29884 THEN
            exp_f := 0;
        ELSIF x =- 29883 THEN
            exp_f := 0;
        ELSIF x =- 29882 THEN
            exp_f := 0;
        ELSIF x =- 29881 THEN
            exp_f := 0;
        ELSIF x =- 29880 THEN
            exp_f := 0;
        ELSIF x =- 29879 THEN
            exp_f := 0;
        ELSIF x =- 29878 THEN
            exp_f := 0;
        ELSIF x =- 29877 THEN
            exp_f := 0;
        ELSIF x =- 29876 THEN
            exp_f := 0;
        ELSIF x =- 29875 THEN
            exp_f := 0;
        ELSIF x =- 29874 THEN
            exp_f := 0;
        ELSIF x =- 29873 THEN
            exp_f := 0;
        ELSIF x =- 29872 THEN
            exp_f := 0;
        ELSIF x =- 29871 THEN
            exp_f := 0;
        ELSIF x =- 29870 THEN
            exp_f := 0;
        ELSIF x =- 29869 THEN
            exp_f := 0;
        ELSIF x =- 29868 THEN
            exp_f := 0;
        ELSIF x =- 29867 THEN
            exp_f := 0;
        ELSIF x =- 29866 THEN
            exp_f := 0;
        ELSIF x =- 29865 THEN
            exp_f := 0;
        ELSIF x =- 29864 THEN
            exp_f := 0;
        ELSIF x =- 29863 THEN
            exp_f := 0;
        ELSIF x =- 29862 THEN
            exp_f := 0;
        ELSIF x =- 29861 THEN
            exp_f := 0;
        ELSIF x =- 29860 THEN
            exp_f := 0;
        ELSIF x =- 29859 THEN
            exp_f := 0;
        ELSIF x =- 29858 THEN
            exp_f := 0;
        ELSIF x =- 29857 THEN
            exp_f := 0;
        ELSIF x =- 29856 THEN
            exp_f := 0;
        ELSIF x =- 29855 THEN
            exp_f := 0;
        ELSIF x =- 29854 THEN
            exp_f := 0;
        ELSIF x =- 29853 THEN
            exp_f := 0;
        ELSIF x =- 29852 THEN
            exp_f := 0;
        ELSIF x =- 29851 THEN
            exp_f := 0;
        ELSIF x =- 29850 THEN
            exp_f := 0;
        ELSIF x =- 29849 THEN
            exp_f := 0;
        ELSIF x =- 29848 THEN
            exp_f := 0;
        ELSIF x =- 29847 THEN
            exp_f := 0;
        ELSIF x =- 29846 THEN
            exp_f := 0;
        ELSIF x =- 29845 THEN
            exp_f := 0;
        ELSIF x =- 29844 THEN
            exp_f := 0;
        ELSIF x =- 29843 THEN
            exp_f := 0;
        ELSIF x =- 29842 THEN
            exp_f := 0;
        ELSIF x =- 29841 THEN
            exp_f := 0;
        ELSIF x =- 29840 THEN
            exp_f := 0;
        ELSIF x =- 29839 THEN
            exp_f := 0;
        ELSIF x =- 29838 THEN
            exp_f := 0;
        ELSIF x =- 29837 THEN
            exp_f := 0;
        ELSIF x =- 29836 THEN
            exp_f := 0;
        ELSIF x =- 29835 THEN
            exp_f := 0;
        ELSIF x =- 29834 THEN
            exp_f := 0;
        ELSIF x =- 29833 THEN
            exp_f := 0;
        ELSIF x =- 29832 THEN
            exp_f := 0;
        ELSIF x =- 29831 THEN
            exp_f := 0;
        ELSIF x =- 29830 THEN
            exp_f := 0;
        ELSIF x =- 29829 THEN
            exp_f := 0;
        ELSIF x =- 29828 THEN
            exp_f := 0;
        ELSIF x =- 29827 THEN
            exp_f := 0;
        ELSIF x =- 29826 THEN
            exp_f := 0;
        ELSIF x =- 29825 THEN
            exp_f := 0;
        ELSIF x =- 29824 THEN
            exp_f := 0;
        ELSIF x =- 29823 THEN
            exp_f := 0;
        ELSIF x =- 29822 THEN
            exp_f := 0;
        ELSIF x =- 29821 THEN
            exp_f := 0;
        ELSIF x =- 29820 THEN
            exp_f := 0;
        ELSIF x =- 29819 THEN
            exp_f := 0;
        ELSIF x =- 29818 THEN
            exp_f := 0;
        ELSIF x =- 29817 THEN
            exp_f := 0;
        ELSIF x =- 29816 THEN
            exp_f := 0;
        ELSIF x =- 29815 THEN
            exp_f := 0;
        ELSIF x =- 29814 THEN
            exp_f := 0;
        ELSIF x =- 29813 THEN
            exp_f := 0;
        ELSIF x =- 29812 THEN
            exp_f := 0;
        ELSIF x =- 29811 THEN
            exp_f := 0;
        ELSIF x =- 29810 THEN
            exp_f := 0;
        ELSIF x =- 29809 THEN
            exp_f := 0;
        ELSIF x =- 29808 THEN
            exp_f := 0;
        ELSIF x =- 29807 THEN
            exp_f := 0;
        ELSIF x =- 29806 THEN
            exp_f := 0;
        ELSIF x =- 29805 THEN
            exp_f := 0;
        ELSIF x =- 29804 THEN
            exp_f := 0;
        ELSIF x =- 29803 THEN
            exp_f := 0;
        ELSIF x =- 29802 THEN
            exp_f := 0;
        ELSIF x =- 29801 THEN
            exp_f := 0;
        ELSIF x =- 29800 THEN
            exp_f := 0;
        ELSIF x =- 29799 THEN
            exp_f := 0;
        ELSIF x =- 29798 THEN
            exp_f := 0;
        ELSIF x =- 29797 THEN
            exp_f := 0;
        ELSIF x =- 29796 THEN
            exp_f := 0;
        ELSIF x =- 29795 THEN
            exp_f := 0;
        ELSIF x =- 29794 THEN
            exp_f := 0;
        ELSIF x =- 29793 THEN
            exp_f := 0;
        ELSIF x =- 29792 THEN
            exp_f := 0;
        ELSIF x =- 29791 THEN
            exp_f := 0;
        ELSIF x =- 29790 THEN
            exp_f := 0;
        ELSIF x =- 29789 THEN
            exp_f := 0;
        ELSIF x =- 29788 THEN
            exp_f := 0;
        ELSIF x =- 29787 THEN
            exp_f := 0;
        ELSIF x =- 29786 THEN
            exp_f := 0;
        ELSIF x =- 29785 THEN
            exp_f := 0;
        ELSIF x =- 29784 THEN
            exp_f := 0;
        ELSIF x =- 29783 THEN
            exp_f := 0;
        ELSIF x =- 29782 THEN
            exp_f := 0;
        ELSIF x =- 29781 THEN
            exp_f := 0;
        ELSIF x =- 29780 THEN
            exp_f := 0;
        ELSIF x =- 29779 THEN
            exp_f := 0;
        ELSIF x =- 29778 THEN
            exp_f := 0;
        ELSIF x =- 29777 THEN
            exp_f := 0;
        ELSIF x =- 29776 THEN
            exp_f := 0;
        ELSIF x =- 29775 THEN
            exp_f := 0;
        ELSIF x =- 29774 THEN
            exp_f := 0;
        ELSIF x =- 29773 THEN
            exp_f := 0;
        ELSIF x =- 29772 THEN
            exp_f := 0;
        ELSIF x =- 29771 THEN
            exp_f := 0;
        ELSIF x =- 29770 THEN
            exp_f := 0;
        ELSIF x =- 29769 THEN
            exp_f := 0;
        ELSIF x =- 29768 THEN
            exp_f := 0;
        ELSIF x =- 29767 THEN
            exp_f := 0;
        ELSIF x =- 29766 THEN
            exp_f := 0;
        ELSIF x =- 29765 THEN
            exp_f := 0;
        ELSIF x =- 29764 THEN
            exp_f := 0;
        ELSIF x =- 29763 THEN
            exp_f := 0;
        ELSIF x =- 29762 THEN
            exp_f := 0;
        ELSIF x =- 29761 THEN
            exp_f := 0;
        ELSIF x =- 29760 THEN
            exp_f := 0;
        ELSIF x =- 29759 THEN
            exp_f := 0;
        ELSIF x =- 29758 THEN
            exp_f := 0;
        ELSIF x =- 29757 THEN
            exp_f := 0;
        ELSIF x =- 29756 THEN
            exp_f := 0;
        ELSIF x =- 29755 THEN
            exp_f := 0;
        ELSIF x =- 29754 THEN
            exp_f := 0;
        ELSIF x =- 29753 THEN
            exp_f := 0;
        ELSIF x =- 29752 THEN
            exp_f := 0;
        ELSIF x =- 29751 THEN
            exp_f := 0;
        ELSIF x =- 29750 THEN
            exp_f := 0;
        ELSIF x =- 29749 THEN
            exp_f := 0;
        ELSIF x =- 29748 THEN
            exp_f := 0;
        ELSIF x =- 29747 THEN
            exp_f := 0;
        ELSIF x =- 29746 THEN
            exp_f := 0;
        ELSIF x =- 29745 THEN
            exp_f := 0;
        ELSIF x =- 29744 THEN
            exp_f := 0;
        ELSIF x =- 29743 THEN
            exp_f := 0;
        ELSIF x =- 29742 THEN
            exp_f := 0;
        ELSIF x =- 29741 THEN
            exp_f := 0;
        ELSIF x =- 29740 THEN
            exp_f := 0;
        ELSIF x =- 29739 THEN
            exp_f := 0;
        ELSIF x =- 29738 THEN
            exp_f := 0;
        ELSIF x =- 29737 THEN
            exp_f := 0;
        ELSIF x =- 29736 THEN
            exp_f := 0;
        ELSIF x =- 29735 THEN
            exp_f := 0;
        ELSIF x =- 29734 THEN
            exp_f := 0;
        ELSIF x =- 29733 THEN
            exp_f := 0;
        ELSIF x =- 29732 THEN
            exp_f := 0;
        ELSIF x =- 29731 THEN
            exp_f := 0;
        ELSIF x =- 29730 THEN
            exp_f := 0;
        ELSIF x =- 29729 THEN
            exp_f := 0;
        ELSIF x =- 29728 THEN
            exp_f := 0;
        ELSIF x =- 29727 THEN
            exp_f := 0;
        ELSIF x =- 29726 THEN
            exp_f := 0;
        ELSIF x =- 29725 THEN
            exp_f := 0;
        ELSIF x =- 29724 THEN
            exp_f := 0;
        ELSIF x =- 29723 THEN
            exp_f := 0;
        ELSIF x =- 29722 THEN
            exp_f := 0;
        ELSIF x =- 29721 THEN
            exp_f := 0;
        ELSIF x =- 29720 THEN
            exp_f := 0;
        ELSIF x =- 29719 THEN
            exp_f := 0;
        ELSIF x =- 29718 THEN
            exp_f := 0;
        ELSIF x =- 29717 THEN
            exp_f := 0;
        ELSIF x =- 29716 THEN
            exp_f := 0;
        ELSIF x =- 29715 THEN
            exp_f := 0;
        ELSIF x =- 29714 THEN
            exp_f := 0;
        ELSIF x =- 29713 THEN
            exp_f := 0;
        ELSIF x =- 29712 THEN
            exp_f := 0;
        ELSIF x =- 29711 THEN
            exp_f := 0;
        ELSIF x =- 29710 THEN
            exp_f := 0;
        ELSIF x =- 29709 THEN
            exp_f := 0;
        ELSIF x =- 29708 THEN
            exp_f := 0;
        ELSIF x =- 29707 THEN
            exp_f := 0;
        ELSIF x =- 29706 THEN
            exp_f := 0;
        ELSIF x =- 29705 THEN
            exp_f := 0;
        ELSIF x =- 29704 THEN
            exp_f := 0;
        ELSIF x =- 29703 THEN
            exp_f := 0;
        ELSIF x =- 29702 THEN
            exp_f := 0;
        ELSIF x =- 29701 THEN
            exp_f := 0;
        ELSIF x =- 29700 THEN
            exp_f := 0;
        ELSIF x =- 29699 THEN
            exp_f := 0;
        ELSIF x =- 29698 THEN
            exp_f := 0;
        ELSIF x =- 29697 THEN
            exp_f := 0;
        ELSIF x =- 29696 THEN
            exp_f := 0;
        ELSIF x =- 29695 THEN
            exp_f := 0;
        ELSIF x =- 29694 THEN
            exp_f := 0;
        ELSIF x =- 29693 THEN
            exp_f := 0;
        ELSIF x =- 29692 THEN
            exp_f := 0;
        ELSIF x =- 29691 THEN
            exp_f := 0;
        ELSIF x =- 29690 THEN
            exp_f := 0;
        ELSIF x =- 29689 THEN
            exp_f := 0;
        ELSIF x =- 29688 THEN
            exp_f := 0;
        ELSIF x =- 29687 THEN
            exp_f := 0;
        ELSIF x =- 29686 THEN
            exp_f := 0;
        ELSIF x =- 29685 THEN
            exp_f := 0;
        ELSIF x =- 29684 THEN
            exp_f := 0;
        ELSIF x =- 29683 THEN
            exp_f := 0;
        ELSIF x =- 29682 THEN
            exp_f := 0;
        ELSIF x =- 29681 THEN
            exp_f := 0;
        ELSIF x =- 29680 THEN
            exp_f := 0;
        ELSIF x =- 29679 THEN
            exp_f := 0;
        ELSIF x =- 29678 THEN
            exp_f := 0;
        ELSIF x =- 29677 THEN
            exp_f := 0;
        ELSIF x =- 29676 THEN
            exp_f := 0;
        ELSIF x =- 29675 THEN
            exp_f := 0;
        ELSIF x =- 29674 THEN
            exp_f := 0;
        ELSIF x =- 29673 THEN
            exp_f := 0;
        ELSIF x =- 29672 THEN
            exp_f := 0;
        ELSIF x =- 29671 THEN
            exp_f := 0;
        ELSIF x =- 29670 THEN
            exp_f := 0;
        ELSIF x =- 29669 THEN
            exp_f := 0;
        ELSIF x =- 29668 THEN
            exp_f := 0;
        ELSIF x =- 29667 THEN
            exp_f := 0;
        ELSIF x =- 29666 THEN
            exp_f := 0;
        ELSIF x =- 29665 THEN
            exp_f := 0;
        ELSIF x =- 29664 THEN
            exp_f := 0;
        ELSIF x =- 29663 THEN
            exp_f := 0;
        ELSIF x =- 29662 THEN
            exp_f := 0;
        ELSIF x =- 29661 THEN
            exp_f := 0;
        ELSIF x =- 29660 THEN
            exp_f := 0;
        ELSIF x =- 29659 THEN
            exp_f := 0;
        ELSIF x =- 29658 THEN
            exp_f := 0;
        ELSIF x =- 29657 THEN
            exp_f := 0;
        ELSIF x =- 29656 THEN
            exp_f := 0;
        ELSIF x =- 29655 THEN
            exp_f := 0;
        ELSIF x =- 29654 THEN
            exp_f := 0;
        ELSIF x =- 29653 THEN
            exp_f := 0;
        ELSIF x =- 29652 THEN
            exp_f := 0;
        ELSIF x =- 29651 THEN
            exp_f := 0;
        ELSIF x =- 29650 THEN
            exp_f := 0;
        ELSIF x =- 29649 THEN
            exp_f := 0;
        ELSIF x =- 29648 THEN
            exp_f := 0;
        ELSIF x =- 29647 THEN
            exp_f := 0;
        ELSIF x =- 29646 THEN
            exp_f := 0;
        ELSIF x =- 29645 THEN
            exp_f := 0;
        ELSIF x =- 29644 THEN
            exp_f := 0;
        ELSIF x =- 29643 THEN
            exp_f := 0;
        ELSIF x =- 29642 THEN
            exp_f := 0;
        ELSIF x =- 29641 THEN
            exp_f := 0;
        ELSIF x =- 29640 THEN
            exp_f := 0;
        ELSIF x =- 29639 THEN
            exp_f := 0;
        ELSIF x =- 29638 THEN
            exp_f := 0;
        ELSIF x =- 29637 THEN
            exp_f := 0;
        ELSIF x =- 29636 THEN
            exp_f := 0;
        ELSIF x =- 29635 THEN
            exp_f := 0;
        ELSIF x =- 29634 THEN
            exp_f := 0;
        ELSIF x =- 29633 THEN
            exp_f := 0;
        ELSIF x =- 29632 THEN
            exp_f := 0;
        ELSIF x =- 29631 THEN
            exp_f := 0;
        ELSIF x =- 29630 THEN
            exp_f := 0;
        ELSIF x =- 29629 THEN
            exp_f := 0;
        ELSIF x =- 29628 THEN
            exp_f := 0;
        ELSIF x =- 29627 THEN
            exp_f := 0;
        ELSIF x =- 29626 THEN
            exp_f := 0;
        ELSIF x =- 29625 THEN
            exp_f := 0;
        ELSIF x =- 29624 THEN
            exp_f := 0;
        ELSIF x =- 29623 THEN
            exp_f := 0;
        ELSIF x =- 29622 THEN
            exp_f := 0;
        ELSIF x =- 29621 THEN
            exp_f := 0;
        ELSIF x =- 29620 THEN
            exp_f := 0;
        ELSIF x =- 29619 THEN
            exp_f := 0;
        ELSIF x =- 29618 THEN
            exp_f := 0;
        ELSIF x =- 29617 THEN
            exp_f := 0;
        ELSIF x =- 29616 THEN
            exp_f := 0;
        ELSIF x =- 29615 THEN
            exp_f := 0;
        ELSIF x =- 29614 THEN
            exp_f := 0;
        ELSIF x =- 29613 THEN
            exp_f := 0;
        ELSIF x =- 29612 THEN
            exp_f := 0;
        ELSIF x =- 29611 THEN
            exp_f := 0;
        ELSIF x =- 29610 THEN
            exp_f := 0;
        ELSIF x =- 29609 THEN
            exp_f := 0;
        ELSIF x =- 29608 THEN
            exp_f := 0;
        ELSIF x =- 29607 THEN
            exp_f := 0;
        ELSIF x =- 29606 THEN
            exp_f := 0;
        ELSIF x =- 29605 THEN
            exp_f := 0;
        ELSIF x =- 29604 THEN
            exp_f := 0;
        ELSIF x =- 29603 THEN
            exp_f := 0;
        ELSIF x =- 29602 THEN
            exp_f := 0;
        ELSIF x =- 29601 THEN
            exp_f := 0;
        ELSIF x =- 29600 THEN
            exp_f := 0;
        ELSIF x =- 29599 THEN
            exp_f := 0;
        ELSIF x =- 29598 THEN
            exp_f := 0;
        ELSIF x =- 29597 THEN
            exp_f := 0;
        ELSIF x =- 29596 THEN
            exp_f := 0;
        ELSIF x =- 29595 THEN
            exp_f := 0;
        ELSIF x =- 29594 THEN
            exp_f := 0;
        ELSIF x =- 29593 THEN
            exp_f := 0;
        ELSIF x =- 29592 THEN
            exp_f := 0;
        ELSIF x =- 29591 THEN
            exp_f := 0;
        ELSIF x =- 29590 THEN
            exp_f := 0;
        ELSIF x =- 29589 THEN
            exp_f := 0;
        ELSIF x =- 29588 THEN
            exp_f := 0;
        ELSIF x =- 29587 THEN
            exp_f := 0;
        ELSIF x =- 29586 THEN
            exp_f := 0;
        ELSIF x =- 29585 THEN
            exp_f := 0;
        ELSIF x =- 29584 THEN
            exp_f := 0;
        ELSIF x =- 29583 THEN
            exp_f := 0;
        ELSIF x =- 29582 THEN
            exp_f := 0;
        ELSIF x =- 29581 THEN
            exp_f := 0;
        ELSIF x =- 29580 THEN
            exp_f := 0;
        ELSIF x =- 29579 THEN
            exp_f := 0;
        ELSIF x =- 29578 THEN
            exp_f := 0;
        ELSIF x =- 29577 THEN
            exp_f := 0;
        ELSIF x =- 29576 THEN
            exp_f := 0;
        ELSIF x =- 29575 THEN
            exp_f := 0;
        ELSIF x =- 29574 THEN
            exp_f := 0;
        ELSIF x =- 29573 THEN
            exp_f := 0;
        ELSIF x =- 29572 THEN
            exp_f := 0;
        ELSIF x =- 29571 THEN
            exp_f := 0;
        ELSIF x =- 29570 THEN
            exp_f := 0;
        ELSIF x =- 29569 THEN
            exp_f := 0;
        ELSIF x =- 29568 THEN
            exp_f := 0;
        ELSIF x =- 29567 THEN
            exp_f := 0;
        ELSIF x =- 29566 THEN
            exp_f := 0;
        ELSIF x =- 29565 THEN
            exp_f := 0;
        ELSIF x =- 29564 THEN
            exp_f := 0;
        ELSIF x =- 29563 THEN
            exp_f := 0;
        ELSIF x =- 29562 THEN
            exp_f := 0;
        ELSIF x =- 29561 THEN
            exp_f := 0;
        ELSIF x =- 29560 THEN
            exp_f := 0;
        ELSIF x =- 29559 THEN
            exp_f := 0;
        ELSIF x =- 29558 THEN
            exp_f := 0;
        ELSIF x =- 29557 THEN
            exp_f := 0;
        ELSIF x =- 29556 THEN
            exp_f := 0;
        ELSIF x =- 29555 THEN
            exp_f := 0;
        ELSIF x =- 29554 THEN
            exp_f := 0;
        ELSIF x =- 29553 THEN
            exp_f := 0;
        ELSIF x =- 29552 THEN
            exp_f := 0;
        ELSIF x =- 29551 THEN
            exp_f := 0;
        ELSIF x =- 29550 THEN
            exp_f := 0;
        ELSIF x =- 29549 THEN
            exp_f := 0;
        ELSIF x =- 29548 THEN
            exp_f := 0;
        ELSIF x =- 29547 THEN
            exp_f := 0;
        ELSIF x =- 29546 THEN
            exp_f := 0;
        ELSIF x =- 29545 THEN
            exp_f := 0;
        ELSIF x =- 29544 THEN
            exp_f := 0;
        ELSIF x =- 29543 THEN
            exp_f := 0;
        ELSIF x =- 29542 THEN
            exp_f := 0;
        ELSIF x =- 29541 THEN
            exp_f := 0;
        ELSIF x =- 29540 THEN
            exp_f := 0;
        ELSIF x =- 29539 THEN
            exp_f := 0;
        ELSIF x =- 29538 THEN
            exp_f := 0;
        ELSIF x =- 29537 THEN
            exp_f := 0;
        ELSIF x =- 29536 THEN
            exp_f := 0;
        ELSIF x =- 29535 THEN
            exp_f := 0;
        ELSIF x =- 29534 THEN
            exp_f := 0;
        ELSIF x =- 29533 THEN
            exp_f := 0;
        ELSIF x =- 29532 THEN
            exp_f := 0;
        ELSIF x =- 29531 THEN
            exp_f := 0;
        ELSIF x =- 29530 THEN
            exp_f := 0;
        ELSIF x =- 29529 THEN
            exp_f := 0;
        ELSIF x =- 29528 THEN
            exp_f := 0;
        ELSIF x =- 29527 THEN
            exp_f := 0;
        ELSIF x =- 29526 THEN
            exp_f := 0;
        ELSIF x =- 29525 THEN
            exp_f := 0;
        ELSIF x =- 29524 THEN
            exp_f := 0;
        ELSIF x =- 29523 THEN
            exp_f := 0;
        ELSIF x =- 29522 THEN
            exp_f := 0;
        ELSIF x =- 29521 THEN
            exp_f := 0;
        ELSIF x =- 29520 THEN
            exp_f := 0;
        ELSIF x =- 29519 THEN
            exp_f := 0;
        ELSIF x =- 29518 THEN
            exp_f := 0;
        ELSIF x =- 29517 THEN
            exp_f := 0;
        ELSIF x =- 29516 THEN
            exp_f := 0;
        ELSIF x =- 29515 THEN
            exp_f := 0;
        ELSIF x =- 29514 THEN
            exp_f := 0;
        ELSIF x =- 29513 THEN
            exp_f := 0;
        ELSIF x =- 29512 THEN
            exp_f := 0;
        ELSIF x =- 29511 THEN
            exp_f := 0;
        ELSIF x =- 29510 THEN
            exp_f := 0;
        ELSIF x =- 29509 THEN
            exp_f := 0;
        ELSIF x =- 29508 THEN
            exp_f := 0;
        ELSIF x =- 29507 THEN
            exp_f := 0;
        ELSIF x =- 29506 THEN
            exp_f := 0;
        ELSIF x =- 29505 THEN
            exp_f := 0;
        ELSIF x =- 29504 THEN
            exp_f := 0;
        ELSIF x =- 29503 THEN
            exp_f := 0;
        ELSIF x =- 29502 THEN
            exp_f := 0;
        ELSIF x =- 29501 THEN
            exp_f := 0;
        ELSIF x =- 29500 THEN
            exp_f := 0;
        ELSIF x =- 29499 THEN
            exp_f := 0;
        ELSIF x =- 29498 THEN
            exp_f := 0;
        ELSIF x =- 29497 THEN
            exp_f := 0;
        ELSIF x =- 29496 THEN
            exp_f := 0;
        ELSIF x =- 29495 THEN
            exp_f := 0;
        ELSIF x =- 29494 THEN
            exp_f := 0;
        ELSIF x =- 29493 THEN
            exp_f := 0;
        ELSIF x =- 29492 THEN
            exp_f := 0;
        ELSIF x =- 29491 THEN
            exp_f := 0;
        ELSIF x =- 29490 THEN
            exp_f := 0;
        ELSIF x =- 29489 THEN
            exp_f := 0;
        ELSIF x =- 29488 THEN
            exp_f := 0;
        ELSIF x =- 29487 THEN
            exp_f := 0;
        ELSIF x =- 29486 THEN
            exp_f := 0;
        ELSIF x =- 29485 THEN
            exp_f := 0;
        ELSIF x =- 29484 THEN
            exp_f := 0;
        ELSIF x =- 29483 THEN
            exp_f := 0;
        ELSIF x =- 29482 THEN
            exp_f := 0;
        ELSIF x =- 29481 THEN
            exp_f := 0;
        ELSIF x =- 29480 THEN
            exp_f := 0;
        ELSIF x =- 29479 THEN
            exp_f := 0;
        ELSIF x =- 29478 THEN
            exp_f := 0;
        ELSIF x =- 29477 THEN
            exp_f := 0;
        ELSIF x =- 29476 THEN
            exp_f := 0;
        ELSIF x =- 29475 THEN
            exp_f := 0;
        ELSIF x =- 29474 THEN
            exp_f := 0;
        ELSIF x =- 29473 THEN
            exp_f := 0;
        ELSIF x =- 29472 THEN
            exp_f := 0;
        ELSIF x =- 29471 THEN
            exp_f := 0;
        ELSIF x =- 29470 THEN
            exp_f := 0;
        ELSIF x =- 29469 THEN
            exp_f := 0;
        ELSIF x =- 29468 THEN
            exp_f := 0;
        ELSIF x =- 29467 THEN
            exp_f := 0;
        ELSIF x =- 29466 THEN
            exp_f := 0;
        ELSIF x =- 29465 THEN
            exp_f := 0;
        ELSIF x =- 29464 THEN
            exp_f := 0;
        ELSIF x =- 29463 THEN
            exp_f := 0;
        ELSIF x =- 29462 THEN
            exp_f := 0;
        ELSIF x =- 29461 THEN
            exp_f := 0;
        ELSIF x =- 29460 THEN
            exp_f := 0;
        ELSIF x =- 29459 THEN
            exp_f := 0;
        ELSIF x =- 29458 THEN
            exp_f := 0;
        ELSIF x =- 29457 THEN
            exp_f := 0;
        ELSIF x =- 29456 THEN
            exp_f := 0;
        ELSIF x =- 29455 THEN
            exp_f := 0;
        ELSIF x =- 29454 THEN
            exp_f := 0;
        ELSIF x =- 29453 THEN
            exp_f := 0;
        ELSIF x =- 29452 THEN
            exp_f := 0;
        ELSIF x =- 29451 THEN
            exp_f := 0;
        ELSIF x =- 29450 THEN
            exp_f := 0;
        ELSIF x =- 29449 THEN
            exp_f := 0;
        ELSIF x =- 29448 THEN
            exp_f := 0;
        ELSIF x =- 29447 THEN
            exp_f := 0;
        ELSIF x =- 29446 THEN
            exp_f := 0;
        ELSIF x =- 29445 THEN
            exp_f := 0;
        ELSIF x =- 29444 THEN
            exp_f := 0;
        ELSIF x =- 29443 THEN
            exp_f := 0;
        ELSIF x =- 29442 THEN
            exp_f := 0;
        ELSIF x =- 29441 THEN
            exp_f := 0;
        ELSIF x =- 29440 THEN
            exp_f := 0;
        ELSIF x =- 29439 THEN
            exp_f := 0;
        ELSIF x =- 29438 THEN
            exp_f := 0;
        ELSIF x =- 29437 THEN
            exp_f := 0;
        ELSIF x =- 29436 THEN
            exp_f := 0;
        ELSIF x =- 29435 THEN
            exp_f := 0;
        ELSIF x =- 29434 THEN
            exp_f := 0;
        ELSIF x =- 29433 THEN
            exp_f := 0;
        ELSIF x =- 29432 THEN
            exp_f := 0;
        ELSIF x =- 29431 THEN
            exp_f := 0;
        ELSIF x =- 29430 THEN
            exp_f := 0;
        ELSIF x =- 29429 THEN
            exp_f := 0;
        ELSIF x =- 29428 THEN
            exp_f := 0;
        ELSIF x =- 29427 THEN
            exp_f := 0;
        ELSIF x =- 29426 THEN
            exp_f := 0;
        ELSIF x =- 29425 THEN
            exp_f := 0;
        ELSIF x =- 29424 THEN
            exp_f := 0;
        ELSIF x =- 29423 THEN
            exp_f := 0;
        ELSIF x =- 29422 THEN
            exp_f := 0;
        ELSIF x =- 29421 THEN
            exp_f := 0;
        ELSIF x =- 29420 THEN
            exp_f := 0;
        ELSIF x =- 29419 THEN
            exp_f := 0;
        ELSIF x =- 29418 THEN
            exp_f := 0;
        ELSIF x =- 29417 THEN
            exp_f := 0;
        ELSIF x =- 29416 THEN
            exp_f := 0;
        ELSIF x =- 29415 THEN
            exp_f := 0;
        ELSIF x =- 29414 THEN
            exp_f := 0;
        ELSIF x =- 29413 THEN
            exp_f := 0;
        ELSIF x =- 29412 THEN
            exp_f := 0;
        ELSIF x =- 29411 THEN
            exp_f := 0;
        ELSIF x =- 29410 THEN
            exp_f := 0;
        ELSIF x =- 29409 THEN
            exp_f := 0;
        ELSIF x =- 29408 THEN
            exp_f := 0;
        ELSIF x =- 29407 THEN
            exp_f := 0;
        ELSIF x =- 29406 THEN
            exp_f := 0;
        ELSIF x =- 29405 THEN
            exp_f := 0;
        ELSIF x =- 29404 THEN
            exp_f := 0;
        ELSIF x =- 29403 THEN
            exp_f := 0;
        ELSIF x =- 29402 THEN
            exp_f := 0;
        ELSIF x =- 29401 THEN
            exp_f := 0;
        ELSIF x =- 29400 THEN
            exp_f := 0;
        ELSIF x =- 29399 THEN
            exp_f := 0;
        ELSIF x =- 29398 THEN
            exp_f := 0;
        ELSIF x =- 29397 THEN
            exp_f := 0;
        ELSIF x =- 29396 THEN
            exp_f := 0;
        ELSIF x =- 29395 THEN
            exp_f := 0;
        ELSIF x =- 29394 THEN
            exp_f := 0;
        ELSIF x =- 29393 THEN
            exp_f := 0;
        ELSIF x =- 29392 THEN
            exp_f := 0;
        ELSIF x =- 29391 THEN
            exp_f := 0;
        ELSIF x =- 29390 THEN
            exp_f := 0;
        ELSIF x =- 29389 THEN
            exp_f := 0;
        ELSIF x =- 29388 THEN
            exp_f := 0;
        ELSIF x =- 29387 THEN
            exp_f := 0;
        ELSIF x =- 29386 THEN
            exp_f := 0;
        ELSIF x =- 29385 THEN
            exp_f := 0;
        ELSIF x =- 29384 THEN
            exp_f := 0;
        ELSIF x =- 29383 THEN
            exp_f := 0;
        ELSIF x =- 29382 THEN
            exp_f := 0;
        ELSIF x =- 29381 THEN
            exp_f := 0;
        ELSIF x =- 29380 THEN
            exp_f := 0;
        ELSIF x =- 29379 THEN
            exp_f := 0;
        ELSIF x =- 29378 THEN
            exp_f := 0;
        ELSIF x =- 29377 THEN
            exp_f := 0;
        ELSIF x =- 29376 THEN
            exp_f := 0;
        ELSIF x =- 29375 THEN
            exp_f := 0;
        ELSIF x =- 29374 THEN
            exp_f := 0;
        ELSIF x =- 29373 THEN
            exp_f := 0;
        ELSIF x =- 29372 THEN
            exp_f := 0;
        ELSIF x =- 29371 THEN
            exp_f := 0;
        ELSIF x =- 29370 THEN
            exp_f := 0;
        ELSIF x =- 29369 THEN
            exp_f := 0;
        ELSIF x =- 29368 THEN
            exp_f := 0;
        ELSIF x =- 29367 THEN
            exp_f := 0;
        ELSIF x =- 29366 THEN
            exp_f := 0;
        ELSIF x =- 29365 THEN
            exp_f := 0;
        ELSIF x =- 29364 THEN
            exp_f := 0;
        ELSIF x =- 29363 THEN
            exp_f := 0;
        ELSIF x =- 29362 THEN
            exp_f := 0;
        ELSIF x =- 29361 THEN
            exp_f := 0;
        ELSIF x =- 29360 THEN
            exp_f := 0;
        ELSIF x =- 29359 THEN
            exp_f := 0;
        ELSIF x =- 29358 THEN
            exp_f := 0;
        ELSIF x =- 29357 THEN
            exp_f := 0;
        ELSIF x =- 29356 THEN
            exp_f := 0;
        ELSIF x =- 29355 THEN
            exp_f := 0;
        ELSIF x =- 29354 THEN
            exp_f := 0;
        ELSIF x =- 29353 THEN
            exp_f := 0;
        ELSIF x =- 29352 THEN
            exp_f := 0;
        ELSIF x =- 29351 THEN
            exp_f := 0;
        ELSIF x =- 29350 THEN
            exp_f := 0;
        ELSIF x =- 29349 THEN
            exp_f := 0;
        ELSIF x =- 29348 THEN
            exp_f := 0;
        ELSIF x =- 29347 THEN
            exp_f := 0;
        ELSIF x =- 29346 THEN
            exp_f := 0;
        ELSIF x =- 29345 THEN
            exp_f := 0;
        ELSIF x =- 29344 THEN
            exp_f := 0;
        ELSIF x =- 29343 THEN
            exp_f := 0;
        ELSIF x =- 29342 THEN
            exp_f := 0;
        ELSIF x =- 29341 THEN
            exp_f := 0;
        ELSIF x =- 29340 THEN
            exp_f := 0;
        ELSIF x =- 29339 THEN
            exp_f := 0;
        ELSIF x =- 29338 THEN
            exp_f := 0;
        ELSIF x =- 29337 THEN
            exp_f := 0;
        ELSIF x =- 29336 THEN
            exp_f := 0;
        ELSIF x =- 29335 THEN
            exp_f := 0;
        ELSIF x =- 29334 THEN
            exp_f := 0;
        ELSIF x =- 29333 THEN
            exp_f := 0;
        ELSIF x =- 29332 THEN
            exp_f := 0;
        ELSIF x =- 29331 THEN
            exp_f := 0;
        ELSIF x =- 29330 THEN
            exp_f := 0;
        ELSIF x =- 29329 THEN
            exp_f := 0;
        ELSIF x =- 29328 THEN
            exp_f := 0;
        ELSIF x =- 29327 THEN
            exp_f := 0;
        ELSIF x =- 29326 THEN
            exp_f := 0;
        ELSIF x =- 29325 THEN
            exp_f := 0;
        ELSIF x =- 29324 THEN
            exp_f := 0;
        ELSIF x =- 29323 THEN
            exp_f := 0;
        ELSIF x =- 29322 THEN
            exp_f := 0;
        ELSIF x =- 29321 THEN
            exp_f := 0;
        ELSIF x =- 29320 THEN
            exp_f := 0;
        ELSIF x =- 29319 THEN
            exp_f := 0;
        ELSIF x =- 29318 THEN
            exp_f := 0;
        ELSIF x =- 29317 THEN
            exp_f := 0;
        ELSIF x =- 29316 THEN
            exp_f := 0;
        ELSIF x =- 29315 THEN
            exp_f := 0;
        ELSIF x =- 29314 THEN
            exp_f := 0;
        ELSIF x =- 29313 THEN
            exp_f := 0;
        ELSIF x =- 29312 THEN
            exp_f := 0;
        ELSIF x =- 29311 THEN
            exp_f := 0;
        ELSIF x =- 29310 THEN
            exp_f := 0;
        ELSIF x =- 29309 THEN
            exp_f := 0;
        ELSIF x =- 29308 THEN
            exp_f := 0;
        ELSIF x =- 29307 THEN
            exp_f := 0;
        ELSIF x =- 29306 THEN
            exp_f := 0;
        ELSIF x =- 29305 THEN
            exp_f := 0;
        ELSIF x =- 29304 THEN
            exp_f := 0;
        ELSIF x =- 29303 THEN
            exp_f := 0;
        ELSIF x =- 29302 THEN
            exp_f := 0;
        ELSIF x =- 29301 THEN
            exp_f := 0;
        ELSIF x =- 29300 THEN
            exp_f := 0;
        ELSIF x =- 29299 THEN
            exp_f := 0;
        ELSIF x =- 29298 THEN
            exp_f := 0;
        ELSIF x =- 29297 THEN
            exp_f := 0;
        ELSIF x =- 29296 THEN
            exp_f := 0;
        ELSIF x =- 29295 THEN
            exp_f := 0;
        ELSIF x =- 29294 THEN
            exp_f := 0;
        ELSIF x =- 29293 THEN
            exp_f := 0;
        ELSIF x =- 29292 THEN
            exp_f := 0;
        ELSIF x =- 29291 THEN
            exp_f := 0;
        ELSIF x =- 29290 THEN
            exp_f := 0;
        ELSIF x =- 29289 THEN
            exp_f := 0;
        ELSIF x =- 29288 THEN
            exp_f := 0;
        ELSIF x =- 29287 THEN
            exp_f := 0;
        ELSIF x =- 29286 THEN
            exp_f := 0;
        ELSIF x =- 29285 THEN
            exp_f := 0;
        ELSIF x =- 29284 THEN
            exp_f := 0;
        ELSIF x =- 29283 THEN
            exp_f := 0;
        ELSIF x =- 29282 THEN
            exp_f := 0;
        ELSIF x =- 29281 THEN
            exp_f := 0;
        ELSIF x =- 29280 THEN
            exp_f := 0;
        ELSIF x =- 29279 THEN
            exp_f := 0;
        ELSIF x =- 29278 THEN
            exp_f := 0;
        ELSIF x =- 29277 THEN
            exp_f := 0;
        ELSIF x =- 29276 THEN
            exp_f := 0;
        ELSIF x =- 29275 THEN
            exp_f := 0;
        ELSIF x =- 29274 THEN
            exp_f := 0;
        ELSIF x =- 29273 THEN
            exp_f := 0;
        ELSIF x =- 29272 THEN
            exp_f := 0;
        ELSIF x =- 29271 THEN
            exp_f := 0;
        ELSIF x =- 29270 THEN
            exp_f := 0;
        ELSIF x =- 29269 THEN
            exp_f := 0;
        ELSIF x =- 29268 THEN
            exp_f := 0;
        ELSIF x =- 29267 THEN
            exp_f := 0;
        ELSIF x =- 29266 THEN
            exp_f := 0;
        ELSIF x =- 29265 THEN
            exp_f := 0;
        ELSIF x =- 29264 THEN
            exp_f := 0;
        ELSIF x =- 29263 THEN
            exp_f := 0;
        ELSIF x =- 29262 THEN
            exp_f := 0;
        ELSIF x =- 29261 THEN
            exp_f := 0;
        ELSIF x =- 29260 THEN
            exp_f := 0;
        ELSIF x =- 29259 THEN
            exp_f := 0;
        ELSIF x =- 29258 THEN
            exp_f := 0;
        ELSIF x =- 29257 THEN
            exp_f := 0;
        ELSIF x =- 29256 THEN
            exp_f := 0;
        ELSIF x =- 29255 THEN
            exp_f := 0;
        ELSIF x =- 29254 THEN
            exp_f := 0;
        ELSIF x =- 29253 THEN
            exp_f := 0;
        ELSIF x =- 29252 THEN
            exp_f := 0;
        ELSIF x =- 29251 THEN
            exp_f := 0;
        ELSIF x =- 29250 THEN
            exp_f := 0;
        ELSIF x =- 29249 THEN
            exp_f := 0;
        ELSIF x =- 29248 THEN
            exp_f := 0;
        ELSIF x =- 29247 THEN
            exp_f := 0;
        ELSIF x =- 29246 THEN
            exp_f := 0;
        ELSIF x =- 29245 THEN
            exp_f := 0;
        ELSIF x =- 29244 THEN
            exp_f := 0;
        ELSIF x =- 29243 THEN
            exp_f := 0;
        ELSIF x =- 29242 THEN
            exp_f := 0;
        ELSIF x =- 29241 THEN
            exp_f := 0;
        ELSIF x =- 29240 THEN
            exp_f := 0;
        ELSIF x =- 29239 THEN
            exp_f := 0;
        ELSIF x =- 29238 THEN
            exp_f := 0;
        ELSIF x =- 29237 THEN
            exp_f := 0;
        ELSIF x =- 29236 THEN
            exp_f := 0;
        ELSIF x =- 29235 THEN
            exp_f := 0;
        ELSIF x =- 29234 THEN
            exp_f := 0;
        ELSIF x =- 29233 THEN
            exp_f := 0;
        ELSIF x =- 29232 THEN
            exp_f := 0;
        ELSIF x =- 29231 THEN
            exp_f := 0;
        ELSIF x =- 29230 THEN
            exp_f := 0;
        ELSIF x =- 29229 THEN
            exp_f := 0;
        ELSIF x =- 29228 THEN
            exp_f := 0;
        ELSIF x =- 29227 THEN
            exp_f := 0;
        ELSIF x =- 29226 THEN
            exp_f := 0;
        ELSIF x =- 29225 THEN
            exp_f := 0;
        ELSIF x =- 29224 THEN
            exp_f := 0;
        ELSIF x =- 29223 THEN
            exp_f := 0;
        ELSIF x =- 29222 THEN
            exp_f := 0;
        ELSIF x =- 29221 THEN
            exp_f := 0;
        ELSIF x =- 29220 THEN
            exp_f := 0;
        ELSIF x =- 29219 THEN
            exp_f := 0;
        ELSIF x =- 29218 THEN
            exp_f := 0;
        ELSIF x =- 29217 THEN
            exp_f := 0;
        ELSIF x =- 29216 THEN
            exp_f := 0;
        ELSIF x =- 29215 THEN
            exp_f := 0;
        ELSIF x =- 29214 THEN
            exp_f := 0;
        ELSIF x =- 29213 THEN
            exp_f := 0;
        ELSIF x =- 29212 THEN
            exp_f := 0;
        ELSIF x =- 29211 THEN
            exp_f := 0;
        ELSIF x =- 29210 THEN
            exp_f := 0;
        ELSIF x =- 29209 THEN
            exp_f := 0;
        ELSIF x =- 29208 THEN
            exp_f := 0;
        ELSIF x =- 29207 THEN
            exp_f := 0;
        ELSIF x =- 29206 THEN
            exp_f := 0;
        ELSIF x =- 29205 THEN
            exp_f := 0;
        ELSIF x =- 29204 THEN
            exp_f := 0;
        ELSIF x =- 29203 THEN
            exp_f := 0;
        ELSIF x =- 29202 THEN
            exp_f := 0;
        ELSIF x =- 29201 THEN
            exp_f := 0;
        ELSIF x =- 29200 THEN
            exp_f := 0;
        ELSIF x =- 29199 THEN
            exp_f := 0;
        ELSIF x =- 29198 THEN
            exp_f := 0;
        ELSIF x =- 29197 THEN
            exp_f := 0;
        ELSIF x =- 29196 THEN
            exp_f := 0;
        ELSIF x =- 29195 THEN
            exp_f := 0;
        ELSIF x =- 29194 THEN
            exp_f := 0;
        ELSIF x =- 29193 THEN
            exp_f := 0;
        ELSIF x =- 29192 THEN
            exp_f := 0;
        ELSIF x =- 29191 THEN
            exp_f := 0;
        ELSIF x =- 29190 THEN
            exp_f := 0;
        ELSIF x =- 29189 THEN
            exp_f := 0;
        ELSIF x =- 29188 THEN
            exp_f := 0;
        ELSIF x =- 29187 THEN
            exp_f := 0;
        ELSIF x =- 29186 THEN
            exp_f := 0;
        ELSIF x =- 29185 THEN
            exp_f := 0;
        ELSIF x =- 29184 THEN
            exp_f := 0;
        ELSIF x =- 29183 THEN
            exp_f := 0;
        ELSIF x =- 29182 THEN
            exp_f := 0;
        ELSIF x =- 29181 THEN
            exp_f := 0;
        ELSIF x =- 29180 THEN
            exp_f := 0;
        ELSIF x =- 29179 THEN
            exp_f := 0;
        ELSIF x =- 29178 THEN
            exp_f := 0;
        ELSIF x =- 29177 THEN
            exp_f := 0;
        ELSIF x =- 29176 THEN
            exp_f := 0;
        ELSIF x =- 29175 THEN
            exp_f := 0;
        ELSIF x =- 29174 THEN
            exp_f := 0;
        ELSIF x =- 29173 THEN
            exp_f := 0;
        ELSIF x =- 29172 THEN
            exp_f := 0;
        ELSIF x =- 29171 THEN
            exp_f := 0;
        ELSIF x =- 29170 THEN
            exp_f := 0;
        ELSIF x =- 29169 THEN
            exp_f := 0;
        ELSIF x =- 29168 THEN
            exp_f := 0;
        ELSIF x =- 29167 THEN
            exp_f := 0;
        ELSIF x =- 29166 THEN
            exp_f := 0;
        ELSIF x =- 29165 THEN
            exp_f := 0;
        ELSIF x =- 29164 THEN
            exp_f := 0;
        ELSIF x =- 29163 THEN
            exp_f := 0;
        ELSIF x =- 29162 THEN
            exp_f := 0;
        ELSIF x =- 29161 THEN
            exp_f := 0;
        ELSIF x =- 29160 THEN
            exp_f := 0;
        ELSIF x =- 29159 THEN
            exp_f := 0;
        ELSIF x =- 29158 THEN
            exp_f := 0;
        ELSIF x =- 29157 THEN
            exp_f := 0;
        ELSIF x =- 29156 THEN
            exp_f := 0;
        ELSIF x =- 29155 THEN
            exp_f := 0;
        ELSIF x =- 29154 THEN
            exp_f := 0;
        ELSIF x =- 29153 THEN
            exp_f := 0;
        ELSIF x =- 29152 THEN
            exp_f := 0;
        ELSIF x =- 29151 THEN
            exp_f := 0;
        ELSIF x =- 29150 THEN
            exp_f := 0;
        ELSIF x =- 29149 THEN
            exp_f := 0;
        ELSIF x =- 29148 THEN
            exp_f := 0;
        ELSIF x =- 29147 THEN
            exp_f := 0;
        ELSIF x =- 29146 THEN
            exp_f := 0;
        ELSIF x =- 29145 THEN
            exp_f := 0;
        ELSIF x =- 29144 THEN
            exp_f := 0;
        ELSIF x =- 29143 THEN
            exp_f := 0;
        ELSIF x =- 29142 THEN
            exp_f := 0;
        ELSIF x =- 29141 THEN
            exp_f := 0;
        ELSIF x =- 29140 THEN
            exp_f := 0;
        ELSIF x =- 29139 THEN
            exp_f := 0;
        ELSIF x =- 29138 THEN
            exp_f := 0;
        ELSIF x =- 29137 THEN
            exp_f := 0;
        ELSIF x =- 29136 THEN
            exp_f := 0;
        ELSIF x =- 29135 THEN
            exp_f := 0;
        ELSIF x =- 29134 THEN
            exp_f := 0;
        ELSIF x =- 29133 THEN
            exp_f := 0;
        ELSIF x =- 29132 THEN
            exp_f := 0;
        ELSIF x =- 29131 THEN
            exp_f := 0;
        ELSIF x =- 29130 THEN
            exp_f := 0;
        ELSIF x =- 29129 THEN
            exp_f := 0;
        ELSIF x =- 29128 THEN
            exp_f := 0;
        ELSIF x =- 29127 THEN
            exp_f := 0;
        ELSIF x =- 29126 THEN
            exp_f := 0;
        ELSIF x =- 29125 THEN
            exp_f := 0;
        ELSIF x =- 29124 THEN
            exp_f := 0;
        ELSIF x =- 29123 THEN
            exp_f := 0;
        ELSIF x =- 29122 THEN
            exp_f := 0;
        ELSIF x =- 29121 THEN
            exp_f := 0;
        ELSIF x =- 29120 THEN
            exp_f := 0;
        ELSIF x =- 29119 THEN
            exp_f := 0;
        ELSIF x =- 29118 THEN
            exp_f := 0;
        ELSIF x =- 29117 THEN
            exp_f := 0;
        ELSIF x =- 29116 THEN
            exp_f := 0;
        ELSIF x =- 29115 THEN
            exp_f := 0;
        ELSIF x =- 29114 THEN
            exp_f := 0;
        ELSIF x =- 29113 THEN
            exp_f := 0;
        ELSIF x =- 29112 THEN
            exp_f := 0;
        ELSIF x =- 29111 THEN
            exp_f := 0;
        ELSIF x =- 29110 THEN
            exp_f := 0;
        ELSIF x =- 29109 THEN
            exp_f := 0;
        ELSIF x =- 29108 THEN
            exp_f := 0;
        ELSIF x =- 29107 THEN
            exp_f := 0;
        ELSIF x =- 29106 THEN
            exp_f := 0;
        ELSIF x =- 29105 THEN
            exp_f := 0;
        ELSIF x =- 29104 THEN
            exp_f := 0;
        ELSIF x =- 29103 THEN
            exp_f := 0;
        ELSIF x =- 29102 THEN
            exp_f := 0;
        ELSIF x =- 29101 THEN
            exp_f := 0;
        ELSIF x =- 29100 THEN
            exp_f := 0;
        ELSIF x =- 29099 THEN
            exp_f := 0;
        ELSIF x =- 29098 THEN
            exp_f := 0;
        ELSIF x =- 29097 THEN
            exp_f := 0;
        ELSIF x =- 29096 THEN
            exp_f := 0;
        ELSIF x =- 29095 THEN
            exp_f := 0;
        ELSIF x =- 29094 THEN
            exp_f := 0;
        ELSIF x =- 29093 THEN
            exp_f := 0;
        ELSIF x =- 29092 THEN
            exp_f := 0;
        ELSIF x =- 29091 THEN
            exp_f := 0;
        ELSIF x =- 29090 THEN
            exp_f := 0;
        ELSIF x =- 29089 THEN
            exp_f := 0;
        ELSIF x =- 29088 THEN
            exp_f := 0;
        ELSIF x =- 29087 THEN
            exp_f := 0;
        ELSIF x =- 29086 THEN
            exp_f := 0;
        ELSIF x =- 29085 THEN
            exp_f := 0;
        ELSIF x =- 29084 THEN
            exp_f := 0;
        ELSIF x =- 29083 THEN
            exp_f := 0;
        ELSIF x =- 29082 THEN
            exp_f := 0;
        ELSIF x =- 29081 THEN
            exp_f := 0;
        ELSIF x =- 29080 THEN
            exp_f := 0;
        ELSIF x =- 29079 THEN
            exp_f := 0;
        ELSIF x =- 29078 THEN
            exp_f := 0;
        ELSIF x =- 29077 THEN
            exp_f := 0;
        ELSIF x =- 29076 THEN
            exp_f := 0;
        ELSIF x =- 29075 THEN
            exp_f := 0;
        ELSIF x =- 29074 THEN
            exp_f := 0;
        ELSIF x =- 29073 THEN
            exp_f := 0;
        ELSIF x =- 29072 THEN
            exp_f := 0;
        ELSIF x =- 29071 THEN
            exp_f := 0;
        ELSIF x =- 29070 THEN
            exp_f := 0;
        ELSIF x =- 29069 THEN
            exp_f := 0;
        ELSIF x =- 29068 THEN
            exp_f := 0;
        ELSIF x =- 29067 THEN
            exp_f := 0;
        ELSIF x =- 29066 THEN
            exp_f := 0;
        ELSIF x =- 29065 THEN
            exp_f := 0;
        ELSIF x =- 29064 THEN
            exp_f := 0;
        ELSIF x =- 29063 THEN
            exp_f := 0;
        ELSIF x =- 29062 THEN
            exp_f := 0;
        ELSIF x =- 29061 THEN
            exp_f := 0;
        ELSIF x =- 29060 THEN
            exp_f := 0;
        ELSIF x =- 29059 THEN
            exp_f := 0;
        ELSIF x =- 29058 THEN
            exp_f := 0;
        ELSIF x =- 29057 THEN
            exp_f := 0;
        ELSIF x =- 29056 THEN
            exp_f := 0;
        ELSIF x =- 29055 THEN
            exp_f := 0;
        ELSIF x =- 29054 THEN
            exp_f := 0;
        ELSIF x =- 29053 THEN
            exp_f := 0;
        ELSIF x =- 29052 THEN
            exp_f := 0;
        ELSIF x =- 29051 THEN
            exp_f := 0;
        ELSIF x =- 29050 THEN
            exp_f := 0;
        ELSIF x =- 29049 THEN
            exp_f := 0;
        ELSIF x =- 29048 THEN
            exp_f := 0;
        ELSIF x =- 29047 THEN
            exp_f := 0;
        ELSIF x =- 29046 THEN
            exp_f := 0;
        ELSIF x =- 29045 THEN
            exp_f := 0;
        ELSIF x =- 29044 THEN
            exp_f := 0;
        ELSIF x =- 29043 THEN
            exp_f := 0;
        ELSIF x =- 29042 THEN
            exp_f := 0;
        ELSIF x =- 29041 THEN
            exp_f := 0;
        ELSIF x =- 29040 THEN
            exp_f := 0;
        ELSIF x =- 29039 THEN
            exp_f := 0;
        ELSIF x =- 29038 THEN
            exp_f := 0;
        ELSIF x =- 29037 THEN
            exp_f := 0;
        ELSIF x =- 29036 THEN
            exp_f := 0;
        ELSIF x =- 29035 THEN
            exp_f := 0;
        ELSIF x =- 29034 THEN
            exp_f := 0;
        ELSIF x =- 29033 THEN
            exp_f := 0;
        ELSIF x =- 29032 THEN
            exp_f := 0;
        ELSIF x =- 29031 THEN
            exp_f := 0;
        ELSIF x =- 29030 THEN
            exp_f := 0;
        ELSIF x =- 29029 THEN
            exp_f := 0;
        ELSIF x =- 29028 THEN
            exp_f := 0;
        ELSIF x =- 29027 THEN
            exp_f := 0;
        ELSIF x =- 29026 THEN
            exp_f := 0;
        ELSIF x =- 29025 THEN
            exp_f := 0;
        ELSIF x =- 29024 THEN
            exp_f := 0;
        ELSIF x =- 29023 THEN
            exp_f := 0;
        ELSIF x =- 29022 THEN
            exp_f := 0;
        ELSIF x =- 29021 THEN
            exp_f := 0;
        ELSIF x =- 29020 THEN
            exp_f := 0;
        ELSIF x =- 29019 THEN
            exp_f := 0;
        ELSIF x =- 29018 THEN
            exp_f := 0;
        ELSIF x =- 29017 THEN
            exp_f := 0;
        ELSIF x =- 29016 THEN
            exp_f := 0;
        ELSIF x =- 29015 THEN
            exp_f := 0;
        ELSIF x =- 29014 THEN
            exp_f := 0;
        ELSIF x =- 29013 THEN
            exp_f := 0;
        ELSIF x =- 29012 THEN
            exp_f := 0;
        ELSIF x =- 29011 THEN
            exp_f := 0;
        ELSIF x =- 29010 THEN
            exp_f := 0;
        ELSIF x =- 29009 THEN
            exp_f := 0;
        ELSIF x =- 29008 THEN
            exp_f := 0;
        ELSIF x =- 29007 THEN
            exp_f := 0;
        ELSIF x =- 29006 THEN
            exp_f := 0;
        ELSIF x =- 29005 THEN
            exp_f := 0;
        ELSIF x =- 29004 THEN
            exp_f := 0;
        ELSIF x =- 29003 THEN
            exp_f := 0;
        ELSIF x =- 29002 THEN
            exp_f := 0;
        ELSIF x =- 29001 THEN
            exp_f := 0;
        ELSIF x =- 29000 THEN
            exp_f := 0;
        ELSIF x =- 28999 THEN
            exp_f := 0;
        ELSIF x =- 28998 THEN
            exp_f := 0;
        ELSIF x =- 28997 THEN
            exp_f := 0;
        ELSIF x =- 28996 THEN
            exp_f := 0;
        ELSIF x =- 28995 THEN
            exp_f := 0;
        ELSIF x =- 28994 THEN
            exp_f := 0;
        ELSIF x =- 28993 THEN
            exp_f := 0;
        ELSIF x =- 28992 THEN
            exp_f := 0;
        ELSIF x =- 28991 THEN
            exp_f := 0;
        ELSIF x =- 28990 THEN
            exp_f := 0;
        ELSIF x =- 28989 THEN
            exp_f := 0;
        ELSIF x =- 28988 THEN
            exp_f := 0;
        ELSIF x =- 28987 THEN
            exp_f := 0;
        ELSIF x =- 28986 THEN
            exp_f := 0;
        ELSIF x =- 28985 THEN
            exp_f := 0;
        ELSIF x =- 28984 THEN
            exp_f := 0;
        ELSIF x =- 28983 THEN
            exp_f := 0;
        ELSIF x =- 28982 THEN
            exp_f := 0;
        ELSIF x =- 28981 THEN
            exp_f := 0;
        ELSIF x =- 28980 THEN
            exp_f := 0;
        ELSIF x =- 28979 THEN
            exp_f := 0;
        ELSIF x =- 28978 THEN
            exp_f := 0;
        ELSIF x =- 28977 THEN
            exp_f := 0;
        ELSIF x =- 28976 THEN
            exp_f := 0;
        ELSIF x =- 28975 THEN
            exp_f := 0;
        ELSIF x =- 28974 THEN
            exp_f := 0;
        ELSIF x =- 28973 THEN
            exp_f := 0;
        ELSIF x =- 28972 THEN
            exp_f := 0;
        ELSIF x =- 28971 THEN
            exp_f := 0;
        ELSIF x =- 28970 THEN
            exp_f := 0;
        ELSIF x =- 28969 THEN
            exp_f := 0;
        ELSIF x =- 28968 THEN
            exp_f := 0;
        ELSIF x =- 28967 THEN
            exp_f := 0;
        ELSIF x =- 28966 THEN
            exp_f := 0;
        ELSIF x =- 28965 THEN
            exp_f := 0;
        ELSIF x =- 28964 THEN
            exp_f := 0;
        ELSIF x =- 28963 THEN
            exp_f := 0;
        ELSIF x =- 28962 THEN
            exp_f := 0;
        ELSIF x =- 28961 THEN
            exp_f := 0;
        ELSIF x =- 28960 THEN
            exp_f := 0;
        ELSIF x =- 28959 THEN
            exp_f := 0;
        ELSIF x =- 28958 THEN
            exp_f := 0;
        ELSIF x =- 28957 THEN
            exp_f := 0;
        ELSIF x =- 28956 THEN
            exp_f := 0;
        ELSIF x =- 28955 THEN
            exp_f := 0;
        ELSIF x =- 28954 THEN
            exp_f := 0;
        ELSIF x =- 28953 THEN
            exp_f := 0;
        ELSIF x =- 28952 THEN
            exp_f := 0;
        ELSIF x =- 28951 THEN
            exp_f := 0;
        ELSIF x =- 28950 THEN
            exp_f := 0;
        ELSIF x =- 28949 THEN
            exp_f := 0;
        ELSIF x =- 28948 THEN
            exp_f := 0;
        ELSIF x =- 28947 THEN
            exp_f := 0;
        ELSIF x =- 28946 THEN
            exp_f := 0;
        ELSIF x =- 28945 THEN
            exp_f := 0;
        ELSIF x =- 28944 THEN
            exp_f := 0;
        ELSIF x =- 28943 THEN
            exp_f := 0;
        ELSIF x =- 28942 THEN
            exp_f := 0;
        ELSIF x =- 28941 THEN
            exp_f := 0;
        ELSIF x =- 28940 THEN
            exp_f := 0;
        ELSIF x =- 28939 THEN
            exp_f := 0;
        ELSIF x =- 28938 THEN
            exp_f := 0;
        ELSIF x =- 28937 THEN
            exp_f := 0;
        ELSIF x =- 28936 THEN
            exp_f := 0;
        ELSIF x =- 28935 THEN
            exp_f := 0;
        ELSIF x =- 28934 THEN
            exp_f := 0;
        ELSIF x =- 28933 THEN
            exp_f := 0;
        ELSIF x =- 28932 THEN
            exp_f := 0;
        ELSIF x =- 28931 THEN
            exp_f := 0;
        ELSIF x =- 28930 THEN
            exp_f := 0;
        ELSIF x =- 28929 THEN
            exp_f := 0;
        ELSIF x =- 28928 THEN
            exp_f := 0;
        ELSIF x =- 28927 THEN
            exp_f := 0;
        ELSIF x =- 28926 THEN
            exp_f := 0;
        ELSIF x =- 28925 THEN
            exp_f := 0;
        ELSIF x =- 28924 THEN
            exp_f := 0;
        ELSIF x =- 28923 THEN
            exp_f := 0;
        ELSIF x =- 28922 THEN
            exp_f := 0;
        ELSIF x =- 28921 THEN
            exp_f := 0;
        ELSIF x =- 28920 THEN
            exp_f := 0;
        ELSIF x =- 28919 THEN
            exp_f := 0;
        ELSIF x =- 28918 THEN
            exp_f := 0;
        ELSIF x =- 28917 THEN
            exp_f := 0;
        ELSIF x =- 28916 THEN
            exp_f := 0;
        ELSIF x =- 28915 THEN
            exp_f := 0;
        ELSIF x =- 28914 THEN
            exp_f := 0;
        ELSIF x =- 28913 THEN
            exp_f := 0;
        ELSIF x =- 28912 THEN
            exp_f := 0;
        ELSIF x =- 28911 THEN
            exp_f := 0;
        ELSIF x =- 28910 THEN
            exp_f := 0;
        ELSIF x =- 28909 THEN
            exp_f := 0;
        ELSIF x =- 28908 THEN
            exp_f := 0;
        ELSIF x =- 28907 THEN
            exp_f := 0;
        ELSIF x =- 28906 THEN
            exp_f := 0;
        ELSIF x =- 28905 THEN
            exp_f := 0;
        ELSIF x =- 28904 THEN
            exp_f := 0;
        ELSIF x =- 28903 THEN
            exp_f := 0;
        ELSIF x =- 28902 THEN
            exp_f := 0;
        ELSIF x =- 28901 THEN
            exp_f := 0;
        ELSIF x =- 28900 THEN
            exp_f := 0;
        ELSIF x =- 28899 THEN
            exp_f := 0;
        ELSIF x =- 28898 THEN
            exp_f := 0;
        ELSIF x =- 28897 THEN
            exp_f := 0;
        ELSIF x =- 28896 THEN
            exp_f := 0;
        ELSIF x =- 28895 THEN
            exp_f := 0;
        ELSIF x =- 28894 THEN
            exp_f := 0;
        ELSIF x =- 28893 THEN
            exp_f := 0;
        ELSIF x =- 28892 THEN
            exp_f := 0;
        ELSIF x =- 28891 THEN
            exp_f := 0;
        ELSIF x =- 28890 THEN
            exp_f := 0;
        ELSIF x =- 28889 THEN
            exp_f := 0;
        ELSIF x =- 28888 THEN
            exp_f := 0;
        ELSIF x =- 28887 THEN
            exp_f := 0;
        ELSIF x =- 28886 THEN
            exp_f := 0;
        ELSIF x =- 28885 THEN
            exp_f := 0;
        ELSIF x =- 28884 THEN
            exp_f := 0;
        ELSIF x =- 28883 THEN
            exp_f := 0;
        ELSIF x =- 28882 THEN
            exp_f := 0;
        ELSIF x =- 28881 THEN
            exp_f := 0;
        ELSIF x =- 28880 THEN
            exp_f := 0;
        ELSIF x =- 28879 THEN
            exp_f := 0;
        ELSIF x =- 28878 THEN
            exp_f := 0;
        ELSIF x =- 28877 THEN
            exp_f := 0;
        ELSIF x =- 28876 THEN
            exp_f := 0;
        ELSIF x =- 28875 THEN
            exp_f := 0;
        ELSIF x =- 28874 THEN
            exp_f := 0;
        ELSIF x =- 28873 THEN
            exp_f := 0;
        ELSIF x =- 28872 THEN
            exp_f := 0;
        ELSIF x =- 28871 THEN
            exp_f := 0;
        ELSIF x =- 28870 THEN
            exp_f := 0;
        ELSIF x =- 28869 THEN
            exp_f := 0;
        ELSIF x =- 28868 THEN
            exp_f := 0;
        ELSIF x =- 28867 THEN
            exp_f := 0;
        ELSIF x =- 28866 THEN
            exp_f := 0;
        ELSIF x =- 28865 THEN
            exp_f := 0;
        ELSIF x =- 28864 THEN
            exp_f := 0;
        ELSIF x =- 28863 THEN
            exp_f := 0;
        ELSIF x =- 28862 THEN
            exp_f := 0;
        ELSIF x =- 28861 THEN
            exp_f := 0;
        ELSIF x =- 28860 THEN
            exp_f := 0;
        ELSIF x =- 28859 THEN
            exp_f := 0;
        ELSIF x =- 28858 THEN
            exp_f := 0;
        ELSIF x =- 28857 THEN
            exp_f := 0;
        ELSIF x =- 28856 THEN
            exp_f := 0;
        ELSIF x =- 28855 THEN
            exp_f := 0;
        ELSIF x =- 28854 THEN
            exp_f := 0;
        ELSIF x =- 28853 THEN
            exp_f := 0;
        ELSIF x =- 28852 THEN
            exp_f := 0;
        ELSIF x =- 28851 THEN
            exp_f := 0;
        ELSIF x =- 28850 THEN
            exp_f := 0;
        ELSIF x =- 28849 THEN
            exp_f := 0;
        ELSIF x =- 28848 THEN
            exp_f := 0;
        ELSIF x =- 28847 THEN
            exp_f := 0;
        ELSIF x =- 28846 THEN
            exp_f := 0;
        ELSIF x =- 28845 THEN
            exp_f := 0;
        ELSIF x =- 28844 THEN
            exp_f := 0;
        ELSIF x =- 28843 THEN
            exp_f := 0;
        ELSIF x =- 28842 THEN
            exp_f := 0;
        ELSIF x =- 28841 THEN
            exp_f := 0;
        ELSIF x =- 28840 THEN
            exp_f := 0;
        ELSIF x =- 28839 THEN
            exp_f := 0;
        ELSIF x =- 28838 THEN
            exp_f := 0;
        ELSIF x =- 28837 THEN
            exp_f := 0;
        ELSIF x =- 28836 THEN
            exp_f := 0;
        ELSIF x =- 28835 THEN
            exp_f := 0;
        ELSIF x =- 28834 THEN
            exp_f := 0;
        ELSIF x =- 28833 THEN
            exp_f := 0;
        ELSIF x =- 28832 THEN
            exp_f := 0;
        ELSIF x =- 28831 THEN
            exp_f := 0;
        ELSIF x =- 28830 THEN
            exp_f := 0;
        ELSIF x =- 28829 THEN
            exp_f := 0;
        ELSIF x =- 28828 THEN
            exp_f := 0;
        ELSIF x =- 28827 THEN
            exp_f := 0;
        ELSIF x =- 28826 THEN
            exp_f := 0;
        ELSIF x =- 28825 THEN
            exp_f := 0;
        ELSIF x =- 28824 THEN
            exp_f := 0;
        ELSIF x =- 28823 THEN
            exp_f := 0;
        ELSIF x =- 28822 THEN
            exp_f := 0;
        ELSIF x =- 28821 THEN
            exp_f := 0;
        ELSIF x =- 28820 THEN
            exp_f := 0;
        ELSIF x =- 28819 THEN
            exp_f := 0;
        ELSIF x =- 28818 THEN
            exp_f := 0;
        ELSIF x =- 28817 THEN
            exp_f := 0;
        ELSIF x =- 28816 THEN
            exp_f := 0;
        ELSIF x =- 28815 THEN
            exp_f := 0;
        ELSIF x =- 28814 THEN
            exp_f := 0;
        ELSIF x =- 28813 THEN
            exp_f := 0;
        ELSIF x =- 28812 THEN
            exp_f := 0;
        ELSIF x =- 28811 THEN
            exp_f := 0;
        ELSIF x =- 28810 THEN
            exp_f := 0;
        ELSIF x =- 28809 THEN
            exp_f := 0;
        ELSIF x =- 28808 THEN
            exp_f := 0;
        ELSIF x =- 28807 THEN
            exp_f := 0;
        ELSIF x =- 28806 THEN
            exp_f := 0;
        ELSIF x =- 28805 THEN
            exp_f := 0;
        ELSIF x =- 28804 THEN
            exp_f := 0;
        ELSIF x =- 28803 THEN
            exp_f := 0;
        ELSIF x =- 28802 THEN
            exp_f := 0;
        ELSIF x =- 28801 THEN
            exp_f := 0;
        ELSIF x =- 28800 THEN
            exp_f := 0;
        ELSIF x =- 28799 THEN
            exp_f := 0;
        ELSIF x =- 28798 THEN
            exp_f := 0;
        ELSIF x =- 28797 THEN
            exp_f := 0;
        ELSIF x =- 28796 THEN
            exp_f := 0;
        ELSIF x =- 28795 THEN
            exp_f := 0;
        ELSIF x =- 28794 THEN
            exp_f := 0;
        ELSIF x =- 28793 THEN
            exp_f := 0;
        ELSIF x =- 28792 THEN
            exp_f := 0;
        ELSIF x =- 28791 THEN
            exp_f := 0;
        ELSIF x =- 28790 THEN
            exp_f := 0;
        ELSIF x =- 28789 THEN
            exp_f := 0;
        ELSIF x =- 28788 THEN
            exp_f := 0;
        ELSIF x =- 28787 THEN
            exp_f := 0;
        ELSIF x =- 28786 THEN
            exp_f := 0;
        ELSIF x =- 28785 THEN
            exp_f := 0;
        ELSIF x =- 28784 THEN
            exp_f := 0;
        ELSIF x =- 28783 THEN
            exp_f := 0;
        ELSIF x =- 28782 THEN
            exp_f := 0;
        ELSIF x =- 28781 THEN
            exp_f := 0;
        ELSIF x =- 28780 THEN
            exp_f := 0;
        ELSIF x =- 28779 THEN
            exp_f := 0;
        ELSIF x =- 28778 THEN
            exp_f := 0;
        ELSIF x =- 28777 THEN
            exp_f := 0;
        ELSIF x =- 28776 THEN
            exp_f := 0;
        ELSIF x =- 28775 THEN
            exp_f := 0;
        ELSIF x =- 28774 THEN
            exp_f := 0;
        ELSIF x =- 28773 THEN
            exp_f := 0;
        ELSIF x =- 28772 THEN
            exp_f := 0;
        ELSIF x =- 28771 THEN
            exp_f := 0;
        ELSIF x =- 28770 THEN
            exp_f := 0;
        ELSIF x =- 28769 THEN
            exp_f := 0;
        ELSIF x =- 28768 THEN
            exp_f := 0;
        ELSIF x =- 28767 THEN
            exp_f := 0;
        ELSIF x =- 28766 THEN
            exp_f := 0;
        ELSIF x =- 28765 THEN
            exp_f := 0;
        ELSIF x =- 28764 THEN
            exp_f := 0;
        ELSIF x =- 28763 THEN
            exp_f := 0;
        ELSIF x =- 28762 THEN
            exp_f := 0;
        ELSIF x =- 28761 THEN
            exp_f := 0;
        ELSIF x =- 28760 THEN
            exp_f := 0;
        ELSIF x =- 28759 THEN
            exp_f := 0;
        ELSIF x =- 28758 THEN
            exp_f := 0;
        ELSIF x =- 28757 THEN
            exp_f := 0;
        ELSIF x =- 28756 THEN
            exp_f := 0;
        ELSIF x =- 28755 THEN
            exp_f := 0;
        ELSIF x =- 28754 THEN
            exp_f := 0;
        ELSIF x =- 28753 THEN
            exp_f := 0;
        ELSIF x =- 28752 THEN
            exp_f := 0;
        ELSIF x =- 28751 THEN
            exp_f := 0;
        ELSIF x =- 28750 THEN
            exp_f := 0;
        ELSIF x =- 28749 THEN
            exp_f := 0;
        ELSIF x =- 28748 THEN
            exp_f := 0;
        ELSIF x =- 28747 THEN
            exp_f := 0;
        ELSIF x =- 28746 THEN
            exp_f := 0;
        ELSIF x =- 28745 THEN
            exp_f := 0;
        ELSIF x =- 28744 THEN
            exp_f := 0;
        ELSIF x =- 28743 THEN
            exp_f := 0;
        ELSIF x =- 28742 THEN
            exp_f := 0;
        ELSIF x =- 28741 THEN
            exp_f := 0;
        ELSIF x =- 28740 THEN
            exp_f := 0;
        ELSIF x =- 28739 THEN
            exp_f := 0;
        ELSIF x =- 28738 THEN
            exp_f := 0;
        ELSIF x =- 28737 THEN
            exp_f := 0;
        ELSIF x =- 28736 THEN
            exp_f := 0;
        ELSIF x =- 28735 THEN
            exp_f := 0;
        ELSIF x =- 28734 THEN
            exp_f := 0;
        ELSIF x =- 28733 THEN
            exp_f := 0;
        ELSIF x =- 28732 THEN
            exp_f := 0;
        ELSIF x =- 28731 THEN
            exp_f := 0;
        ELSIF x =- 28730 THEN
            exp_f := 0;
        ELSIF x =- 28729 THEN
            exp_f := 0;
        ELSIF x =- 28728 THEN
            exp_f := 0;
        ELSIF x =- 28727 THEN
            exp_f := 0;
        ELSIF x =- 28726 THEN
            exp_f := 0;
        ELSIF x =- 28725 THEN
            exp_f := 0;
        ELSIF x =- 28724 THEN
            exp_f := 0;
        ELSIF x =- 28723 THEN
            exp_f := 0;
        ELSIF x =- 28722 THEN
            exp_f := 0;
        ELSIF x =- 28721 THEN
            exp_f := 0;
        ELSIF x =- 28720 THEN
            exp_f := 0;
        ELSIF x =- 28719 THEN
            exp_f := 0;
        ELSIF x =- 28718 THEN
            exp_f := 0;
        ELSIF x =- 28717 THEN
            exp_f := 0;
        ELSIF x =- 28716 THEN
            exp_f := 0;
        ELSIF x =- 28715 THEN
            exp_f := 0;
        ELSIF x =- 28714 THEN
            exp_f := 0;
        ELSIF x =- 28713 THEN
            exp_f := 0;
        ELSIF x =- 28712 THEN
            exp_f := 0;
        ELSIF x =- 28711 THEN
            exp_f := 0;
        ELSIF x =- 28710 THEN
            exp_f := 0;
        ELSIF x =- 28709 THEN
            exp_f := 0;
        ELSIF x =- 28708 THEN
            exp_f := 0;
        ELSIF x =- 28707 THEN
            exp_f := 0;
        ELSIF x =- 28706 THEN
            exp_f := 0;
        ELSIF x =- 28705 THEN
            exp_f := 0;
        ELSIF x =- 28704 THEN
            exp_f := 0;
        ELSIF x =- 28703 THEN
            exp_f := 0;
        ELSIF x =- 28702 THEN
            exp_f := 0;
        ELSIF x =- 28701 THEN
            exp_f := 0;
        ELSIF x =- 28700 THEN
            exp_f := 0;
        ELSIF x =- 28699 THEN
            exp_f := 0;
        ELSIF x =- 28698 THEN
            exp_f := 0;
        ELSIF x =- 28697 THEN
            exp_f := 0;
        ELSIF x =- 28696 THEN
            exp_f := 0;
        ELSIF x =- 28695 THEN
            exp_f := 0;
        ELSIF x =- 28694 THEN
            exp_f := 0;
        ELSIF x =- 28693 THEN
            exp_f := 0;
        ELSIF x =- 28692 THEN
            exp_f := 0;
        ELSIF x =- 28691 THEN
            exp_f := 0;
        ELSIF x =- 28690 THEN
            exp_f := 0;
        ELSIF x =- 28689 THEN
            exp_f := 0;
        ELSIF x =- 28688 THEN
            exp_f := 0;
        ELSIF x =- 28687 THEN
            exp_f := 0;
        ELSIF x =- 28686 THEN
            exp_f := 0;
        ELSIF x =- 28685 THEN
            exp_f := 0;
        ELSIF x =- 28684 THEN
            exp_f := 0;
        ELSIF x =- 28683 THEN
            exp_f := 0;
        ELSIF x =- 28682 THEN
            exp_f := 0;
        ELSIF x =- 28681 THEN
            exp_f := 0;
        ELSIF x =- 28680 THEN
            exp_f := 0;
        ELSIF x =- 28679 THEN
            exp_f := 0;
        ELSIF x =- 28678 THEN
            exp_f := 0;
        ELSIF x =- 28677 THEN
            exp_f := 0;
        ELSIF x =- 28676 THEN
            exp_f := 0;
        ELSIF x =- 28675 THEN
            exp_f := 0;
        ELSIF x =- 28674 THEN
            exp_f := 0;
        ELSIF x =- 28673 THEN
            exp_f := 0;
        ELSIF x =- 28672 THEN
            exp_f := 0;
        ELSIF x =- 28671 THEN
            exp_f := 0;
        ELSIF x =- 28670 THEN
            exp_f := 0;
        ELSIF x =- 28669 THEN
            exp_f := 0;
        ELSIF x =- 28668 THEN
            exp_f := 0;
        ELSIF x =- 28667 THEN
            exp_f := 0;
        ELSIF x =- 28666 THEN
            exp_f := 0;
        ELSIF x =- 28665 THEN
            exp_f := 0;
        ELSIF x =- 28664 THEN
            exp_f := 0;
        ELSIF x =- 28663 THEN
            exp_f := 0;
        ELSIF x =- 28662 THEN
            exp_f := 0;
        ELSIF x =- 28661 THEN
            exp_f := 0;
        ELSIF x =- 28660 THEN
            exp_f := 0;
        ELSIF x =- 28659 THEN
            exp_f := 0;
        ELSIF x =- 28658 THEN
            exp_f := 0;
        ELSIF x =- 28657 THEN
            exp_f := 0;
        ELSIF x =- 28656 THEN
            exp_f := 0;
        ELSIF x =- 28655 THEN
            exp_f := 0;
        ELSIF x =- 28654 THEN
            exp_f := 0;
        ELSIF x =- 28653 THEN
            exp_f := 0;
        ELSIF x =- 28652 THEN
            exp_f := 0;
        ELSIF x =- 28651 THEN
            exp_f := 0;
        ELSIF x =- 28650 THEN
            exp_f := 0;
        ELSIF x =- 28649 THEN
            exp_f := 0;
        ELSIF x =- 28648 THEN
            exp_f := 0;
        ELSIF x =- 28647 THEN
            exp_f := 0;
        ELSIF x =- 28646 THEN
            exp_f := 0;
        ELSIF x =- 28645 THEN
            exp_f := 0;
        ELSIF x =- 28644 THEN
            exp_f := 0;
        ELSIF x =- 28643 THEN
            exp_f := 0;
        ELSIF x =- 28642 THEN
            exp_f := 0;
        ELSIF x =- 28641 THEN
            exp_f := 0;
        ELSIF x =- 28640 THEN
            exp_f := 0;
        ELSIF x =- 28639 THEN
            exp_f := 0;
        ELSIF x =- 28638 THEN
            exp_f := 0;
        ELSIF x =- 28637 THEN
            exp_f := 0;
        ELSIF x =- 28636 THEN
            exp_f := 0;
        ELSIF x =- 28635 THEN
            exp_f := 0;
        ELSIF x =- 28634 THEN
            exp_f := 0;
        ELSIF x =- 28633 THEN
            exp_f := 0;
        ELSIF x =- 28632 THEN
            exp_f := 0;
        ELSIF x =- 28631 THEN
            exp_f := 0;
        ELSIF x =- 28630 THEN
            exp_f := 0;
        ELSIF x =- 28629 THEN
            exp_f := 0;
        ELSIF x =- 28628 THEN
            exp_f := 0;
        ELSIF x =- 28627 THEN
            exp_f := 0;
        ELSIF x =- 28626 THEN
            exp_f := 0;
        ELSIF x =- 28625 THEN
            exp_f := 0;
        ELSIF x =- 28624 THEN
            exp_f := 0;
        ELSIF x =- 28623 THEN
            exp_f := 0;
        ELSIF x =- 28622 THEN
            exp_f := 0;
        ELSIF x =- 28621 THEN
            exp_f := 0;
        ELSIF x =- 28620 THEN
            exp_f := 0;
        ELSIF x =- 28619 THEN
            exp_f := 0;
        ELSIF x =- 28618 THEN
            exp_f := 0;
        ELSIF x =- 28617 THEN
            exp_f := 0;
        ELSIF x =- 28616 THEN
            exp_f := 0;
        ELSIF x =- 28615 THEN
            exp_f := 0;
        ELSIF x =- 28614 THEN
            exp_f := 0;
        ELSIF x =- 28613 THEN
            exp_f := 0;
        ELSIF x =- 28612 THEN
            exp_f := 0;
        ELSIF x =- 28611 THEN
            exp_f := 0;
        ELSIF x =- 28610 THEN
            exp_f := 0;
        ELSIF x =- 28609 THEN
            exp_f := 0;
        ELSIF x =- 28608 THEN
            exp_f := 0;
        ELSIF x =- 28607 THEN
            exp_f := 0;
        ELSIF x =- 28606 THEN
            exp_f := 0;
        ELSIF x =- 28605 THEN
            exp_f := 0;
        ELSIF x =- 28604 THEN
            exp_f := 0;
        ELSIF x =- 28603 THEN
            exp_f := 0;
        ELSIF x =- 28602 THEN
            exp_f := 0;
        ELSIF x =- 28601 THEN
            exp_f := 0;
        ELSIF x =- 28600 THEN
            exp_f := 0;
        ELSIF x =- 28599 THEN
            exp_f := 0;
        ELSIF x =- 28598 THEN
            exp_f := 0;
        ELSIF x =- 28597 THEN
            exp_f := 0;
        ELSIF x =- 28596 THEN
            exp_f := 0;
        ELSIF x =- 28595 THEN
            exp_f := 0;
        ELSIF x =- 28594 THEN
            exp_f := 0;
        ELSIF x =- 28593 THEN
            exp_f := 0;
        ELSIF x =- 28592 THEN
            exp_f := 0;
        ELSIF x =- 28591 THEN
            exp_f := 0;
        ELSIF x =- 28590 THEN
            exp_f := 0;
        ELSIF x =- 28589 THEN
            exp_f := 0;
        ELSIF x =- 28588 THEN
            exp_f := 0;
        ELSIF x =- 28587 THEN
            exp_f := 0;
        ELSIF x =- 28586 THEN
            exp_f := 0;
        ELSIF x =- 28585 THEN
            exp_f := 0;
        ELSIF x =- 28584 THEN
            exp_f := 0;
        ELSIF x =- 28583 THEN
            exp_f := 0;
        ELSIF x =- 28582 THEN
            exp_f := 0;
        ELSIF x =- 28581 THEN
            exp_f := 0;
        ELSIF x =- 28580 THEN
            exp_f := 0;
        ELSIF x =- 28579 THEN
            exp_f := 0;
        ELSIF x =- 28578 THEN
            exp_f := 0;
        ELSIF x =- 28577 THEN
            exp_f := 0;
        ELSIF x =- 28576 THEN
            exp_f := 0;
        ELSIF x =- 28575 THEN
            exp_f := 0;
        ELSIF x =- 28574 THEN
            exp_f := 0;
        ELSIF x =- 28573 THEN
            exp_f := 0;
        ELSIF x =- 28572 THEN
            exp_f := 0;
        ELSIF x =- 28571 THEN
            exp_f := 0;
        ELSIF x =- 28570 THEN
            exp_f := 0;
        ELSIF x =- 28569 THEN
            exp_f := 0;
        ELSIF x =- 28568 THEN
            exp_f := 0;
        ELSIF x =- 28567 THEN
            exp_f := 0;
        ELSIF x =- 28566 THEN
            exp_f := 0;
        ELSIF x =- 28565 THEN
            exp_f := 0;
        ELSIF x =- 28564 THEN
            exp_f := 0;
        ELSIF x =- 28563 THEN
            exp_f := 0;
        ELSIF x =- 28562 THEN
            exp_f := 0;
        ELSIF x =- 28561 THEN
            exp_f := 0;
        ELSIF x =- 28560 THEN
            exp_f := 0;
        ELSIF x =- 28559 THEN
            exp_f := 0;
        ELSIF x =- 28558 THEN
            exp_f := 0;
        ELSIF x =- 28557 THEN
            exp_f := 0;
        ELSIF x =- 28556 THEN
            exp_f := 0;
        ELSIF x =- 28555 THEN
            exp_f := 0;
        ELSIF x =- 28554 THEN
            exp_f := 0;
        ELSIF x =- 28553 THEN
            exp_f := 0;
        ELSIF x =- 28552 THEN
            exp_f := 0;
        ELSIF x =- 28551 THEN
            exp_f := 0;
        ELSIF x =- 28550 THEN
            exp_f := 0;
        ELSIF x =- 28549 THEN
            exp_f := 0;
        ELSIF x =- 28548 THEN
            exp_f := 0;
        ELSIF x =- 28547 THEN
            exp_f := 0;
        ELSIF x =- 28546 THEN
            exp_f := 0;
        ELSIF x =- 28545 THEN
            exp_f := 0;
        ELSIF x =- 28544 THEN
            exp_f := 0;
        ELSIF x =- 28543 THEN
            exp_f := 0;
        ELSIF x =- 28542 THEN
            exp_f := 0;
        ELSIF x =- 28541 THEN
            exp_f := 0;
        ELSIF x =- 28540 THEN
            exp_f := 0;
        ELSIF x =- 28539 THEN
            exp_f := 0;
        ELSIF x =- 28538 THEN
            exp_f := 0;
        ELSIF x =- 28537 THEN
            exp_f := 0;
        ELSIF x =- 28536 THEN
            exp_f := 0;
        ELSIF x =- 28535 THEN
            exp_f := 0;
        ELSIF x =- 28534 THEN
            exp_f := 0;
        ELSIF x =- 28533 THEN
            exp_f := 0;
        ELSIF x =- 28532 THEN
            exp_f := 0;
        ELSIF x =- 28531 THEN
            exp_f := 0;
        ELSIF x =- 28530 THEN
            exp_f := 0;
        ELSIF x =- 28529 THEN
            exp_f := 0;
        ELSIF x =- 28528 THEN
            exp_f := 0;
        ELSIF x =- 28527 THEN
            exp_f := 0;
        ELSIF x =- 28526 THEN
            exp_f := 0;
        ELSIF x =- 28525 THEN
            exp_f := 0;
        ELSIF x =- 28524 THEN
            exp_f := 0;
        ELSIF x =- 28523 THEN
            exp_f := 0;
        ELSIF x =- 28522 THEN
            exp_f := 0;
        ELSIF x =- 28521 THEN
            exp_f := 0;
        ELSIF x =- 28520 THEN
            exp_f := 0;
        ELSIF x =- 28519 THEN
            exp_f := 0;
        ELSIF x =- 28518 THEN
            exp_f := 0;
        ELSIF x =- 28517 THEN
            exp_f := 0;
        ELSIF x =- 28516 THEN
            exp_f := 0;
        ELSIF x =- 28515 THEN
            exp_f := 0;
        ELSIF x =- 28514 THEN
            exp_f := 0;
        ELSIF x =- 28513 THEN
            exp_f := 0;
        ELSIF x =- 28512 THEN
            exp_f := 0;
        ELSIF x =- 28511 THEN
            exp_f := 0;
        ELSIF x =- 28510 THEN
            exp_f := 0;
        ELSIF x =- 28509 THEN
            exp_f := 0;
        ELSIF x =- 28508 THEN
            exp_f := 0;
        ELSIF x =- 28507 THEN
            exp_f := 0;
        ELSIF x =- 28506 THEN
            exp_f := 0;
        ELSIF x =- 28505 THEN
            exp_f := 0;
        ELSIF x =- 28504 THEN
            exp_f := 0;
        ELSIF x =- 28503 THEN
            exp_f := 0;
        ELSIF x =- 28502 THEN
            exp_f := 0;
        ELSIF x =- 28501 THEN
            exp_f := 0;
        ELSIF x =- 28500 THEN
            exp_f := 0;
        ELSIF x =- 28499 THEN
            exp_f := 0;
        ELSIF x =- 28498 THEN
            exp_f := 0;
        ELSIF x =- 28497 THEN
            exp_f := 0;
        ELSIF x =- 28496 THEN
            exp_f := 0;
        ELSIF x =- 28495 THEN
            exp_f := 0;
        ELSIF x =- 28494 THEN
            exp_f := 0;
        ELSIF x =- 28493 THEN
            exp_f := 0;
        ELSIF x =- 28492 THEN
            exp_f := 0;
        ELSIF x =- 28491 THEN
            exp_f := 0;
        ELSIF x =- 28490 THEN
            exp_f := 0;
        ELSIF x =- 28489 THEN
            exp_f := 0;
        ELSIF x =- 28488 THEN
            exp_f := 0;
        ELSIF x =- 28487 THEN
            exp_f := 0;
        ELSIF x =- 28486 THEN
            exp_f := 0;
        ELSIF x =- 28485 THEN
            exp_f := 0;
        ELSIF x =- 28484 THEN
            exp_f := 0;
        ELSIF x =- 28483 THEN
            exp_f := 0;
        ELSIF x =- 28482 THEN
            exp_f := 0;
        ELSIF x =- 28481 THEN
            exp_f := 0;
        ELSIF x =- 28480 THEN
            exp_f := 0;
        ELSIF x =- 28479 THEN
            exp_f := 0;
        ELSIF x =- 28478 THEN
            exp_f := 0;
        ELSIF x =- 28477 THEN
            exp_f := 0;
        ELSIF x =- 28476 THEN
            exp_f := 0;
        ELSIF x =- 28475 THEN
            exp_f := 0;
        ELSIF x =- 28474 THEN
            exp_f := 0;
        ELSIF x =- 28473 THEN
            exp_f := 0;
        ELSIF x =- 28472 THEN
            exp_f := 0;
        ELSIF x =- 28471 THEN
            exp_f := 0;
        ELSIF x =- 28470 THEN
            exp_f := 0;
        ELSIF x =- 28469 THEN
            exp_f := 0;
        ELSIF x =- 28468 THEN
            exp_f := 0;
        ELSIF x =- 28467 THEN
            exp_f := 0;
        ELSIF x =- 28466 THEN
            exp_f := 0;
        ELSIF x =- 28465 THEN
            exp_f := 0;
        ELSIF x =- 28464 THEN
            exp_f := 0;
        ELSIF x =- 28463 THEN
            exp_f := 0;
        ELSIF x =- 28462 THEN
            exp_f := 0;
        ELSIF x =- 28461 THEN
            exp_f := 0;
        ELSIF x =- 28460 THEN
            exp_f := 0;
        ELSIF x =- 28459 THEN
            exp_f := 0;
        ELSIF x =- 28458 THEN
            exp_f := 0;
        ELSIF x =- 28457 THEN
            exp_f := 0;
        ELSIF x =- 28456 THEN
            exp_f := 0;
        ELSIF x =- 28455 THEN
            exp_f := 0;
        ELSIF x =- 28454 THEN
            exp_f := 0;
        ELSIF x =- 28453 THEN
            exp_f := 0;
        ELSIF x =- 28452 THEN
            exp_f := 0;
        ELSIF x =- 28451 THEN
            exp_f := 0;
        ELSIF x =- 28450 THEN
            exp_f := 0;
        ELSIF x =- 28449 THEN
            exp_f := 0;
        ELSIF x =- 28448 THEN
            exp_f := 0;
        ELSIF x =- 28447 THEN
            exp_f := 0;
        ELSIF x =- 28446 THEN
            exp_f := 0;
        ELSIF x =- 28445 THEN
            exp_f := 0;
        ELSIF x =- 28444 THEN
            exp_f := 0;
        ELSIF x =- 28443 THEN
            exp_f := 0;
        ELSIF x =- 28442 THEN
            exp_f := 0;
        ELSIF x =- 28441 THEN
            exp_f := 0;
        ELSIF x =- 28440 THEN
            exp_f := 0;
        ELSIF x =- 28439 THEN
            exp_f := 0;
        ELSIF x =- 28438 THEN
            exp_f := 0;
        ELSIF x =- 28437 THEN
            exp_f := 0;
        ELSIF x =- 28436 THEN
            exp_f := 0;
        ELSIF x =- 28435 THEN
            exp_f := 0;
        ELSIF x =- 28434 THEN
            exp_f := 0;
        ELSIF x =- 28433 THEN
            exp_f := 0;
        ELSIF x =- 28432 THEN
            exp_f := 0;
        ELSIF x =- 28431 THEN
            exp_f := 0;
        ELSIF x =- 28430 THEN
            exp_f := 0;
        ELSIF x =- 28429 THEN
            exp_f := 0;
        ELSIF x =- 28428 THEN
            exp_f := 0;
        ELSIF x =- 28427 THEN
            exp_f := 0;
        ELSIF x =- 28426 THEN
            exp_f := 0;
        ELSIF x =- 28425 THEN
            exp_f := 0;
        ELSIF x =- 28424 THEN
            exp_f := 0;
        ELSIF x =- 28423 THEN
            exp_f := 0;
        ELSIF x =- 28422 THEN
            exp_f := 0;
        ELSIF x =- 28421 THEN
            exp_f := 0;
        ELSIF x =- 28420 THEN
            exp_f := 0;
        ELSIF x =- 28419 THEN
            exp_f := 0;
        ELSIF x =- 28418 THEN
            exp_f := 0;
        ELSIF x =- 28417 THEN
            exp_f := 0;
        ELSIF x =- 28416 THEN
            exp_f := 0;
        ELSIF x =- 28415 THEN
            exp_f := 0;
        ELSIF x =- 28414 THEN
            exp_f := 0;
        ELSIF x =- 28413 THEN
            exp_f := 0;
        ELSIF x =- 28412 THEN
            exp_f := 0;
        ELSIF x =- 28411 THEN
            exp_f := 0;
        ELSIF x =- 28410 THEN
            exp_f := 0;
        ELSIF x =- 28409 THEN
            exp_f := 0;
        ELSIF x =- 28408 THEN
            exp_f := 0;
        ELSIF x =- 28407 THEN
            exp_f := 0;
        ELSIF x =- 28406 THEN
            exp_f := 0;
        ELSIF x =- 28405 THEN
            exp_f := 0;
        ELSIF x =- 28404 THEN
            exp_f := 0;
        ELSIF x =- 28403 THEN
            exp_f := 0;
        ELSIF x =- 28402 THEN
            exp_f := 0;
        ELSIF x =- 28401 THEN
            exp_f := 0;
        ELSIF x =- 28400 THEN
            exp_f := 0;
        ELSIF x =- 28399 THEN
            exp_f := 0;
        ELSIF x =- 28398 THEN
            exp_f := 0;
        ELSIF x =- 28397 THEN
            exp_f := 0;
        ELSIF x =- 28396 THEN
            exp_f := 0;
        ELSIF x =- 28395 THEN
            exp_f := 0;
        ELSIF x =- 28394 THEN
            exp_f := 0;
        ELSIF x =- 28393 THEN
            exp_f := 0;
        ELSIF x =- 28392 THEN
            exp_f := 0;
        ELSIF x =- 28391 THEN
            exp_f := 0;
        ELSIF x =- 28390 THEN
            exp_f := 0;
        ELSIF x =- 28389 THEN
            exp_f := 0;
        ELSIF x =- 28388 THEN
            exp_f := 0;
        ELSIF x =- 28387 THEN
            exp_f := 0;
        ELSIF x =- 28386 THEN
            exp_f := 0;
        ELSIF x =- 28385 THEN
            exp_f := 0;
        ELSIF x =- 28384 THEN
            exp_f := 0;
        ELSIF x =- 28383 THEN
            exp_f := 0;
        ELSIF x =- 28382 THEN
            exp_f := 0;
        ELSIF x =- 28381 THEN
            exp_f := 0;
        ELSIF x =- 28380 THEN
            exp_f := 0;
        ELSIF x =- 28379 THEN
            exp_f := 0;
        ELSIF x =- 28378 THEN
            exp_f := 0;
        ELSIF x =- 28377 THEN
            exp_f := 0;
        ELSIF x =- 28376 THEN
            exp_f := 0;
        ELSIF x =- 28375 THEN
            exp_f := 0;
        ELSIF x =- 28374 THEN
            exp_f := 0;
        ELSIF x =- 28373 THEN
            exp_f := 0;
        ELSIF x =- 28372 THEN
            exp_f := 0;
        ELSIF x =- 28371 THEN
            exp_f := 0;
        ELSIF x =- 28370 THEN
            exp_f := 0;
        ELSIF x =- 28369 THEN
            exp_f := 0;
        ELSIF x =- 28368 THEN
            exp_f := 0;
        ELSIF x =- 28367 THEN
            exp_f := 0;
        ELSIF x =- 28366 THEN
            exp_f := 0;
        ELSIF x =- 28365 THEN
            exp_f := 0;
        ELSIF x =- 28364 THEN
            exp_f := 0;
        ELSIF x =- 28363 THEN
            exp_f := 0;
        ELSIF x =- 28362 THEN
            exp_f := 0;
        ELSIF x =- 28361 THEN
            exp_f := 0;
        ELSIF x =- 28360 THEN
            exp_f := 0;
        ELSIF x =- 28359 THEN
            exp_f := 0;
        ELSIF x =- 28358 THEN
            exp_f := 0;
        ELSIF x =- 28357 THEN
            exp_f := 0;
        ELSIF x =- 28356 THEN
            exp_f := 0;
        ELSIF x =- 28355 THEN
            exp_f := 0;
        ELSIF x =- 28354 THEN
            exp_f := 0;
        ELSIF x =- 28353 THEN
            exp_f := 0;
        ELSIF x =- 28352 THEN
            exp_f := 0;
        ELSIF x =- 28351 THEN
            exp_f := 0;
        ELSIF x =- 28350 THEN
            exp_f := 0;
        ELSIF x =- 28349 THEN
            exp_f := 0;
        ELSIF x =- 28348 THEN
            exp_f := 0;
        ELSIF x =- 28347 THEN
            exp_f := 0;
        ELSIF x =- 28346 THEN
            exp_f := 0;
        ELSIF x =- 28345 THEN
            exp_f := 0;
        ELSIF x =- 28344 THEN
            exp_f := 0;
        ELSIF x =- 28343 THEN
            exp_f := 0;
        ELSIF x =- 28342 THEN
            exp_f := 0;
        ELSIF x =- 28341 THEN
            exp_f := 0;
        ELSIF x =- 28340 THEN
            exp_f := 0;
        ELSIF x =- 28339 THEN
            exp_f := 0;
        ELSIF x =- 28338 THEN
            exp_f := 0;
        ELSIF x =- 28337 THEN
            exp_f := 0;
        ELSIF x =- 28336 THEN
            exp_f := 0;
        ELSIF x =- 28335 THEN
            exp_f := 0;
        ELSIF x =- 28334 THEN
            exp_f := 0;
        ELSIF x =- 28333 THEN
            exp_f := 0;
        ELSIF x =- 28332 THEN
            exp_f := 0;
        ELSIF x =- 28331 THEN
            exp_f := 0;
        ELSIF x =- 28330 THEN
            exp_f := 0;
        ELSIF x =- 28329 THEN
            exp_f := 0;
        ELSIF x =- 28328 THEN
            exp_f := 0;
        ELSIF x =- 28327 THEN
            exp_f := 0;
        ELSIF x =- 28326 THEN
            exp_f := 0;
        ELSIF x =- 28325 THEN
            exp_f := 0;
        ELSIF x =- 28324 THEN
            exp_f := 0;
        ELSIF x =- 28323 THEN
            exp_f := 0;
        ELSIF x =- 28322 THEN
            exp_f := 0;
        ELSIF x =- 28321 THEN
            exp_f := 0;
        ELSIF x =- 28320 THEN
            exp_f := 0;
        ELSIF x =- 28319 THEN
            exp_f := 0;
        ELSIF x =- 28318 THEN
            exp_f := 0;
        ELSIF x =- 28317 THEN
            exp_f := 0;
        ELSIF x =- 28316 THEN
            exp_f := 0;
        ELSIF x =- 28315 THEN
            exp_f := 0;
        ELSIF x =- 28314 THEN
            exp_f := 0;
        ELSIF x =- 28313 THEN
            exp_f := 0;
        ELSIF x =- 28312 THEN
            exp_f := 0;
        ELSIF x =- 28311 THEN
            exp_f := 0;
        ELSIF x =- 28310 THEN
            exp_f := 0;
        ELSIF x =- 28309 THEN
            exp_f := 0;
        ELSIF x =- 28308 THEN
            exp_f := 0;
        ELSIF x =- 28307 THEN
            exp_f := 0;
        ELSIF x =- 28306 THEN
            exp_f := 0;
        ELSIF x =- 28305 THEN
            exp_f := 0;
        ELSIF x =- 28304 THEN
            exp_f := 0;
        ELSIF x =- 28303 THEN
            exp_f := 0;
        ELSIF x =- 28302 THEN
            exp_f := 0;
        ELSIF x =- 28301 THEN
            exp_f := 0;
        ELSIF x =- 28300 THEN
            exp_f := 0;
        ELSIF x =- 28299 THEN
            exp_f := 0;
        ELSIF x =- 28298 THEN
            exp_f := 0;
        ELSIF x =- 28297 THEN
            exp_f := 0;
        ELSIF x =- 28296 THEN
            exp_f := 0;
        ELSIF x =- 28295 THEN
            exp_f := 0;
        ELSIF x =- 28294 THEN
            exp_f := 0;
        ELSIF x =- 28293 THEN
            exp_f := 0;
        ELSIF x =- 28292 THEN
            exp_f := 0;
        ELSIF x =- 28291 THEN
            exp_f := 0;
        ELSIF x =- 28290 THEN
            exp_f := 0;
        ELSIF x =- 28289 THEN
            exp_f := 0;
        ELSIF x =- 28288 THEN
            exp_f := 0;
        ELSIF x =- 28287 THEN
            exp_f := 0;
        ELSIF x =- 28286 THEN
            exp_f := 0;
        ELSIF x =- 28285 THEN
            exp_f := 0;
        ELSIF x =- 28284 THEN
            exp_f := 0;
        ELSIF x =- 28283 THEN
            exp_f := 0;
        ELSIF x =- 28282 THEN
            exp_f := 0;
        ELSIF x =- 28281 THEN
            exp_f := 0;
        ELSIF x =- 28280 THEN
            exp_f := 0;
        ELSIF x =- 28279 THEN
            exp_f := 0;
        ELSIF x =- 28278 THEN
            exp_f := 0;
        ELSIF x =- 28277 THEN
            exp_f := 0;
        ELSIF x =- 28276 THEN
            exp_f := 0;
        ELSIF x =- 28275 THEN
            exp_f := 0;
        ELSIF x =- 28274 THEN
            exp_f := 0;
        ELSIF x =- 28273 THEN
            exp_f := 0;
        ELSIF x =- 28272 THEN
            exp_f := 0;
        ELSIF x =- 28271 THEN
            exp_f := 0;
        ELSIF x =- 28270 THEN
            exp_f := 0;
        ELSIF x =- 28269 THEN
            exp_f := 0;
        ELSIF x =- 28268 THEN
            exp_f := 0;
        ELSIF x =- 28267 THEN
            exp_f := 0;
        ELSIF x =- 28266 THEN
            exp_f := 0;
        ELSIF x =- 28265 THEN
            exp_f := 0;
        ELSIF x =- 28264 THEN
            exp_f := 0;
        ELSIF x =- 28263 THEN
            exp_f := 0;
        ELSIF x =- 28262 THEN
            exp_f := 0;
        ELSIF x =- 28261 THEN
            exp_f := 0;
        ELSIF x =- 28260 THEN
            exp_f := 0;
        ELSIF x =- 28259 THEN
            exp_f := 0;
        ELSIF x =- 28258 THEN
            exp_f := 0;
        ELSIF x =- 28257 THEN
            exp_f := 0;
        ELSIF x =- 28256 THEN
            exp_f := 0;
        ELSIF x =- 28255 THEN
            exp_f := 0;
        ELSIF x =- 28254 THEN
            exp_f := 0;
        ELSIF x =- 28253 THEN
            exp_f := 0;
        ELSIF x =- 28252 THEN
            exp_f := 0;
        ELSIF x =- 28251 THEN
            exp_f := 0;
        ELSIF x =- 28250 THEN
            exp_f := 0;
        ELSIF x =- 28249 THEN
            exp_f := 0;
        ELSIF x =- 28248 THEN
            exp_f := 0;
        ELSIF x =- 28247 THEN
            exp_f := 0;
        ELSIF x =- 28246 THEN
            exp_f := 0;
        ELSIF x =- 28245 THEN
            exp_f := 0;
        ELSIF x =- 28244 THEN
            exp_f := 0;
        ELSIF x =- 28243 THEN
            exp_f := 0;
        ELSIF x =- 28242 THEN
            exp_f := 0;
        ELSIF x =- 28241 THEN
            exp_f := 0;
        ELSIF x =- 28240 THEN
            exp_f := 0;
        ELSIF x =- 28239 THEN
            exp_f := 0;
        ELSIF x =- 28238 THEN
            exp_f := 0;
        ELSIF x =- 28237 THEN
            exp_f := 0;
        ELSIF x =- 28236 THEN
            exp_f := 0;
        ELSIF x =- 28235 THEN
            exp_f := 0;
        ELSIF x =- 28234 THEN
            exp_f := 0;
        ELSIF x =- 28233 THEN
            exp_f := 0;
        ELSIF x =- 28232 THEN
            exp_f := 0;
        ELSIF x =- 28231 THEN
            exp_f := 0;
        ELSIF x =- 28230 THEN
            exp_f := 0;
        ELSIF x =- 28229 THEN
            exp_f := 0;
        ELSIF x =- 28228 THEN
            exp_f := 0;
        ELSIF x =- 28227 THEN
            exp_f := 0;
        ELSIF x =- 28226 THEN
            exp_f := 0;
        ELSIF x =- 28225 THEN
            exp_f := 0;
        ELSIF x =- 28224 THEN
            exp_f := 0;
        ELSIF x =- 28223 THEN
            exp_f := 0;
        ELSIF x =- 28222 THEN
            exp_f := 0;
        ELSIF x =- 28221 THEN
            exp_f := 0;
        ELSIF x =- 28220 THEN
            exp_f := 0;
        ELSIF x =- 28219 THEN
            exp_f := 0;
        ELSIF x =- 28218 THEN
            exp_f := 0;
        ELSIF x =- 28217 THEN
            exp_f := 0;
        ELSIF x =- 28216 THEN
            exp_f := 0;
        ELSIF x =- 28215 THEN
            exp_f := 0;
        ELSIF x =- 28214 THEN
            exp_f := 0;
        ELSIF x =- 28213 THEN
            exp_f := 0;
        ELSIF x =- 28212 THEN
            exp_f := 0;
        ELSIF x =- 28211 THEN
            exp_f := 0;
        ELSIF x =- 28210 THEN
            exp_f := 0;
        ELSIF x =- 28209 THEN
            exp_f := 0;
        ELSIF x =- 28208 THEN
            exp_f := 0;
        ELSIF x =- 28207 THEN
            exp_f := 0;
        ELSIF x =- 28206 THEN
            exp_f := 0;
        ELSIF x =- 28205 THEN
            exp_f := 0;
        ELSIF x =- 28204 THEN
            exp_f := 0;
        ELSIF x =- 28203 THEN
            exp_f := 0;
        ELSIF x =- 28202 THEN
            exp_f := 0;
        ELSIF x =- 28201 THEN
            exp_f := 0;
        ELSIF x =- 28200 THEN
            exp_f := 0;
        ELSIF x =- 28199 THEN
            exp_f := 0;
        ELSIF x =- 28198 THEN
            exp_f := 0;
        ELSIF x =- 28197 THEN
            exp_f := 0;
        ELSIF x =- 28196 THEN
            exp_f := 0;
        ELSIF x =- 28195 THEN
            exp_f := 0;
        ELSIF x =- 28194 THEN
            exp_f := 0;
        ELSIF x =- 28193 THEN
            exp_f := 0;
        ELSIF x =- 28192 THEN
            exp_f := 0;
        ELSIF x =- 28191 THEN
            exp_f := 0;
        ELSIF x =- 28190 THEN
            exp_f := 0;
        ELSIF x =- 28189 THEN
            exp_f := 0;
        ELSIF x =- 28188 THEN
            exp_f := 0;
        ELSIF x =- 28187 THEN
            exp_f := 0;
        ELSIF x =- 28186 THEN
            exp_f := 0;
        ELSIF x =- 28185 THEN
            exp_f := 0;
        ELSIF x =- 28184 THEN
            exp_f := 0;
        ELSIF x =- 28183 THEN
            exp_f := 0;
        ELSIF x =- 28182 THEN
            exp_f := 0;
        ELSIF x =- 28181 THEN
            exp_f := 0;
        ELSIF x =- 28180 THEN
            exp_f := 0;
        ELSIF x =- 28179 THEN
            exp_f := 0;
        ELSIF x =- 28178 THEN
            exp_f := 0;
        ELSIF x =- 28177 THEN
            exp_f := 0;
        ELSIF x =- 28176 THEN
            exp_f := 0;
        ELSIF x =- 28175 THEN
            exp_f := 0;
        ELSIF x =- 28174 THEN
            exp_f := 0;
        ELSIF x =- 28173 THEN
            exp_f := 0;
        ELSIF x =- 28172 THEN
            exp_f := 0;
        ELSIF x =- 28171 THEN
            exp_f := 0;
        ELSIF x =- 28170 THEN
            exp_f := 0;
        ELSIF x =- 28169 THEN
            exp_f := 0;
        ELSIF x =- 28168 THEN
            exp_f := 0;
        ELSIF x =- 28167 THEN
            exp_f := 0;
        ELSIF x =- 28166 THEN
            exp_f := 0;
        ELSIF x =- 28165 THEN
            exp_f := 0;
        ELSIF x =- 28164 THEN
            exp_f := 0;
        ELSIF x =- 28163 THEN
            exp_f := 0;
        ELSIF x =- 28162 THEN
            exp_f := 0;
        ELSIF x =- 28161 THEN
            exp_f := 0;
        ELSIF x =- 28160 THEN
            exp_f := 0;
        ELSIF x =- 28159 THEN
            exp_f := 0;
        ELSIF x =- 28158 THEN
            exp_f := 0;
        ELSIF x =- 28157 THEN
            exp_f := 0;
        ELSIF x =- 28156 THEN
            exp_f := 0;
        ELSIF x =- 28155 THEN
            exp_f := 0;
        ELSIF x =- 28154 THEN
            exp_f := 0;
        ELSIF x =- 28153 THEN
            exp_f := 0;
        ELSIF x =- 28152 THEN
            exp_f := 0;
        ELSIF x =- 28151 THEN
            exp_f := 0;
        ELSIF x =- 28150 THEN
            exp_f := 0;
        ELSIF x =- 28149 THEN
            exp_f := 0;
        ELSIF x =- 28148 THEN
            exp_f := 0;
        ELSIF x =- 28147 THEN
            exp_f := 0;
        ELSIF x =- 28146 THEN
            exp_f := 0;
        ELSIF x =- 28145 THEN
            exp_f := 0;
        ELSIF x =- 28144 THEN
            exp_f := 0;
        ELSIF x =- 28143 THEN
            exp_f := 0;
        ELSIF x =- 28142 THEN
            exp_f := 0;
        ELSIF x =- 28141 THEN
            exp_f := 0;
        ELSIF x =- 28140 THEN
            exp_f := 0;
        ELSIF x =- 28139 THEN
            exp_f := 0;
        ELSIF x =- 28138 THEN
            exp_f := 0;
        ELSIF x =- 28137 THEN
            exp_f := 0;
        ELSIF x =- 28136 THEN
            exp_f := 0;
        ELSIF x =- 28135 THEN
            exp_f := 0;
        ELSIF x =- 28134 THEN
            exp_f := 0;
        ELSIF x =- 28133 THEN
            exp_f := 0;
        ELSIF x =- 28132 THEN
            exp_f := 0;
        ELSIF x =- 28131 THEN
            exp_f := 0;
        ELSIF x =- 28130 THEN
            exp_f := 0;
        ELSIF x =- 28129 THEN
            exp_f := 0;
        ELSIF x =- 28128 THEN
            exp_f := 0;
        ELSIF x =- 28127 THEN
            exp_f := 0;
        ELSIF x =- 28126 THEN
            exp_f := 0;
        ELSIF x =- 28125 THEN
            exp_f := 0;
        ELSIF x =- 28124 THEN
            exp_f := 0;
        ELSIF x =- 28123 THEN
            exp_f := 0;
        ELSIF x =- 28122 THEN
            exp_f := 0;
        ELSIF x =- 28121 THEN
            exp_f := 0;
        ELSIF x =- 28120 THEN
            exp_f := 0;
        ELSIF x =- 28119 THEN
            exp_f := 0;
        ELSIF x =- 28118 THEN
            exp_f := 0;
        ELSIF x =- 28117 THEN
            exp_f := 0;
        ELSIF x =- 28116 THEN
            exp_f := 0;
        ELSIF x =- 28115 THEN
            exp_f := 0;
        ELSIF x =- 28114 THEN
            exp_f := 0;
        ELSIF x =- 28113 THEN
            exp_f := 0;
        ELSIF x =- 28112 THEN
            exp_f := 0;
        ELSIF x =- 28111 THEN
            exp_f := 0;
        ELSIF x =- 28110 THEN
            exp_f := 0;
        ELSIF x =- 28109 THEN
            exp_f := 0;
        ELSIF x =- 28108 THEN
            exp_f := 0;
        ELSIF x =- 28107 THEN
            exp_f := 0;
        ELSIF x =- 28106 THEN
            exp_f := 0;
        ELSIF x =- 28105 THEN
            exp_f := 0;
        ELSIF x =- 28104 THEN
            exp_f := 0;
        ELSIF x =- 28103 THEN
            exp_f := 0;
        ELSIF x =- 28102 THEN
            exp_f := 0;
        ELSIF x =- 28101 THEN
            exp_f := 0;
        ELSIF x =- 28100 THEN
            exp_f := 0;
        ELSIF x =- 28099 THEN
            exp_f := 0;
        ELSIF x =- 28098 THEN
            exp_f := 0;
        ELSIF x =- 28097 THEN
            exp_f := 0;
        ELSIF x =- 28096 THEN
            exp_f := 0;
        ELSIF x =- 28095 THEN
            exp_f := 0;
        ELSIF x =- 28094 THEN
            exp_f := 0;
        ELSIF x =- 28093 THEN
            exp_f := 0;
        ELSIF x =- 28092 THEN
            exp_f := 0;
        ELSIF x =- 28091 THEN
            exp_f := 0;
        ELSIF x =- 28090 THEN
            exp_f := 0;
        ELSIF x =- 28089 THEN
            exp_f := 0;
        ELSIF x =- 28088 THEN
            exp_f := 0;
        ELSIF x =- 28087 THEN
            exp_f := 0;
        ELSIF x =- 28086 THEN
            exp_f := 0;
        ELSIF x =- 28085 THEN
            exp_f := 0;
        ELSIF x =- 28084 THEN
            exp_f := 0;
        ELSIF x =- 28083 THEN
            exp_f := 0;
        ELSIF x =- 28082 THEN
            exp_f := 0;
        ELSIF x =- 28081 THEN
            exp_f := 0;
        ELSIF x =- 28080 THEN
            exp_f := 0;
        ELSIF x =- 28079 THEN
            exp_f := 0;
        ELSIF x =- 28078 THEN
            exp_f := 0;
        ELSIF x =- 28077 THEN
            exp_f := 0;
        ELSIF x =- 28076 THEN
            exp_f := 0;
        ELSIF x =- 28075 THEN
            exp_f := 0;
        ELSIF x =- 28074 THEN
            exp_f := 0;
        ELSIF x =- 28073 THEN
            exp_f := 0;
        ELSIF x =- 28072 THEN
            exp_f := 0;
        ELSIF x =- 28071 THEN
            exp_f := 0;
        ELSIF x =- 28070 THEN
            exp_f := 0;
        ELSIF x =- 28069 THEN
            exp_f := 0;
        ELSIF x =- 28068 THEN
            exp_f := 0;
        ELSIF x =- 28067 THEN
            exp_f := 0;
        ELSIF x =- 28066 THEN
            exp_f := 0;
        ELSIF x =- 28065 THEN
            exp_f := 0;
        ELSIF x =- 28064 THEN
            exp_f := 0;
        ELSIF x =- 28063 THEN
            exp_f := 0;
        ELSIF x =- 28062 THEN
            exp_f := 0;
        ELSIF x =- 28061 THEN
            exp_f := 0;
        ELSIF x =- 28060 THEN
            exp_f := 0;
        ELSIF x =- 28059 THEN
            exp_f := 0;
        ELSIF x =- 28058 THEN
            exp_f := 0;
        ELSIF x =- 28057 THEN
            exp_f := 0;
        ELSIF x =- 28056 THEN
            exp_f := 0;
        ELSIF x =- 28055 THEN
            exp_f := 0;
        ELSIF x =- 28054 THEN
            exp_f := 0;
        ELSIF x =- 28053 THEN
            exp_f := 0;
        ELSIF x =- 28052 THEN
            exp_f := 0;
        ELSIF x =- 28051 THEN
            exp_f := 0;
        ELSIF x =- 28050 THEN
            exp_f := 0;
        ELSIF x =- 28049 THEN
            exp_f := 0;
        ELSIF x =- 28048 THEN
            exp_f := 0;
        ELSIF x =- 28047 THEN
            exp_f := 0;
        ELSIF x =- 28046 THEN
            exp_f := 0;
        ELSIF x =- 28045 THEN
            exp_f := 0;
        ELSIF x =- 28044 THEN
            exp_f := 0;
        ELSIF x =- 28043 THEN
            exp_f := 0;
        ELSIF x =- 28042 THEN
            exp_f := 0;
        ELSIF x =- 28041 THEN
            exp_f := 0;
        ELSIF x =- 28040 THEN
            exp_f := 0;
        ELSIF x =- 28039 THEN
            exp_f := 0;
        ELSIF x =- 28038 THEN
            exp_f := 0;
        ELSIF x =- 28037 THEN
            exp_f := 0;
        ELSIF x =- 28036 THEN
            exp_f := 0;
        ELSIF x =- 28035 THEN
            exp_f := 0;
        ELSIF x =- 28034 THEN
            exp_f := 0;
        ELSIF x =- 28033 THEN
            exp_f := 0;
        ELSIF x =- 28032 THEN
            exp_f := 0;
        ELSIF x =- 28031 THEN
            exp_f := 0;
        ELSIF x =- 28030 THEN
            exp_f := 0;
        ELSIF x =- 28029 THEN
            exp_f := 0;
        ELSIF x =- 28028 THEN
            exp_f := 0;
        ELSIF x =- 28027 THEN
            exp_f := 0;
        ELSIF x =- 28026 THEN
            exp_f := 0;
        ELSIF x =- 28025 THEN
            exp_f := 0;
        ELSIF x =- 28024 THEN
            exp_f := 0;
        ELSIF x =- 28023 THEN
            exp_f := 0;
        ELSIF x =- 28022 THEN
            exp_f := 0;
        ELSIF x =- 28021 THEN
            exp_f := 0;
        ELSIF x =- 28020 THEN
            exp_f := 0;
        ELSIF x =- 28019 THEN
            exp_f := 0;
        ELSIF x =- 28018 THEN
            exp_f := 0;
        ELSIF x =- 28017 THEN
            exp_f := 0;
        ELSIF x =- 28016 THEN
            exp_f := 0;
        ELSIF x =- 28015 THEN
            exp_f := 0;
        ELSIF x =- 28014 THEN
            exp_f := 0;
        ELSIF x =- 28013 THEN
            exp_f := 0;
        ELSIF x =- 28012 THEN
            exp_f := 0;
        ELSIF x =- 28011 THEN
            exp_f := 0;
        ELSIF x =- 28010 THEN
            exp_f := 0;
        ELSIF x =- 28009 THEN
            exp_f := 0;
        ELSIF x =- 28008 THEN
            exp_f := 0;
        ELSIF x =- 28007 THEN
            exp_f := 0;
        ELSIF x =- 28006 THEN
            exp_f := 0;
        ELSIF x =- 28005 THEN
            exp_f := 0;
        ELSIF x =- 28004 THEN
            exp_f := 0;
        ELSIF x =- 28003 THEN
            exp_f := 0;
        ELSIF x =- 28002 THEN
            exp_f := 0;
        ELSIF x =- 28001 THEN
            exp_f := 0;
        ELSIF x =- 28000 THEN
            exp_f := 0;
        ELSIF x =- 27999 THEN
            exp_f := 0;
        ELSIF x =- 27998 THEN
            exp_f := 0;
        ELSIF x =- 27997 THEN
            exp_f := 0;
        ELSIF x =- 27996 THEN
            exp_f := 0;
        ELSIF x =- 27995 THEN
            exp_f := 0;
        ELSIF x =- 27994 THEN
            exp_f := 0;
        ELSIF x =- 27993 THEN
            exp_f := 0;
        ELSIF x =- 27992 THEN
            exp_f := 0;
        ELSIF x =- 27991 THEN
            exp_f := 0;
        ELSIF x =- 27990 THEN
            exp_f := 0;
        ELSIF x =- 27989 THEN
            exp_f := 0;
        ELSIF x =- 27988 THEN
            exp_f := 0;
        ELSIF x =- 27987 THEN
            exp_f := 0;
        ELSIF x =- 27986 THEN
            exp_f := 0;
        ELSIF x =- 27985 THEN
            exp_f := 0;
        ELSIF x =- 27984 THEN
            exp_f := 0;
        ELSIF x =- 27983 THEN
            exp_f := 0;
        ELSIF x =- 27982 THEN
            exp_f := 0;
        ELSIF x =- 27981 THEN
            exp_f := 0;
        ELSIF x =- 27980 THEN
            exp_f := 0;
        ELSIF x =- 27979 THEN
            exp_f := 0;
        ELSIF x =- 27978 THEN
            exp_f := 0;
        ELSIF x =- 27977 THEN
            exp_f := 0;
        ELSIF x =- 27976 THEN
            exp_f := 0;
        ELSIF x =- 27975 THEN
            exp_f := 0;
        ELSIF x =- 27974 THEN
            exp_f := 0;
        ELSIF x =- 27973 THEN
            exp_f := 0;
        ELSIF x =- 27972 THEN
            exp_f := 0;
        ELSIF x =- 27971 THEN
            exp_f := 0;
        ELSIF x =- 27970 THEN
            exp_f := 0;
        ELSIF x =- 27969 THEN
            exp_f := 0;
        ELSIF x =- 27968 THEN
            exp_f := 0;
        ELSIF x =- 27967 THEN
            exp_f := 0;
        ELSIF x =- 27966 THEN
            exp_f := 0;
        ELSIF x =- 27965 THEN
            exp_f := 0;
        ELSIF x =- 27964 THEN
            exp_f := 0;
        ELSIF x =- 27963 THEN
            exp_f := 0;
        ELSIF x =- 27962 THEN
            exp_f := 0;
        ELSIF x =- 27961 THEN
            exp_f := 0;
        ELSIF x =- 27960 THEN
            exp_f := 0;
        ELSIF x =- 27959 THEN
            exp_f := 0;
        ELSIF x =- 27958 THEN
            exp_f := 0;
        ELSIF x =- 27957 THEN
            exp_f := 0;
        ELSIF x =- 27956 THEN
            exp_f := 0;
        ELSIF x =- 27955 THEN
            exp_f := 0;
        ELSIF x =- 27954 THEN
            exp_f := 0;
        ELSIF x =- 27953 THEN
            exp_f := 0;
        ELSIF x =- 27952 THEN
            exp_f := 0;
        ELSIF x =- 27951 THEN
            exp_f := 0;
        ELSIF x =- 27950 THEN
            exp_f := 0;
        ELSIF x =- 27949 THEN
            exp_f := 0;
        ELSIF x =- 27948 THEN
            exp_f := 0;
        ELSIF x =- 27947 THEN
            exp_f := 0;
        ELSIF x =- 27946 THEN
            exp_f := 0;
        ELSIF x =- 27945 THEN
            exp_f := 0;
        ELSIF x =- 27944 THEN
            exp_f := 0;
        ELSIF x =- 27943 THEN
            exp_f := 0;
        ELSIF x =- 27942 THEN
            exp_f := 0;
        ELSIF x =- 27941 THEN
            exp_f := 0;
        ELSIF x =- 27940 THEN
            exp_f := 0;
        ELSIF x =- 27939 THEN
            exp_f := 0;
        ELSIF x =- 27938 THEN
            exp_f := 0;
        ELSIF x =- 27937 THEN
            exp_f := 0;
        ELSIF x =- 27936 THEN
            exp_f := 0;
        ELSIF x =- 27935 THEN
            exp_f := 0;
        ELSIF x =- 27934 THEN
            exp_f := 0;
        ELSIF x =- 27933 THEN
            exp_f := 0;
        ELSIF x =- 27932 THEN
            exp_f := 0;
        ELSIF x =- 27931 THEN
            exp_f := 0;
        ELSIF x =- 27930 THEN
            exp_f := 0;
        ELSIF x =- 27929 THEN
            exp_f := 0;
        ELSIF x =- 27928 THEN
            exp_f := 0;
        ELSIF x =- 27927 THEN
            exp_f := 0;
        ELSIF x =- 27926 THEN
            exp_f := 0;
        ELSIF x =- 27925 THEN
            exp_f := 0;
        ELSIF x =- 27924 THEN
            exp_f := 0;
        ELSIF x =- 27923 THEN
            exp_f := 0;
        ELSIF x =- 27922 THEN
            exp_f := 0;
        ELSIF x =- 27921 THEN
            exp_f := 0;
        ELSIF x =- 27920 THEN
            exp_f := 0;
        ELSIF x =- 27919 THEN
            exp_f := 0;
        ELSIF x =- 27918 THEN
            exp_f := 0;
        ELSIF x =- 27917 THEN
            exp_f := 0;
        ELSIF x =- 27916 THEN
            exp_f := 0;
        ELSIF x =- 27915 THEN
            exp_f := 0;
        ELSIF x =- 27914 THEN
            exp_f := 0;
        ELSIF x =- 27913 THEN
            exp_f := 0;
        ELSIF x =- 27912 THEN
            exp_f := 0;
        ELSIF x =- 27911 THEN
            exp_f := 0;
        ELSIF x =- 27910 THEN
            exp_f := 0;
        ELSIF x =- 27909 THEN
            exp_f := 0;
        ELSIF x =- 27908 THEN
            exp_f := 0;
        ELSIF x =- 27907 THEN
            exp_f := 0;
        ELSIF x =- 27906 THEN
            exp_f := 0;
        ELSIF x =- 27905 THEN
            exp_f := 0;
        ELSIF x =- 27904 THEN
            exp_f := 0;
        ELSIF x =- 27903 THEN
            exp_f := 0;
        ELSIF x =- 27902 THEN
            exp_f := 0;
        ELSIF x =- 27901 THEN
            exp_f := 0;
        ELSIF x =- 27900 THEN
            exp_f := 0;
        ELSIF x =- 27899 THEN
            exp_f := 0;
        ELSIF x =- 27898 THEN
            exp_f := 0;
        ELSIF x =- 27897 THEN
            exp_f := 0;
        ELSIF x =- 27896 THEN
            exp_f := 0;
        ELSIF x =- 27895 THEN
            exp_f := 0;
        ELSIF x =- 27894 THEN
            exp_f := 0;
        ELSIF x =- 27893 THEN
            exp_f := 0;
        ELSIF x =- 27892 THEN
            exp_f := 0;
        ELSIF x =- 27891 THEN
            exp_f := 0;
        ELSIF x =- 27890 THEN
            exp_f := 0;
        ELSIF x =- 27889 THEN
            exp_f := 0;
        ELSIF x =- 27888 THEN
            exp_f := 0;
        ELSIF x =- 27887 THEN
            exp_f := 0;
        ELSIF x =- 27886 THEN
            exp_f := 0;
        ELSIF x =- 27885 THEN
            exp_f := 0;
        ELSIF x =- 27884 THEN
            exp_f := 0;
        ELSIF x =- 27883 THEN
            exp_f := 0;
        ELSIF x =- 27882 THEN
            exp_f := 0;
        ELSIF x =- 27881 THEN
            exp_f := 0;
        ELSIF x =- 27880 THEN
            exp_f := 0;
        ELSIF x =- 27879 THEN
            exp_f := 0;
        ELSIF x =- 27878 THEN
            exp_f := 0;
        ELSIF x =- 27877 THEN
            exp_f := 0;
        ELSIF x =- 27876 THEN
            exp_f := 0;
        ELSIF x =- 27875 THEN
            exp_f := 0;
        ELSIF x =- 27874 THEN
            exp_f := 0;
        ELSIF x =- 27873 THEN
            exp_f := 0;
        ELSIF x =- 27872 THEN
            exp_f := 0;
        ELSIF x =- 27871 THEN
            exp_f := 0;
        ELSIF x =- 27870 THEN
            exp_f := 0;
        ELSIF x =- 27869 THEN
            exp_f := 0;
        ELSIF x =- 27868 THEN
            exp_f := 0;
        ELSIF x =- 27867 THEN
            exp_f := 0;
        ELSIF x =- 27866 THEN
            exp_f := 0;
        ELSIF x =- 27865 THEN
            exp_f := 0;
        ELSIF x =- 27864 THEN
            exp_f := 0;
        ELSIF x =- 27863 THEN
            exp_f := 0;
        ELSIF x =- 27862 THEN
            exp_f := 0;
        ELSIF x =- 27861 THEN
            exp_f := 0;
        ELSIF x =- 27860 THEN
            exp_f := 0;
        ELSIF x =- 27859 THEN
            exp_f := 0;
        ELSIF x =- 27858 THEN
            exp_f := 0;
        ELSIF x =- 27857 THEN
            exp_f := 0;
        ELSIF x =- 27856 THEN
            exp_f := 0;
        ELSIF x =- 27855 THEN
            exp_f := 0;
        ELSIF x =- 27854 THEN
            exp_f := 0;
        ELSIF x =- 27853 THEN
            exp_f := 0;
        ELSIF x =- 27852 THEN
            exp_f := 0;
        ELSIF x =- 27851 THEN
            exp_f := 0;
        ELSIF x =- 27850 THEN
            exp_f := 0;
        ELSIF x =- 27849 THEN
            exp_f := 0;
        ELSIF x =- 27848 THEN
            exp_f := 0;
        ELSIF x =- 27847 THEN
            exp_f := 0;
        ELSIF x =- 27846 THEN
            exp_f := 0;
        ELSIF x =- 27845 THEN
            exp_f := 0;
        ELSIF x =- 27844 THEN
            exp_f := 0;
        ELSIF x =- 27843 THEN
            exp_f := 0;
        ELSIF x =- 27842 THEN
            exp_f := 0;
        ELSIF x =- 27841 THEN
            exp_f := 0;
        ELSIF x =- 27840 THEN
            exp_f := 0;
        ELSIF x =- 27839 THEN
            exp_f := 0;
        ELSIF x =- 27838 THEN
            exp_f := 0;
        ELSIF x =- 27837 THEN
            exp_f := 0;
        ELSIF x =- 27836 THEN
            exp_f := 0;
        ELSIF x =- 27835 THEN
            exp_f := 0;
        ELSIF x =- 27834 THEN
            exp_f := 0;
        ELSIF x =- 27833 THEN
            exp_f := 0;
        ELSIF x =- 27832 THEN
            exp_f := 0;
        ELSIF x =- 27831 THEN
            exp_f := 0;
        ELSIF x =- 27830 THEN
            exp_f := 0;
        ELSIF x =- 27829 THEN
            exp_f := 0;
        ELSIF x =- 27828 THEN
            exp_f := 0;
        ELSIF x =- 27827 THEN
            exp_f := 0;
        ELSIF x =- 27826 THEN
            exp_f := 0;
        ELSIF x =- 27825 THEN
            exp_f := 0;
        ELSIF x =- 27824 THEN
            exp_f := 0;
        ELSIF x =- 27823 THEN
            exp_f := 0;
        ELSIF x =- 27822 THEN
            exp_f := 0;
        ELSIF x =- 27821 THEN
            exp_f := 0;
        ELSIF x =- 27820 THEN
            exp_f := 0;
        ELSIF x =- 27819 THEN
            exp_f := 0;
        ELSIF x =- 27818 THEN
            exp_f := 0;
        ELSIF x =- 27817 THEN
            exp_f := 0;
        ELSIF x =- 27816 THEN
            exp_f := 0;
        ELSIF x =- 27815 THEN
            exp_f := 0;
        ELSIF x =- 27814 THEN
            exp_f := 0;
        ELSIF x =- 27813 THEN
            exp_f := 0;
        ELSIF x =- 27812 THEN
            exp_f := 0;
        ELSIF x =- 27811 THEN
            exp_f := 0;
        ELSIF x =- 27810 THEN
            exp_f := 0;
        ELSIF x =- 27809 THEN
            exp_f := 0;
        ELSIF x =- 27808 THEN
            exp_f := 0;
        ELSIF x =- 27807 THEN
            exp_f := 0;
        ELSIF x =- 27806 THEN
            exp_f := 0;
        ELSIF x =- 27805 THEN
            exp_f := 0;
        ELSIF x =- 27804 THEN
            exp_f := 0;
        ELSIF x =- 27803 THEN
            exp_f := 0;
        ELSIF x =- 27802 THEN
            exp_f := 0;
        ELSIF x =- 27801 THEN
            exp_f := 0;
        ELSIF x =- 27800 THEN
            exp_f := 0;
        ELSIF x =- 27799 THEN
            exp_f := 0;
        ELSIF x =- 27798 THEN
            exp_f := 0;
        ELSIF x =- 27797 THEN
            exp_f := 0;
        ELSIF x =- 27796 THEN
            exp_f := 0;
        ELSIF x =- 27795 THEN
            exp_f := 0;
        ELSIF x =- 27794 THEN
            exp_f := 0;
        ELSIF x =- 27793 THEN
            exp_f := 0;
        ELSIF x =- 27792 THEN
            exp_f := 0;
        ELSIF x =- 27791 THEN
            exp_f := 0;
        ELSIF x =- 27790 THEN
            exp_f := 0;
        ELSIF x =- 27789 THEN
            exp_f := 0;
        ELSIF x =- 27788 THEN
            exp_f := 0;
        ELSIF x =- 27787 THEN
            exp_f := 0;
        ELSIF x =- 27786 THEN
            exp_f := 0;
        ELSIF x =- 27785 THEN
            exp_f := 0;
        ELSIF x =- 27784 THEN
            exp_f := 0;
        ELSIF x =- 27783 THEN
            exp_f := 0;
        ELSIF x =- 27782 THEN
            exp_f := 0;
        ELSIF x =- 27781 THEN
            exp_f := 0;
        ELSIF x =- 27780 THEN
            exp_f := 0;
        ELSIF x =- 27779 THEN
            exp_f := 0;
        ELSIF x =- 27778 THEN
            exp_f := 0;
        ELSIF x =- 27777 THEN
            exp_f := 0;
        ELSIF x =- 27776 THEN
            exp_f := 0;
        ELSIF x =- 27775 THEN
            exp_f := 0;
        ELSIF x =- 27774 THEN
            exp_f := 0;
        ELSIF x =- 27773 THEN
            exp_f := 0;
        ELSIF x =- 27772 THEN
            exp_f := 0;
        ELSIF x =- 27771 THEN
            exp_f := 0;
        ELSIF x =- 27770 THEN
            exp_f := 0;
        ELSIF x =- 27769 THEN
            exp_f := 0;
        ELSIF x =- 27768 THEN
            exp_f := 0;
        ELSIF x =- 27767 THEN
            exp_f := 0;
        ELSIF x =- 27766 THEN
            exp_f := 0;
        ELSIF x =- 27765 THEN
            exp_f := 0;
        ELSIF x =- 27764 THEN
            exp_f := 0;
        ELSIF x =- 27763 THEN
            exp_f := 0;
        ELSIF x =- 27762 THEN
            exp_f := 0;
        ELSIF x =- 27761 THEN
            exp_f := 0;
        ELSIF x =- 27760 THEN
            exp_f := 0;
        ELSIF x =- 27759 THEN
            exp_f := 0;
        ELSIF x =- 27758 THEN
            exp_f := 0;
        ELSIF x =- 27757 THEN
            exp_f := 0;
        ELSIF x =- 27756 THEN
            exp_f := 0;
        ELSIF x =- 27755 THEN
            exp_f := 0;
        ELSIF x =- 27754 THEN
            exp_f := 0;
        ELSIF x =- 27753 THEN
            exp_f := 0;
        ELSIF x =- 27752 THEN
            exp_f := 0;
        ELSIF x =- 27751 THEN
            exp_f := 0;
        ELSIF x =- 27750 THEN
            exp_f := 0;
        ELSIF x =- 27749 THEN
            exp_f := 0;
        ELSIF x =- 27748 THEN
            exp_f := 0;
        ELSIF x =- 27747 THEN
            exp_f := 0;
        ELSIF x =- 27746 THEN
            exp_f := 0;
        ELSIF x =- 27745 THEN
            exp_f := 0;
        ELSIF x =- 27744 THEN
            exp_f := 0;
        ELSIF x =- 27743 THEN
            exp_f := 0;
        ELSIF x =- 27742 THEN
            exp_f := 0;
        ELSIF x =- 27741 THEN
            exp_f := 0;
        ELSIF x =- 27740 THEN
            exp_f := 0;
        ELSIF x =- 27739 THEN
            exp_f := 0;
        ELSIF x =- 27738 THEN
            exp_f := 0;
        ELSIF x =- 27737 THEN
            exp_f := 0;
        ELSIF x =- 27736 THEN
            exp_f := 0;
        ELSIF x =- 27735 THEN
            exp_f := 0;
        ELSIF x =- 27734 THEN
            exp_f := 0;
        ELSIF x =- 27733 THEN
            exp_f := 0;
        ELSIF x =- 27732 THEN
            exp_f := 0;
        ELSIF x =- 27731 THEN
            exp_f := 0;
        ELSIF x =- 27730 THEN
            exp_f := 0;
        ELSIF x =- 27729 THEN
            exp_f := 0;
        ELSIF x =- 27728 THEN
            exp_f := 0;
        ELSIF x =- 27727 THEN
            exp_f := 0;
        ELSIF x =- 27726 THEN
            exp_f := 0;
        ELSIF x =- 27725 THEN
            exp_f := 0;
        ELSIF x =- 27724 THEN
            exp_f := 0;
        ELSIF x =- 27723 THEN
            exp_f := 0;
        ELSIF x =- 27722 THEN
            exp_f := 0;
        ELSIF x =- 27721 THEN
            exp_f := 0;
        ELSIF x =- 27720 THEN
            exp_f := 0;
        ELSIF x =- 27719 THEN
            exp_f := 0;
        ELSIF x =- 27718 THEN
            exp_f := 0;
        ELSIF x =- 27717 THEN
            exp_f := 0;
        ELSIF x =- 27716 THEN
            exp_f := 0;
        ELSIF x =- 27715 THEN
            exp_f := 0;
        ELSIF x =- 27714 THEN
            exp_f := 0;
        ELSIF x =- 27713 THEN
            exp_f := 0;
        ELSIF x =- 27712 THEN
            exp_f := 0;
        ELSIF x =- 27711 THEN
            exp_f := 0;
        ELSIF x =- 27710 THEN
            exp_f := 0;
        ELSIF x =- 27709 THEN
            exp_f := 0;
        ELSIF x =- 27708 THEN
            exp_f := 0;
        ELSIF x =- 27707 THEN
            exp_f := 0;
        ELSIF x =- 27706 THEN
            exp_f := 0;
        ELSIF x =- 27705 THEN
            exp_f := 0;
        ELSIF x =- 27704 THEN
            exp_f := 0;
        ELSIF x =- 27703 THEN
            exp_f := 0;
        ELSIF x =- 27702 THEN
            exp_f := 0;
        ELSIF x =- 27701 THEN
            exp_f := 0;
        ELSIF x =- 27700 THEN
            exp_f := 0;
        ELSIF x =- 27699 THEN
            exp_f := 0;
        ELSIF x =- 27698 THEN
            exp_f := 0;
        ELSIF x =- 27697 THEN
            exp_f := 0;
        ELSIF x =- 27696 THEN
            exp_f := 0;
        ELSIF x =- 27695 THEN
            exp_f := 0;
        ELSIF x =- 27694 THEN
            exp_f := 0;
        ELSIF x =- 27693 THEN
            exp_f := 0;
        ELSIF x =- 27692 THEN
            exp_f := 0;
        ELSIF x =- 27691 THEN
            exp_f := 0;
        ELSIF x =- 27690 THEN
            exp_f := 0;
        ELSIF x =- 27689 THEN
            exp_f := 0;
        ELSIF x =- 27688 THEN
            exp_f := 0;
        ELSIF x =- 27687 THEN
            exp_f := 0;
        ELSIF x =- 27686 THEN
            exp_f := 0;
        ELSIF x =- 27685 THEN
            exp_f := 0;
        ELSIF x =- 27684 THEN
            exp_f := 0;
        ELSIF x =- 27683 THEN
            exp_f := 0;
        ELSIF x =- 27682 THEN
            exp_f := 0;
        ELSIF x =- 27681 THEN
            exp_f := 0;
        ELSIF x =- 27680 THEN
            exp_f := 0;
        ELSIF x =- 27679 THEN
            exp_f := 0;
        ELSIF x =- 27678 THEN
            exp_f := 0;
        ELSIF x =- 27677 THEN
            exp_f := 0;
        ELSIF x =- 27676 THEN
            exp_f := 0;
        ELSIF x =- 27675 THEN
            exp_f := 0;
        ELSIF x =- 27674 THEN
            exp_f := 0;
        ELSIF x =- 27673 THEN
            exp_f := 0;
        ELSIF x =- 27672 THEN
            exp_f := 0;
        ELSIF x =- 27671 THEN
            exp_f := 0;
        ELSIF x =- 27670 THEN
            exp_f := 0;
        ELSIF x =- 27669 THEN
            exp_f := 0;
        ELSIF x =- 27668 THEN
            exp_f := 0;
        ELSIF x =- 27667 THEN
            exp_f := 0;
        ELSIF x =- 27666 THEN
            exp_f := 0;
        ELSIF x =- 27665 THEN
            exp_f := 0;
        ELSIF x =- 27664 THEN
            exp_f := 0;
        ELSIF x =- 27663 THEN
            exp_f := 0;
        ELSIF x =- 27662 THEN
            exp_f := 0;
        ELSIF x =- 27661 THEN
            exp_f := 0;
        ELSIF x =- 27660 THEN
            exp_f := 0;
        ELSIF x =- 27659 THEN
            exp_f := 0;
        ELSIF x =- 27658 THEN
            exp_f := 0;
        ELSIF x =- 27657 THEN
            exp_f := 0;
        ELSIF x =- 27656 THEN
            exp_f := 0;
        ELSIF x =- 27655 THEN
            exp_f := 0;
        ELSIF x =- 27654 THEN
            exp_f := 0;
        ELSIF x =- 27653 THEN
            exp_f := 0;
        ELSIF x =- 27652 THEN
            exp_f := 0;
        ELSIF x =- 27651 THEN
            exp_f := 0;
        ELSIF x =- 27650 THEN
            exp_f := 0;
        ELSIF x =- 27649 THEN
            exp_f := 0;
        ELSIF x =- 27648 THEN
            exp_f := 0;
        ELSIF x =- 27647 THEN
            exp_f := 0;
        ELSIF x =- 27646 THEN
            exp_f := 0;
        ELSIF x =- 27645 THEN
            exp_f := 0;
        ELSIF x =- 27644 THEN
            exp_f := 0;
        ELSIF x =- 27643 THEN
            exp_f := 0;
        ELSIF x =- 27642 THEN
            exp_f := 0;
        ELSIF x =- 27641 THEN
            exp_f := 0;
        ELSIF x =- 27640 THEN
            exp_f := 0;
        ELSIF x =- 27639 THEN
            exp_f := 0;
        ELSIF x =- 27638 THEN
            exp_f := 0;
        ELSIF x =- 27637 THEN
            exp_f := 0;
        ELSIF x =- 27636 THEN
            exp_f := 0;
        ELSIF x =- 27635 THEN
            exp_f := 0;
        ELSIF x =- 27634 THEN
            exp_f := 0;
        ELSIF x =- 27633 THEN
            exp_f := 0;
        ELSIF x =- 27632 THEN
            exp_f := 0;
        ELSIF x =- 27631 THEN
            exp_f := 0;
        ELSIF x =- 27630 THEN
            exp_f := 0;
        ELSIF x =- 27629 THEN
            exp_f := 0;
        ELSIF x =- 27628 THEN
            exp_f := 0;
        ELSIF x =- 27627 THEN
            exp_f := 0;
        ELSIF x =- 27626 THEN
            exp_f := 0;
        ELSIF x =- 27625 THEN
            exp_f := 0;
        ELSIF x =- 27624 THEN
            exp_f := 0;
        ELSIF x =- 27623 THEN
            exp_f := 0;
        ELSIF x =- 27622 THEN
            exp_f := 0;
        ELSIF x =- 27621 THEN
            exp_f := 0;
        ELSIF x =- 27620 THEN
            exp_f := 0;
        ELSIF x =- 27619 THEN
            exp_f := 0;
        ELSIF x =- 27618 THEN
            exp_f := 0;
        ELSIF x =- 27617 THEN
            exp_f := 0;
        ELSIF x =- 27616 THEN
            exp_f := 0;
        ELSIF x =- 27615 THEN
            exp_f := 0;
        ELSIF x =- 27614 THEN
            exp_f := 0;
        ELSIF x =- 27613 THEN
            exp_f := 0;
        ELSIF x =- 27612 THEN
            exp_f := 0;
        ELSIF x =- 27611 THEN
            exp_f := 0;
        ELSIF x =- 27610 THEN
            exp_f := 0;
        ELSIF x =- 27609 THEN
            exp_f := 0;
        ELSIF x =- 27608 THEN
            exp_f := 0;
        ELSIF x =- 27607 THEN
            exp_f := 0;
        ELSIF x =- 27606 THEN
            exp_f := 0;
        ELSIF x =- 27605 THEN
            exp_f := 0;
        ELSIF x =- 27604 THEN
            exp_f := 0;
        ELSIF x =- 27603 THEN
            exp_f := 0;
        ELSIF x =- 27602 THEN
            exp_f := 0;
        ELSIF x =- 27601 THEN
            exp_f := 0;
        ELSIF x =- 27600 THEN
            exp_f := 0;
        ELSIF x =- 27599 THEN
            exp_f := 0;
        ELSIF x =- 27598 THEN
            exp_f := 0;
        ELSIF x =- 27597 THEN
            exp_f := 0;
        ELSIF x =- 27596 THEN
            exp_f := 0;
        ELSIF x =- 27595 THEN
            exp_f := 0;
        ELSIF x =- 27594 THEN
            exp_f := 0;
        ELSIF x =- 27593 THEN
            exp_f := 0;
        ELSIF x =- 27592 THEN
            exp_f := 0;
        ELSIF x =- 27591 THEN
            exp_f := 0;
        ELSIF x =- 27590 THEN
            exp_f := 0;
        ELSIF x =- 27589 THEN
            exp_f := 0;
        ELSIF x =- 27588 THEN
            exp_f := 0;
        ELSIF x =- 27587 THEN
            exp_f := 0;
        ELSIF x =- 27586 THEN
            exp_f := 0;
        ELSIF x =- 27585 THEN
            exp_f := 0;
        ELSIF x =- 27584 THEN
            exp_f := 0;
        ELSIF x =- 27583 THEN
            exp_f := 0;
        ELSIF x =- 27582 THEN
            exp_f := 0;
        ELSIF x =- 27581 THEN
            exp_f := 0;
        ELSIF x =- 27580 THEN
            exp_f := 0;
        ELSIF x =- 27579 THEN
            exp_f := 0;
        ELSIF x =- 27578 THEN
            exp_f := 0;
        ELSIF x =- 27577 THEN
            exp_f := 0;
        ELSIF x =- 27576 THEN
            exp_f := 0;
        ELSIF x =- 27575 THEN
            exp_f := 0;
        ELSIF x =- 27574 THEN
            exp_f := 0;
        ELSIF x =- 27573 THEN
            exp_f := 0;
        ELSIF x =- 27572 THEN
            exp_f := 0;
        ELSIF x =- 27571 THEN
            exp_f := 0;
        ELSIF x =- 27570 THEN
            exp_f := 0;
        ELSIF x =- 27569 THEN
            exp_f := 0;
        ELSIF x =- 27568 THEN
            exp_f := 0;
        ELSIF x =- 27567 THEN
            exp_f := 0;
        ELSIF x =- 27566 THEN
            exp_f := 0;
        ELSIF x =- 27565 THEN
            exp_f := 0;
        ELSIF x =- 27564 THEN
            exp_f := 0;
        ELSIF x =- 27563 THEN
            exp_f := 0;
        ELSIF x =- 27562 THEN
            exp_f := 0;
        ELSIF x =- 27561 THEN
            exp_f := 0;
        ELSIF x =- 27560 THEN
            exp_f := 0;
        ELSIF x =- 27559 THEN
            exp_f := 0;
        ELSIF x =- 27558 THEN
            exp_f := 0;
        ELSIF x =- 27557 THEN
            exp_f := 0;
        ELSIF x =- 27556 THEN
            exp_f := 0;
        ELSIF x =- 27555 THEN
            exp_f := 0;
        ELSIF x =- 27554 THEN
            exp_f := 0;
        ELSIF x =- 27553 THEN
            exp_f := 0;
        ELSIF x =- 27552 THEN
            exp_f := 0;
        ELSIF x =- 27551 THEN
            exp_f := 0;
        ELSIF x =- 27550 THEN
            exp_f := 0;
        ELSIF x =- 27549 THEN
            exp_f := 0;
        ELSIF x =- 27548 THEN
            exp_f := 0;
        ELSIF x =- 27547 THEN
            exp_f := 0;
        ELSIF x =- 27546 THEN
            exp_f := 0;
        ELSIF x =- 27545 THEN
            exp_f := 0;
        ELSIF x =- 27544 THEN
            exp_f := 0;
        ELSIF x =- 27543 THEN
            exp_f := 0;
        ELSIF x =- 27542 THEN
            exp_f := 0;
        ELSIF x =- 27541 THEN
            exp_f := 0;
        ELSIF x =- 27540 THEN
            exp_f := 0;
        ELSIF x =- 27539 THEN
            exp_f := 0;
        ELSIF x =- 27538 THEN
            exp_f := 0;
        ELSIF x =- 27537 THEN
            exp_f := 0;
        ELSIF x =- 27536 THEN
            exp_f := 0;
        ELSIF x =- 27535 THEN
            exp_f := 0;
        ELSIF x =- 27534 THEN
            exp_f := 0;
        ELSIF x =- 27533 THEN
            exp_f := 0;
        ELSIF x =- 27532 THEN
            exp_f := 0;
        ELSIF x =- 27531 THEN
            exp_f := 0;
        ELSIF x =- 27530 THEN
            exp_f := 0;
        ELSIF x =- 27529 THEN
            exp_f := 0;
        ELSIF x =- 27528 THEN
            exp_f := 0;
        ELSIF x =- 27527 THEN
            exp_f := 0;
        ELSIF x =- 27526 THEN
            exp_f := 0;
        ELSIF x =- 27525 THEN
            exp_f := 0;
        ELSIF x =- 27524 THEN
            exp_f := 0;
        ELSIF x =- 27523 THEN
            exp_f := 0;
        ELSIF x =- 27522 THEN
            exp_f := 0;
        ELSIF x =- 27521 THEN
            exp_f := 0;
        ELSIF x =- 27520 THEN
            exp_f := 0;
        ELSIF x =- 27519 THEN
            exp_f := 0;
        ELSIF x =- 27518 THEN
            exp_f := 0;
        ELSIF x =- 27517 THEN
            exp_f := 0;
        ELSIF x =- 27516 THEN
            exp_f := 0;
        ELSIF x =- 27515 THEN
            exp_f := 0;
        ELSIF x =- 27514 THEN
            exp_f := 0;
        ELSIF x =- 27513 THEN
            exp_f := 0;
        ELSIF x =- 27512 THEN
            exp_f := 0;
        ELSIF x =- 27511 THEN
            exp_f := 0;
        ELSIF x =- 27510 THEN
            exp_f := 0;
        ELSIF x =- 27509 THEN
            exp_f := 0;
        ELSIF x =- 27508 THEN
            exp_f := 0;
        ELSIF x =- 27507 THEN
            exp_f := 0;
        ELSIF x =- 27506 THEN
            exp_f := 0;
        ELSIF x =- 27505 THEN
            exp_f := 0;
        ELSIF x =- 27504 THEN
            exp_f := 0;
        ELSIF x =- 27503 THEN
            exp_f := 0;
        ELSIF x =- 27502 THEN
            exp_f := 0;
        ELSIF x =- 27501 THEN
            exp_f := 0;
        ELSIF x =- 27500 THEN
            exp_f := 0;
        ELSIF x =- 27499 THEN
            exp_f := 0;
        ELSIF x =- 27498 THEN
            exp_f := 0;
        ELSIF x =- 27497 THEN
            exp_f := 0;
        ELSIF x =- 27496 THEN
            exp_f := 0;
        ELSIF x =- 27495 THEN
            exp_f := 0;
        ELSIF x =- 27494 THEN
            exp_f := 0;
        ELSIF x =- 27493 THEN
            exp_f := 0;
        ELSIF x =- 27492 THEN
            exp_f := 0;
        ELSIF x =- 27491 THEN
            exp_f := 0;
        ELSIF x =- 27490 THEN
            exp_f := 0;
        ELSIF x =- 27489 THEN
            exp_f := 0;
        ELSIF x =- 27488 THEN
            exp_f := 0;
        ELSIF x =- 27487 THEN
            exp_f := 0;
        ELSIF x =- 27486 THEN
            exp_f := 0;
        ELSIF x =- 27485 THEN
            exp_f := 0;
        ELSIF x =- 27484 THEN
            exp_f := 0;
        ELSIF x =- 27483 THEN
            exp_f := 0;
        ELSIF x =- 27482 THEN
            exp_f := 0;
        ELSIF x =- 27481 THEN
            exp_f := 0;
        ELSIF x =- 27480 THEN
            exp_f := 0;
        ELSIF x =- 27479 THEN
            exp_f := 0;
        ELSIF x =- 27478 THEN
            exp_f := 0;
        ELSIF x =- 27477 THEN
            exp_f := 0;
        ELSIF x =- 27476 THEN
            exp_f := 0;
        ELSIF x =- 27475 THEN
            exp_f := 0;
        ELSIF x =- 27474 THEN
            exp_f := 0;
        ELSIF x =- 27473 THEN
            exp_f := 0;
        ELSIF x =- 27472 THEN
            exp_f := 0;
        ELSIF x =- 27471 THEN
            exp_f := 0;
        ELSIF x =- 27470 THEN
            exp_f := 0;
        ELSIF x =- 27469 THEN
            exp_f := 0;
        ELSIF x =- 27468 THEN
            exp_f := 0;
        ELSIF x =- 27467 THEN
            exp_f := 0;
        ELSIF x =- 27466 THEN
            exp_f := 0;
        ELSIF x =- 27465 THEN
            exp_f := 0;
        ELSIF x =- 27464 THEN
            exp_f := 0;
        ELSIF x =- 27463 THEN
            exp_f := 0;
        ELSIF x =- 27462 THEN
            exp_f := 0;
        ELSIF x =- 27461 THEN
            exp_f := 0;
        ELSIF x =- 27460 THEN
            exp_f := 0;
        ELSIF x =- 27459 THEN
            exp_f := 0;
        ELSIF x =- 27458 THEN
            exp_f := 0;
        ELSIF x =- 27457 THEN
            exp_f := 0;
        ELSIF x =- 27456 THEN
            exp_f := 0;
        ELSIF x =- 27455 THEN
            exp_f := 0;
        ELSIF x =- 27454 THEN
            exp_f := 0;
        ELSIF x =- 27453 THEN
            exp_f := 0;
        ELSIF x =- 27452 THEN
            exp_f := 0;
        ELSIF x =- 27451 THEN
            exp_f := 0;
        ELSIF x =- 27450 THEN
            exp_f := 0;
        ELSIF x =- 27449 THEN
            exp_f := 0;
        ELSIF x =- 27448 THEN
            exp_f := 0;
        ELSIF x =- 27447 THEN
            exp_f := 0;
        ELSIF x =- 27446 THEN
            exp_f := 0;
        ELSIF x =- 27445 THEN
            exp_f := 0;
        ELSIF x =- 27444 THEN
            exp_f := 0;
        ELSIF x =- 27443 THEN
            exp_f := 0;
        ELSIF x =- 27442 THEN
            exp_f := 0;
        ELSIF x =- 27441 THEN
            exp_f := 0;
        ELSIF x =- 27440 THEN
            exp_f := 0;
        ELSIF x =- 27439 THEN
            exp_f := 0;
        ELSIF x =- 27438 THEN
            exp_f := 0;
        ELSIF x =- 27437 THEN
            exp_f := 0;
        ELSIF x =- 27436 THEN
            exp_f := 0;
        ELSIF x =- 27435 THEN
            exp_f := 0;
        ELSIF x =- 27434 THEN
            exp_f := 0;
        ELSIF x =- 27433 THEN
            exp_f := 0;
        ELSIF x =- 27432 THEN
            exp_f := 0;
        ELSIF x =- 27431 THEN
            exp_f := 0;
        ELSIF x =- 27430 THEN
            exp_f := 0;
        ELSIF x =- 27429 THEN
            exp_f := 0;
        ELSIF x =- 27428 THEN
            exp_f := 0;
        ELSIF x =- 27427 THEN
            exp_f := 0;
        ELSIF x =- 27426 THEN
            exp_f := 0;
        ELSIF x =- 27425 THEN
            exp_f := 0;
        ELSIF x =- 27424 THEN
            exp_f := 0;
        ELSIF x =- 27423 THEN
            exp_f := 0;
        ELSIF x =- 27422 THEN
            exp_f := 0;
        ELSIF x =- 27421 THEN
            exp_f := 0;
        ELSIF x =- 27420 THEN
            exp_f := 0;
        ELSIF x =- 27419 THEN
            exp_f := 0;
        ELSIF x =- 27418 THEN
            exp_f := 0;
        ELSIF x =- 27417 THEN
            exp_f := 0;
        ELSIF x =- 27416 THEN
            exp_f := 0;
        ELSIF x =- 27415 THEN
            exp_f := 0;
        ELSIF x =- 27414 THEN
            exp_f := 0;
        ELSIF x =- 27413 THEN
            exp_f := 0;
        ELSIF x =- 27412 THEN
            exp_f := 0;
        ELSIF x =- 27411 THEN
            exp_f := 0;
        ELSIF x =- 27410 THEN
            exp_f := 0;
        ELSIF x =- 27409 THEN
            exp_f := 0;
        ELSIF x =- 27408 THEN
            exp_f := 0;
        ELSIF x =- 27407 THEN
            exp_f := 0;
        ELSIF x =- 27406 THEN
            exp_f := 0;
        ELSIF x =- 27405 THEN
            exp_f := 0;
        ELSIF x =- 27404 THEN
            exp_f := 0;
        ELSIF x =- 27403 THEN
            exp_f := 0;
        ELSIF x =- 27402 THEN
            exp_f := 0;
        ELSIF x =- 27401 THEN
            exp_f := 0;
        ELSIF x =- 27400 THEN
            exp_f := 0;
        ELSIF x =- 27399 THEN
            exp_f := 0;
        ELSIF x =- 27398 THEN
            exp_f := 0;
        ELSIF x =- 27397 THEN
            exp_f := 0;
        ELSIF x =- 27396 THEN
            exp_f := 0;
        ELSIF x =- 27395 THEN
            exp_f := 0;
        ELSIF x =- 27394 THEN
            exp_f := 0;
        ELSIF x =- 27393 THEN
            exp_f := 0;
        ELSIF x =- 27392 THEN
            exp_f := 0;
        ELSIF x =- 27391 THEN
            exp_f := 0;
        ELSIF x =- 27390 THEN
            exp_f := 0;
        ELSIF x =- 27389 THEN
            exp_f := 0;
        ELSIF x =- 27388 THEN
            exp_f := 0;
        ELSIF x =- 27387 THEN
            exp_f := 0;
        ELSIF x =- 27386 THEN
            exp_f := 0;
        ELSIF x =- 27385 THEN
            exp_f := 0;
        ELSIF x =- 27384 THEN
            exp_f := 0;
        ELSIF x =- 27383 THEN
            exp_f := 0;
        ELSIF x =- 27382 THEN
            exp_f := 0;
        ELSIF x =- 27381 THEN
            exp_f := 0;
        ELSIF x =- 27380 THEN
            exp_f := 0;
        ELSIF x =- 27379 THEN
            exp_f := 0;
        ELSIF x =- 27378 THEN
            exp_f := 0;
        ELSIF x =- 27377 THEN
            exp_f := 0;
        ELSIF x =- 27376 THEN
            exp_f := 0;
        ELSIF x =- 27375 THEN
            exp_f := 0;
        ELSIF x =- 27374 THEN
            exp_f := 0;
        ELSIF x =- 27373 THEN
            exp_f := 0;
        ELSIF x =- 27372 THEN
            exp_f := 0;
        ELSIF x =- 27371 THEN
            exp_f := 0;
        ELSIF x =- 27370 THEN
            exp_f := 0;
        ELSIF x =- 27369 THEN
            exp_f := 0;
        ELSIF x =- 27368 THEN
            exp_f := 0;
        ELSIF x =- 27367 THEN
            exp_f := 0;
        ELSIF x =- 27366 THEN
            exp_f := 0;
        ELSIF x =- 27365 THEN
            exp_f := 0;
        ELSIF x =- 27364 THEN
            exp_f := 0;
        ELSIF x =- 27363 THEN
            exp_f := 0;
        ELSIF x =- 27362 THEN
            exp_f := 0;
        ELSIF x =- 27361 THEN
            exp_f := 0;
        ELSIF x =- 27360 THEN
            exp_f := 0;
        ELSIF x =- 27359 THEN
            exp_f := 0;
        ELSIF x =- 27358 THEN
            exp_f := 0;
        ELSIF x =- 27357 THEN
            exp_f := 0;
        ELSIF x =- 27356 THEN
            exp_f := 0;
        ELSIF x =- 27355 THEN
            exp_f := 0;
        ELSIF x =- 27354 THEN
            exp_f := 0;
        ELSIF x =- 27353 THEN
            exp_f := 0;
        ELSIF x =- 27352 THEN
            exp_f := 0;
        ELSIF x =- 27351 THEN
            exp_f := 0;
        ELSIF x =- 27350 THEN
            exp_f := 0;
        ELSIF x =- 27349 THEN
            exp_f := 0;
        ELSIF x =- 27348 THEN
            exp_f := 0;
        ELSIF x =- 27347 THEN
            exp_f := 0;
        ELSIF x =- 27346 THEN
            exp_f := 0;
        ELSIF x =- 27345 THEN
            exp_f := 0;
        ELSIF x =- 27344 THEN
            exp_f := 0;
        ELSIF x =- 27343 THEN
            exp_f := 0;
        ELSIF x =- 27342 THEN
            exp_f := 0;
        ELSIF x =- 27341 THEN
            exp_f := 0;
        ELSIF x =- 27340 THEN
            exp_f := 0;
        ELSIF x =- 27339 THEN
            exp_f := 0;
        ELSIF x =- 27338 THEN
            exp_f := 0;
        ELSIF x =- 27337 THEN
            exp_f := 0;
        ELSIF x =- 27336 THEN
            exp_f := 0;
        ELSIF x =- 27335 THEN
            exp_f := 0;
        ELSIF x =- 27334 THEN
            exp_f := 0;
        ELSIF x =- 27333 THEN
            exp_f := 0;
        ELSIF x =- 27332 THEN
            exp_f := 0;
        ELSIF x =- 27331 THEN
            exp_f := 0;
        ELSIF x =- 27330 THEN
            exp_f := 0;
        ELSIF x =- 27329 THEN
            exp_f := 0;
        ELSIF x =- 27328 THEN
            exp_f := 0;
        ELSIF x =- 27327 THEN
            exp_f := 0;
        ELSIF x =- 27326 THEN
            exp_f := 0;
        ELSIF x =- 27325 THEN
            exp_f := 0;
        ELSIF x =- 27324 THEN
            exp_f := 0;
        ELSIF x =- 27323 THEN
            exp_f := 0;
        ELSIF x =- 27322 THEN
            exp_f := 0;
        ELSIF x =- 27321 THEN
            exp_f := 0;
        ELSIF x =- 27320 THEN
            exp_f := 0;
        ELSIF x =- 27319 THEN
            exp_f := 0;
        ELSIF x =- 27318 THEN
            exp_f := 0;
        ELSIF x =- 27317 THEN
            exp_f := 0;
        ELSIF x =- 27316 THEN
            exp_f := 0;
        ELSIF x =- 27315 THEN
            exp_f := 0;
        ELSIF x =- 27314 THEN
            exp_f := 0;
        ELSIF x =- 27313 THEN
            exp_f := 0;
        ELSIF x =- 27312 THEN
            exp_f := 0;
        ELSIF x =- 27311 THEN
            exp_f := 0;
        ELSIF x =- 27310 THEN
            exp_f := 0;
        ELSIF x =- 27309 THEN
            exp_f := 0;
        ELSIF x =- 27308 THEN
            exp_f := 0;
        ELSIF x =- 27307 THEN
            exp_f := 0;
        ELSIF x =- 27306 THEN
            exp_f := 0;
        ELSIF x =- 27305 THEN
            exp_f := 0;
        ELSIF x =- 27304 THEN
            exp_f := 0;
        ELSIF x =- 27303 THEN
            exp_f := 0;
        ELSIF x =- 27302 THEN
            exp_f := 0;
        ELSIF x =- 27301 THEN
            exp_f := 0;
        ELSIF x =- 27300 THEN
            exp_f := 0;
        ELSIF x =- 27299 THEN
            exp_f := 0;
        ELSIF x =- 27298 THEN
            exp_f := 0;
        ELSIF x =- 27297 THEN
            exp_f := 0;
        ELSIF x =- 27296 THEN
            exp_f := 0;
        ELSIF x =- 27295 THEN
            exp_f := 0;
        ELSIF x =- 27294 THEN
            exp_f := 0;
        ELSIF x =- 27293 THEN
            exp_f := 0;
        ELSIF x =- 27292 THEN
            exp_f := 0;
        ELSIF x =- 27291 THEN
            exp_f := 0;
        ELSIF x =- 27290 THEN
            exp_f := 0;
        ELSIF x =- 27289 THEN
            exp_f := 0;
        ELSIF x =- 27288 THEN
            exp_f := 0;
        ELSIF x =- 27287 THEN
            exp_f := 0;
        ELSIF x =- 27286 THEN
            exp_f := 0;
        ELSIF x =- 27285 THEN
            exp_f := 0;
        ELSIF x =- 27284 THEN
            exp_f := 0;
        ELSIF x =- 27283 THEN
            exp_f := 0;
        ELSIF x =- 27282 THEN
            exp_f := 0;
        ELSIF x =- 27281 THEN
            exp_f := 0;
        ELSIF x =- 27280 THEN
            exp_f := 0;
        ELSIF x =- 27279 THEN
            exp_f := 0;
        ELSIF x =- 27278 THEN
            exp_f := 0;
        ELSIF x =- 27277 THEN
            exp_f := 0;
        ELSIF x =- 27276 THEN
            exp_f := 0;
        ELSIF x =- 27275 THEN
            exp_f := 0;
        ELSIF x =- 27274 THEN
            exp_f := 0;
        ELSIF x =- 27273 THEN
            exp_f := 0;
        ELSIF x =- 27272 THEN
            exp_f := 0;
        ELSIF x =- 27271 THEN
            exp_f := 0;
        ELSIF x =- 27270 THEN
            exp_f := 0;
        ELSIF x =- 27269 THEN
            exp_f := 0;
        ELSIF x =- 27268 THEN
            exp_f := 0;
        ELSIF x =- 27267 THEN
            exp_f := 0;
        ELSIF x =- 27266 THEN
            exp_f := 0;
        ELSIF x =- 27265 THEN
            exp_f := 0;
        ELSIF x =- 27264 THEN
            exp_f := 0;
        ELSIF x =- 27263 THEN
            exp_f := 0;
        ELSIF x =- 27262 THEN
            exp_f := 0;
        ELSIF x =- 27261 THEN
            exp_f := 0;
        ELSIF x =- 27260 THEN
            exp_f := 0;
        ELSIF x =- 27259 THEN
            exp_f := 0;
        ELSIF x =- 27258 THEN
            exp_f := 0;
        ELSIF x =- 27257 THEN
            exp_f := 0;
        ELSIF x =- 27256 THEN
            exp_f := 0;
        ELSIF x =- 27255 THEN
            exp_f := 0;
        ELSIF x =- 27254 THEN
            exp_f := 0;
        ELSIF x =- 27253 THEN
            exp_f := 0;
        ELSIF x =- 27252 THEN
            exp_f := 0;
        ELSIF x =- 27251 THEN
            exp_f := 0;
        ELSIF x =- 27250 THEN
            exp_f := 0;
        ELSIF x =- 27249 THEN
            exp_f := 0;
        ELSIF x =- 27248 THEN
            exp_f := 0;
        ELSIF x =- 27247 THEN
            exp_f := 0;
        ELSIF x =- 27246 THEN
            exp_f := 0;
        ELSIF x =- 27245 THEN
            exp_f := 0;
        ELSIF x =- 27244 THEN
            exp_f := 0;
        ELSIF x =- 27243 THEN
            exp_f := 0;
        ELSIF x =- 27242 THEN
            exp_f := 0;
        ELSIF x =- 27241 THEN
            exp_f := 0;
        ELSIF x =- 27240 THEN
            exp_f := 0;
        ELSIF x =- 27239 THEN
            exp_f := 0;
        ELSIF x =- 27238 THEN
            exp_f := 0;
        ELSIF x =- 27237 THEN
            exp_f := 0;
        ELSIF x =- 27236 THEN
            exp_f := 0;
        ELSIF x =- 27235 THEN
            exp_f := 0;
        ELSIF x =- 27234 THEN
            exp_f := 0;
        ELSIF x =- 27233 THEN
            exp_f := 0;
        ELSIF x =- 27232 THEN
            exp_f := 0;
        ELSIF x =- 27231 THEN
            exp_f := 0;
        ELSIF x =- 27230 THEN
            exp_f := 0;
        ELSIF x =- 27229 THEN
            exp_f := 0;
        ELSIF x =- 27228 THEN
            exp_f := 0;
        ELSIF x =- 27227 THEN
            exp_f := 0;
        ELSIF x =- 27226 THEN
            exp_f := 0;
        ELSIF x =- 27225 THEN
            exp_f := 0;
        ELSIF x =- 27224 THEN
            exp_f := 0;
        ELSIF x =- 27223 THEN
            exp_f := 0;
        ELSIF x =- 27222 THEN
            exp_f := 0;
        ELSIF x =- 27221 THEN
            exp_f := 0;
        ELSIF x =- 27220 THEN
            exp_f := 0;
        ELSIF x =- 27219 THEN
            exp_f := 0;
        ELSIF x =- 27218 THEN
            exp_f := 0;
        ELSIF x =- 27217 THEN
            exp_f := 0;
        ELSIF x =- 27216 THEN
            exp_f := 0;
        ELSIF x =- 27215 THEN
            exp_f := 0;
        ELSIF x =- 27214 THEN
            exp_f := 0;
        ELSIF x =- 27213 THEN
            exp_f := 0;
        ELSIF x =- 27212 THEN
            exp_f := 0;
        ELSIF x =- 27211 THEN
            exp_f := 0;
        ELSIF x =- 27210 THEN
            exp_f := 0;
        ELSIF x =- 27209 THEN
            exp_f := 0;
        ELSIF x =- 27208 THEN
            exp_f := 0;
        ELSIF x =- 27207 THEN
            exp_f := 0;
        ELSIF x =- 27206 THEN
            exp_f := 0;
        ELSIF x =- 27205 THEN
            exp_f := 0;
        ELSIF x =- 27204 THEN
            exp_f := 0;
        ELSIF x =- 27203 THEN
            exp_f := 0;
        ELSIF x =- 27202 THEN
            exp_f := 0;
        ELSIF x =- 27201 THEN
            exp_f := 0;
        ELSIF x =- 27200 THEN
            exp_f := 0;
        ELSIF x =- 27199 THEN
            exp_f := 0;
        ELSIF x =- 27198 THEN
            exp_f := 0;
        ELSIF x =- 27197 THEN
            exp_f := 0;
        ELSIF x =- 27196 THEN
            exp_f := 0;
        ELSIF x =- 27195 THEN
            exp_f := 0;
        ELSIF x =- 27194 THEN
            exp_f := 0;
        ELSIF x =- 27193 THEN
            exp_f := 0;
        ELSIF x =- 27192 THEN
            exp_f := 0;
        ELSIF x =- 27191 THEN
            exp_f := 0;
        ELSIF x =- 27190 THEN
            exp_f := 0;
        ELSIF x =- 27189 THEN
            exp_f := 0;
        ELSIF x =- 27188 THEN
            exp_f := 0;
        ELSIF x =- 27187 THEN
            exp_f := 0;
        ELSIF x =- 27186 THEN
            exp_f := 0;
        ELSIF x =- 27185 THEN
            exp_f := 0;
        ELSIF x =- 27184 THEN
            exp_f := 0;
        ELSIF x =- 27183 THEN
            exp_f := 0;
        ELSIF x =- 27182 THEN
            exp_f := 0;
        ELSIF x =- 27181 THEN
            exp_f := 0;
        ELSIF x =- 27180 THEN
            exp_f := 0;
        ELSIF x =- 27179 THEN
            exp_f := 0;
        ELSIF x =- 27178 THEN
            exp_f := 0;
        ELSIF x =- 27177 THEN
            exp_f := 0;
        ELSIF x =- 27176 THEN
            exp_f := 0;
        ELSIF x =- 27175 THEN
            exp_f := 0;
        ELSIF x =- 27174 THEN
            exp_f := 0;
        ELSIF x =- 27173 THEN
            exp_f := 0;
        ELSIF x =- 27172 THEN
            exp_f := 0;
        ELSIF x =- 27171 THEN
            exp_f := 0;
        ELSIF x =- 27170 THEN
            exp_f := 0;
        ELSIF x =- 27169 THEN
            exp_f := 0;
        ELSIF x =- 27168 THEN
            exp_f := 0;
        ELSIF x =- 27167 THEN
            exp_f := 0;
        ELSIF x =- 27166 THEN
            exp_f := 0;
        ELSIF x =- 27165 THEN
            exp_f := 0;
        ELSIF x =- 27164 THEN
            exp_f := 0;
        ELSIF x =- 27163 THEN
            exp_f := 0;
        ELSIF x =- 27162 THEN
            exp_f := 0;
        ELSIF x =- 27161 THEN
            exp_f := 0;
        ELSIF x =- 27160 THEN
            exp_f := 0;
        ELSIF x =- 27159 THEN
            exp_f := 0;
        ELSIF x =- 27158 THEN
            exp_f := 0;
        ELSIF x =- 27157 THEN
            exp_f := 0;
        ELSIF x =- 27156 THEN
            exp_f := 0;
        ELSIF x =- 27155 THEN
            exp_f := 0;
        ELSIF x =- 27154 THEN
            exp_f := 0;
        ELSIF x =- 27153 THEN
            exp_f := 0;
        ELSIF x =- 27152 THEN
            exp_f := 0;
        ELSIF x =- 27151 THEN
            exp_f := 0;
        ELSIF x =- 27150 THEN
            exp_f := 0;
        ELSIF x =- 27149 THEN
            exp_f := 0;
        ELSIF x =- 27148 THEN
            exp_f := 0;
        ELSIF x =- 27147 THEN
            exp_f := 0;
        ELSIF x =- 27146 THEN
            exp_f := 0;
        ELSIF x =- 27145 THEN
            exp_f := 0;
        ELSIF x =- 27144 THEN
            exp_f := 0;
        ELSIF x =- 27143 THEN
            exp_f := 0;
        ELSIF x =- 27142 THEN
            exp_f := 0;
        ELSIF x =- 27141 THEN
            exp_f := 0;
        ELSIF x =- 27140 THEN
            exp_f := 0;
        ELSIF x =- 27139 THEN
            exp_f := 0;
        ELSIF x =- 27138 THEN
            exp_f := 0;
        ELSIF x =- 27137 THEN
            exp_f := 0;
        ELSIF x =- 27136 THEN
            exp_f := 0;
        ELSIF x =- 27135 THEN
            exp_f := 0;
        ELSIF x =- 27134 THEN
            exp_f := 0;
        ELSIF x =- 27133 THEN
            exp_f := 0;
        ELSIF x =- 27132 THEN
            exp_f := 0;
        ELSIF x =- 27131 THEN
            exp_f := 0;
        ELSIF x =- 27130 THEN
            exp_f := 0;
        ELSIF x =- 27129 THEN
            exp_f := 0;
        ELSIF x =- 27128 THEN
            exp_f := 0;
        ELSIF x =- 27127 THEN
            exp_f := 0;
        ELSIF x =- 27126 THEN
            exp_f := 0;
        ELSIF x =- 27125 THEN
            exp_f := 0;
        ELSIF x =- 27124 THEN
            exp_f := 0;
        ELSIF x =- 27123 THEN
            exp_f := 0;
        ELSIF x =- 27122 THEN
            exp_f := 0;
        ELSIF x =- 27121 THEN
            exp_f := 0;
        ELSIF x =- 27120 THEN
            exp_f := 0;
        ELSIF x =- 27119 THEN
            exp_f := 0;
        ELSIF x =- 27118 THEN
            exp_f := 0;
        ELSIF x =- 27117 THEN
            exp_f := 0;
        ELSIF x =- 27116 THEN
            exp_f := 0;
        ELSIF x =- 27115 THEN
            exp_f := 0;
        ELSIF x =- 27114 THEN
            exp_f := 0;
        ELSIF x =- 27113 THEN
            exp_f := 0;
        ELSIF x =- 27112 THEN
            exp_f := 0;
        ELSIF x =- 27111 THEN
            exp_f := 0;
        ELSIF x =- 27110 THEN
            exp_f := 0;
        ELSIF x =- 27109 THEN
            exp_f := 0;
        ELSIF x =- 27108 THEN
            exp_f := 0;
        ELSIF x =- 27107 THEN
            exp_f := 0;
        ELSIF x =- 27106 THEN
            exp_f := 0;
        ELSIF x =- 27105 THEN
            exp_f := 0;
        ELSIF x =- 27104 THEN
            exp_f := 0;
        ELSIF x =- 27103 THEN
            exp_f := 0;
        ELSIF x =- 27102 THEN
            exp_f := 0;
        ELSIF x =- 27101 THEN
            exp_f := 0;
        ELSIF x =- 27100 THEN
            exp_f := 0;
        ELSIF x =- 27099 THEN
            exp_f := 0;
        ELSIF x =- 27098 THEN
            exp_f := 0;
        ELSIF x =- 27097 THEN
            exp_f := 0;
        ELSIF x =- 27096 THEN
            exp_f := 0;
        ELSIF x =- 27095 THEN
            exp_f := 0;
        ELSIF x =- 27094 THEN
            exp_f := 0;
        ELSIF x =- 27093 THEN
            exp_f := 0;
        ELSIF x =- 27092 THEN
            exp_f := 0;
        ELSIF x =- 27091 THEN
            exp_f := 0;
        ELSIF x =- 27090 THEN
            exp_f := 0;
        ELSIF x =- 27089 THEN
            exp_f := 0;
        ELSIF x =- 27088 THEN
            exp_f := 0;
        ELSIF x =- 27087 THEN
            exp_f := 0;
        ELSIF x =- 27086 THEN
            exp_f := 0;
        ELSIF x =- 27085 THEN
            exp_f := 0;
        ELSIF x =- 27084 THEN
            exp_f := 0;
        ELSIF x =- 27083 THEN
            exp_f := 0;
        ELSIF x =- 27082 THEN
            exp_f := 0;
        ELSIF x =- 27081 THEN
            exp_f := 0;
        ELSIF x =- 27080 THEN
            exp_f := 0;
        ELSIF x =- 27079 THEN
            exp_f := 0;
        ELSIF x =- 27078 THEN
            exp_f := 0;
        ELSIF x =- 27077 THEN
            exp_f := 0;
        ELSIF x =- 27076 THEN
            exp_f := 0;
        ELSIF x =- 27075 THEN
            exp_f := 0;
        ELSIF x =- 27074 THEN
            exp_f := 0;
        ELSIF x =- 27073 THEN
            exp_f := 0;
        ELSIF x =- 27072 THEN
            exp_f := 0;
        ELSIF x =- 27071 THEN
            exp_f := 0;
        ELSIF x =- 27070 THEN
            exp_f := 0;
        ELSIF x =- 27069 THEN
            exp_f := 0;
        ELSIF x =- 27068 THEN
            exp_f := 0;
        ELSIF x =- 27067 THEN
            exp_f := 0;
        ELSIF x =- 27066 THEN
            exp_f := 0;
        ELSIF x =- 27065 THEN
            exp_f := 0;
        ELSIF x =- 27064 THEN
            exp_f := 0;
        ELSIF x =- 27063 THEN
            exp_f := 0;
        ELSIF x =- 27062 THEN
            exp_f := 0;
        ELSIF x =- 27061 THEN
            exp_f := 0;
        ELSIF x =- 27060 THEN
            exp_f := 0;
        ELSIF x =- 27059 THEN
            exp_f := 0;
        ELSIF x =- 27058 THEN
            exp_f := 0;
        ELSIF x =- 27057 THEN
            exp_f := 0;
        ELSIF x =- 27056 THEN
            exp_f := 0;
        ELSIF x =- 27055 THEN
            exp_f := 0;
        ELSIF x =- 27054 THEN
            exp_f := 0;
        ELSIF x =- 27053 THEN
            exp_f := 0;
        ELSIF x =- 27052 THEN
            exp_f := 0;
        ELSIF x =- 27051 THEN
            exp_f := 0;
        ELSIF x =- 27050 THEN
            exp_f := 0;
        ELSIF x =- 27049 THEN
            exp_f := 0;
        ELSIF x =- 27048 THEN
            exp_f := 0;
        ELSIF x =- 27047 THEN
            exp_f := 0;
        ELSIF x =- 27046 THEN
            exp_f := 0;
        ELSIF x =- 27045 THEN
            exp_f := 0;
        ELSIF x =- 27044 THEN
            exp_f := 0;
        ELSIF x =- 27043 THEN
            exp_f := 0;
        ELSIF x =- 27042 THEN
            exp_f := 0;
        ELSIF x =- 27041 THEN
            exp_f := 0;
        ELSIF x =- 27040 THEN
            exp_f := 0;
        ELSIF x =- 27039 THEN
            exp_f := 0;
        ELSIF x =- 27038 THEN
            exp_f := 0;
        ELSIF x =- 27037 THEN
            exp_f := 0;
        ELSIF x =- 27036 THEN
            exp_f := 0;
        ELSIF x =- 27035 THEN
            exp_f := 0;
        ELSIF x =- 27034 THEN
            exp_f := 0;
        ELSIF x =- 27033 THEN
            exp_f := 0;
        ELSIF x =- 27032 THEN
            exp_f := 0;
        ELSIF x =- 27031 THEN
            exp_f := 0;
        ELSIF x =- 27030 THEN
            exp_f := 0;
        ELSIF x =- 27029 THEN
            exp_f := 0;
        ELSIF x =- 27028 THEN
            exp_f := 0;
        ELSIF x =- 27027 THEN
            exp_f := 0;
        ELSIF x =- 27026 THEN
            exp_f := 0;
        ELSIF x =- 27025 THEN
            exp_f := 0;
        ELSIF x =- 27024 THEN
            exp_f := 0;
        ELSIF x =- 27023 THEN
            exp_f := 0;
        ELSIF x =- 27022 THEN
            exp_f := 0;
        ELSIF x =- 27021 THEN
            exp_f := 0;
        ELSIF x =- 27020 THEN
            exp_f := 0;
        ELSIF x =- 27019 THEN
            exp_f := 0;
        ELSIF x =- 27018 THEN
            exp_f := 0;
        ELSIF x =- 27017 THEN
            exp_f := 0;
        ELSIF x =- 27016 THEN
            exp_f := 0;
        ELSIF x =- 27015 THEN
            exp_f := 0;
        ELSIF x =- 27014 THEN
            exp_f := 0;
        ELSIF x =- 27013 THEN
            exp_f := 0;
        ELSIF x =- 27012 THEN
            exp_f := 0;
        ELSIF x =- 27011 THEN
            exp_f := 0;
        ELSIF x =- 27010 THEN
            exp_f := 0;
        ELSIF x =- 27009 THEN
            exp_f := 0;
        ELSIF x =- 27008 THEN
            exp_f := 0;
        ELSIF x =- 27007 THEN
            exp_f := 0;
        ELSIF x =- 27006 THEN
            exp_f := 0;
        ELSIF x =- 27005 THEN
            exp_f := 0;
        ELSIF x =- 27004 THEN
            exp_f := 0;
        ELSIF x =- 27003 THEN
            exp_f := 0;
        ELSIF x =- 27002 THEN
            exp_f := 0;
        ELSIF x =- 27001 THEN
            exp_f := 0;
        ELSIF x =- 27000 THEN
            exp_f := 0;
        ELSIF x =- 26999 THEN
            exp_f := 0;
        ELSIF x =- 26998 THEN
            exp_f := 0;
        ELSIF x =- 26997 THEN
            exp_f := 0;
        ELSIF x =- 26996 THEN
            exp_f := 0;
        ELSIF x =- 26995 THEN
            exp_f := 0;
        ELSIF x =- 26994 THEN
            exp_f := 0;
        ELSIF x =- 26993 THEN
            exp_f := 0;
        ELSIF x =- 26992 THEN
            exp_f := 0;
        ELSIF x =- 26991 THEN
            exp_f := 0;
        ELSIF x =- 26990 THEN
            exp_f := 0;
        ELSIF x =- 26989 THEN
            exp_f := 0;
        ELSIF x =- 26988 THEN
            exp_f := 0;
        ELSIF x =- 26987 THEN
            exp_f := 0;
        ELSIF x =- 26986 THEN
            exp_f := 0;
        ELSIF x =- 26985 THEN
            exp_f := 0;
        ELSIF x =- 26984 THEN
            exp_f := 0;
        ELSIF x =- 26983 THEN
            exp_f := 0;
        ELSIF x =- 26982 THEN
            exp_f := 0;
        ELSIF x =- 26981 THEN
            exp_f := 0;
        ELSIF x =- 26980 THEN
            exp_f := 0;
        ELSIF x =- 26979 THEN
            exp_f := 0;
        ELSIF x =- 26978 THEN
            exp_f := 0;
        ELSIF x =- 26977 THEN
            exp_f := 0;
        ELSIF x =- 26976 THEN
            exp_f := 0;
        ELSIF x =- 26975 THEN
            exp_f := 0;
        ELSIF x =- 26974 THEN
            exp_f := 0;
        ELSIF x =- 26973 THEN
            exp_f := 0;
        ELSIF x =- 26972 THEN
            exp_f := 0;
        ELSIF x =- 26971 THEN
            exp_f := 0;
        ELSIF x =- 26970 THEN
            exp_f := 0;
        ELSIF x =- 26969 THEN
            exp_f := 0;
        ELSIF x =- 26968 THEN
            exp_f := 0;
        ELSIF x =- 26967 THEN
            exp_f := 0;
        ELSIF x =- 26966 THEN
            exp_f := 0;
        ELSIF x =- 26965 THEN
            exp_f := 0;
        ELSIF x =- 26964 THEN
            exp_f := 0;
        ELSIF x =- 26963 THEN
            exp_f := 0;
        ELSIF x =- 26962 THEN
            exp_f := 0;
        ELSIF x =- 26961 THEN
            exp_f := 0;
        ELSIF x =- 26960 THEN
            exp_f := 0;
        ELSIF x =- 26959 THEN
            exp_f := 0;
        ELSIF x =- 26958 THEN
            exp_f := 0;
        ELSIF x =- 26957 THEN
            exp_f := 0;
        ELSIF x =- 26956 THEN
            exp_f := 0;
        ELSIF x =- 26955 THEN
            exp_f := 0;
        ELSIF x =- 26954 THEN
            exp_f := 0;
        ELSIF x =- 26953 THEN
            exp_f := 0;
        ELSIF x =- 26952 THEN
            exp_f := 0;
        ELSIF x =- 26951 THEN
            exp_f := 0;
        ELSIF x =- 26950 THEN
            exp_f := 0;
        ELSIF x =- 26949 THEN
            exp_f := 0;
        ELSIF x =- 26948 THEN
            exp_f := 0;
        ELSIF x =- 26947 THEN
            exp_f := 0;
        ELSIF x =- 26946 THEN
            exp_f := 0;
        ELSIF x =- 26945 THEN
            exp_f := 0;
        ELSIF x =- 26944 THEN
            exp_f := 0;
        ELSIF x =- 26943 THEN
            exp_f := 0;
        ELSIF x =- 26942 THEN
            exp_f := 0;
        ELSIF x =- 26941 THEN
            exp_f := 0;
        ELSIF x =- 26940 THEN
            exp_f := 0;
        ELSIF x =- 26939 THEN
            exp_f := 0;
        ELSIF x =- 26938 THEN
            exp_f := 0;
        ELSIF x =- 26937 THEN
            exp_f := 0;
        ELSIF x =- 26936 THEN
            exp_f := 0;
        ELSIF x =- 26935 THEN
            exp_f := 0;
        ELSIF x =- 26934 THEN
            exp_f := 0;
        ELSIF x =- 26933 THEN
            exp_f := 0;
        ELSIF x =- 26932 THEN
            exp_f := 0;
        ELSIF x =- 26931 THEN
            exp_f := 0;
        ELSIF x =- 26930 THEN
            exp_f := 0;
        ELSIF x =- 26929 THEN
            exp_f := 0;
        ELSIF x =- 26928 THEN
            exp_f := 0;
        ELSIF x =- 26927 THEN
            exp_f := 0;
        ELSIF x =- 26926 THEN
            exp_f := 0;
        ELSIF x =- 26925 THEN
            exp_f := 0;
        ELSIF x =- 26924 THEN
            exp_f := 0;
        ELSIF x =- 26923 THEN
            exp_f := 0;
        ELSIF x =- 26922 THEN
            exp_f := 0;
        ELSIF x =- 26921 THEN
            exp_f := 0;
        ELSIF x =- 26920 THEN
            exp_f := 0;
        ELSIF x =- 26919 THEN
            exp_f := 0;
        ELSIF x =- 26918 THEN
            exp_f := 0;
        ELSIF x =- 26917 THEN
            exp_f := 0;
        ELSIF x =- 26916 THEN
            exp_f := 0;
        ELSIF x =- 26915 THEN
            exp_f := 0;
        ELSIF x =- 26914 THEN
            exp_f := 0;
        ELSIF x =- 26913 THEN
            exp_f := 0;
        ELSIF x =- 26912 THEN
            exp_f := 0;
        ELSIF x =- 26911 THEN
            exp_f := 0;
        ELSIF x =- 26910 THEN
            exp_f := 0;
        ELSIF x =- 26909 THEN
            exp_f := 0;
        ELSIF x =- 26908 THEN
            exp_f := 0;
        ELSIF x =- 26907 THEN
            exp_f := 0;
        ELSIF x =- 26906 THEN
            exp_f := 0;
        ELSIF x =- 26905 THEN
            exp_f := 0;
        ELSIF x =- 26904 THEN
            exp_f := 0;
        ELSIF x =- 26903 THEN
            exp_f := 0;
        ELSIF x =- 26902 THEN
            exp_f := 0;
        ELSIF x =- 26901 THEN
            exp_f := 0;
        ELSIF x =- 26900 THEN
            exp_f := 0;
        ELSIF x =- 26899 THEN
            exp_f := 0;
        ELSIF x =- 26898 THEN
            exp_f := 0;
        ELSIF x =- 26897 THEN
            exp_f := 0;
        ELSIF x =- 26896 THEN
            exp_f := 0;
        ELSIF x =- 26895 THEN
            exp_f := 0;
        ELSIF x =- 26894 THEN
            exp_f := 0;
        ELSIF x =- 26893 THEN
            exp_f := 0;
        ELSIF x =- 26892 THEN
            exp_f := 0;
        ELSIF x =- 26891 THEN
            exp_f := 0;
        ELSIF x =- 26890 THEN
            exp_f := 0;
        ELSIF x =- 26889 THEN
            exp_f := 0;
        ELSIF x =- 26888 THEN
            exp_f := 0;
        ELSIF x =- 26887 THEN
            exp_f := 0;
        ELSIF x =- 26886 THEN
            exp_f := 0;
        ELSIF x =- 26885 THEN
            exp_f := 0;
        ELSIF x =- 26884 THEN
            exp_f := 0;
        ELSIF x =- 26883 THEN
            exp_f := 0;
        ELSIF x =- 26882 THEN
            exp_f := 0;
        ELSIF x =- 26881 THEN
            exp_f := 0;
        ELSIF x =- 26880 THEN
            exp_f := 0;
        ELSIF x =- 26879 THEN
            exp_f := 0;
        ELSIF x =- 26878 THEN
            exp_f := 0;
        ELSIF x =- 26877 THEN
            exp_f := 0;
        ELSIF x =- 26876 THEN
            exp_f := 0;
        ELSIF x =- 26875 THEN
            exp_f := 0;
        ELSIF x =- 26874 THEN
            exp_f := 0;
        ELSIF x =- 26873 THEN
            exp_f := 0;
        ELSIF x =- 26872 THEN
            exp_f := 0;
        ELSIF x =- 26871 THEN
            exp_f := 0;
        ELSIF x =- 26870 THEN
            exp_f := 0;
        ELSIF x =- 26869 THEN
            exp_f := 0;
        ELSIF x =- 26868 THEN
            exp_f := 0;
        ELSIF x =- 26867 THEN
            exp_f := 0;
        ELSIF x =- 26866 THEN
            exp_f := 0;
        ELSIF x =- 26865 THEN
            exp_f := 0;
        ELSIF x =- 26864 THEN
            exp_f := 0;
        ELSIF x =- 26863 THEN
            exp_f := 0;
        ELSIF x =- 26862 THEN
            exp_f := 0;
        ELSIF x =- 26861 THEN
            exp_f := 0;
        ELSIF x =- 26860 THEN
            exp_f := 0;
        ELSIF x =- 26859 THEN
            exp_f := 0;
        ELSIF x =- 26858 THEN
            exp_f := 0;
        ELSIF x =- 26857 THEN
            exp_f := 0;
        ELSIF x =- 26856 THEN
            exp_f := 0;
        ELSIF x =- 26855 THEN
            exp_f := 0;
        ELSIF x =- 26854 THEN
            exp_f := 0;
        ELSIF x =- 26853 THEN
            exp_f := 0;
        ELSIF x =- 26852 THEN
            exp_f := 0;
        ELSIF x =- 26851 THEN
            exp_f := 0;
        ELSIF x =- 26850 THEN
            exp_f := 0;
        ELSIF x =- 26849 THEN
            exp_f := 0;
        ELSIF x =- 26848 THEN
            exp_f := 0;
        ELSIF x =- 26847 THEN
            exp_f := 0;
        ELSIF x =- 26846 THEN
            exp_f := 0;
        ELSIF x =- 26845 THEN
            exp_f := 0;
        ELSIF x =- 26844 THEN
            exp_f := 0;
        ELSIF x =- 26843 THEN
            exp_f := 0;
        ELSIF x =- 26842 THEN
            exp_f := 0;
        ELSIF x =- 26841 THEN
            exp_f := 0;
        ELSIF x =- 26840 THEN
            exp_f := 0;
        ELSIF x =- 26839 THEN
            exp_f := 0;
        ELSIF x =- 26838 THEN
            exp_f := 0;
        ELSIF x =- 26837 THEN
            exp_f := 0;
        ELSIF x =- 26836 THEN
            exp_f := 0;
        ELSIF x =- 26835 THEN
            exp_f := 0;
        ELSIF x =- 26834 THEN
            exp_f := 0;
        ELSIF x =- 26833 THEN
            exp_f := 0;
        ELSIF x =- 26832 THEN
            exp_f := 0;
        ELSIF x =- 26831 THEN
            exp_f := 0;
        ELSIF x =- 26830 THEN
            exp_f := 0;
        ELSIF x =- 26829 THEN
            exp_f := 0;
        ELSIF x =- 26828 THEN
            exp_f := 0;
        ELSIF x =- 26827 THEN
            exp_f := 0;
        ELSIF x =- 26826 THEN
            exp_f := 0;
        ELSIF x =- 26825 THEN
            exp_f := 0;
        ELSIF x =- 26824 THEN
            exp_f := 0;
        ELSIF x =- 26823 THEN
            exp_f := 0;
        ELSIF x =- 26822 THEN
            exp_f := 0;
        ELSIF x =- 26821 THEN
            exp_f := 0;
        ELSIF x =- 26820 THEN
            exp_f := 0;
        ELSIF x =- 26819 THEN
            exp_f := 0;
        ELSIF x =- 26818 THEN
            exp_f := 0;
        ELSIF x =- 26817 THEN
            exp_f := 0;
        ELSIF x =- 26816 THEN
            exp_f := 0;
        ELSIF x =- 26815 THEN
            exp_f := 0;
        ELSIF x =- 26814 THEN
            exp_f := 0;
        ELSIF x =- 26813 THEN
            exp_f := 0;
        ELSIF x =- 26812 THEN
            exp_f := 0;
        ELSIF x =- 26811 THEN
            exp_f := 0;
        ELSIF x =- 26810 THEN
            exp_f := 0;
        ELSIF x =- 26809 THEN
            exp_f := 0;
        ELSIF x =- 26808 THEN
            exp_f := 0;
        ELSIF x =- 26807 THEN
            exp_f := 0;
        ELSIF x =- 26806 THEN
            exp_f := 0;
        ELSIF x =- 26805 THEN
            exp_f := 0;
        ELSIF x =- 26804 THEN
            exp_f := 0;
        ELSIF x =- 26803 THEN
            exp_f := 0;
        ELSIF x =- 26802 THEN
            exp_f := 0;
        ELSIF x =- 26801 THEN
            exp_f := 0;
        ELSIF x =- 26800 THEN
            exp_f := 0;
        ELSIF x =- 26799 THEN
            exp_f := 0;
        ELSIF x =- 26798 THEN
            exp_f := 0;
        ELSIF x =- 26797 THEN
            exp_f := 0;
        ELSIF x =- 26796 THEN
            exp_f := 0;
        ELSIF x =- 26795 THEN
            exp_f := 0;
        ELSIF x =- 26794 THEN
            exp_f := 0;
        ELSIF x =- 26793 THEN
            exp_f := 0;
        ELSIF x =- 26792 THEN
            exp_f := 0;
        ELSIF x =- 26791 THEN
            exp_f := 0;
        ELSIF x =- 26790 THEN
            exp_f := 0;
        ELSIF x =- 26789 THEN
            exp_f := 0;
        ELSIF x =- 26788 THEN
            exp_f := 0;
        ELSIF x =- 26787 THEN
            exp_f := 0;
        ELSIF x =- 26786 THEN
            exp_f := 0;
        ELSIF x =- 26785 THEN
            exp_f := 0;
        ELSIF x =- 26784 THEN
            exp_f := 0;
        ELSIF x =- 26783 THEN
            exp_f := 0;
        ELSIF x =- 26782 THEN
            exp_f := 0;
        ELSIF x =- 26781 THEN
            exp_f := 0;
        ELSIF x =- 26780 THEN
            exp_f := 0;
        ELSIF x =- 26779 THEN
            exp_f := 0;
        ELSIF x =- 26778 THEN
            exp_f := 0;
        ELSIF x =- 26777 THEN
            exp_f := 0;
        ELSIF x =- 26776 THEN
            exp_f := 0;
        ELSIF x =- 26775 THEN
            exp_f := 0;
        ELSIF x =- 26774 THEN
            exp_f := 0;
        ELSIF x =- 26773 THEN
            exp_f := 0;
        ELSIF x =- 26772 THEN
            exp_f := 0;
        ELSIF x =- 26771 THEN
            exp_f := 0;
        ELSIF x =- 26770 THEN
            exp_f := 0;
        ELSIF x =- 26769 THEN
            exp_f := 0;
        ELSIF x =- 26768 THEN
            exp_f := 0;
        ELSIF x =- 26767 THEN
            exp_f := 0;
        ELSIF x =- 26766 THEN
            exp_f := 0;
        ELSIF x =- 26765 THEN
            exp_f := 0;
        ELSIF x =- 26764 THEN
            exp_f := 0;
        ELSIF x =- 26763 THEN
            exp_f := 0;
        ELSIF x =- 26762 THEN
            exp_f := 0;
        ELSIF x =- 26761 THEN
            exp_f := 0;
        ELSIF x =- 26760 THEN
            exp_f := 0;
        ELSIF x =- 26759 THEN
            exp_f := 0;
        ELSIF x =- 26758 THEN
            exp_f := 0;
        ELSIF x =- 26757 THEN
            exp_f := 0;
        ELSIF x =- 26756 THEN
            exp_f := 0;
        ELSIF x =- 26755 THEN
            exp_f := 0;
        ELSIF x =- 26754 THEN
            exp_f := 0;
        ELSIF x =- 26753 THEN
            exp_f := 0;
        ELSIF x =- 26752 THEN
            exp_f := 0;
        ELSIF x =- 26751 THEN
            exp_f := 0;
        ELSIF x =- 26750 THEN
            exp_f := 0;
        ELSIF x =- 26749 THEN
            exp_f := 0;
        ELSIF x =- 26748 THEN
            exp_f := 0;
        ELSIF x =- 26747 THEN
            exp_f := 0;
        ELSIF x =- 26746 THEN
            exp_f := 0;
        ELSIF x =- 26745 THEN
            exp_f := 0;
        ELSIF x =- 26744 THEN
            exp_f := 0;
        ELSIF x =- 26743 THEN
            exp_f := 0;
        ELSIF x =- 26742 THEN
            exp_f := 0;
        ELSIF x =- 26741 THEN
            exp_f := 0;
        ELSIF x =- 26740 THEN
            exp_f := 0;
        ELSIF x =- 26739 THEN
            exp_f := 0;
        ELSIF x =- 26738 THEN
            exp_f := 0;
        ELSIF x =- 26737 THEN
            exp_f := 0;
        ELSIF x =- 26736 THEN
            exp_f := 0;
        ELSIF x =- 26735 THEN
            exp_f := 0;
        ELSIF x =- 26734 THEN
            exp_f := 0;
        ELSIF x =- 26733 THEN
            exp_f := 0;
        ELSIF x =- 26732 THEN
            exp_f := 0;
        ELSIF x =- 26731 THEN
            exp_f := 0;
        ELSIF x =- 26730 THEN
            exp_f := 0;
        ELSIF x =- 26729 THEN
            exp_f := 0;
        ELSIF x =- 26728 THEN
            exp_f := 0;
        ELSIF x =- 26727 THEN
            exp_f := 0;
        ELSIF x =- 26726 THEN
            exp_f := 0;
        ELSIF x =- 26725 THEN
            exp_f := 0;
        ELSIF x =- 26724 THEN
            exp_f := 0;
        ELSIF x =- 26723 THEN
            exp_f := 0;
        ELSIF x =- 26722 THEN
            exp_f := 0;
        ELSIF x =- 26721 THEN
            exp_f := 0;
        ELSIF x =- 26720 THEN
            exp_f := 0;
        ELSIF x =- 26719 THEN
            exp_f := 0;
        ELSIF x =- 26718 THEN
            exp_f := 0;
        ELSIF x =- 26717 THEN
            exp_f := 0;
        ELSIF x =- 26716 THEN
            exp_f := 0;
        ELSIF x =- 26715 THEN
            exp_f := 0;
        ELSIF x =- 26714 THEN
            exp_f := 0;
        ELSIF x =- 26713 THEN
            exp_f := 0;
        ELSIF x =- 26712 THEN
            exp_f := 0;
        ELSIF x =- 26711 THEN
            exp_f := 0;
        ELSIF x =- 26710 THEN
            exp_f := 0;
        ELSIF x =- 26709 THEN
            exp_f := 0;
        ELSIF x =- 26708 THEN
            exp_f := 0;
        ELSIF x =- 26707 THEN
            exp_f := 0;
        ELSIF x =- 26706 THEN
            exp_f := 0;
        ELSIF x =- 26705 THEN
            exp_f := 0;
        ELSIF x =- 26704 THEN
            exp_f := 0;
        ELSIF x =- 26703 THEN
            exp_f := 0;
        ELSIF x =- 26702 THEN
            exp_f := 0;
        ELSIF x =- 26701 THEN
            exp_f := 0;
        ELSIF x =- 26700 THEN
            exp_f := 0;
        ELSIF x =- 26699 THEN
            exp_f := 0;
        ELSIF x =- 26698 THEN
            exp_f := 0;
        ELSIF x =- 26697 THEN
            exp_f := 0;
        ELSIF x =- 26696 THEN
            exp_f := 0;
        ELSIF x =- 26695 THEN
            exp_f := 0;
        ELSIF x =- 26694 THEN
            exp_f := 0;
        ELSIF x =- 26693 THEN
            exp_f := 0;
        ELSIF x =- 26692 THEN
            exp_f := 0;
        ELSIF x =- 26691 THEN
            exp_f := 0;
        ELSIF x =- 26690 THEN
            exp_f := 0;
        ELSIF x =- 26689 THEN
            exp_f := 0;
        ELSIF x =- 26688 THEN
            exp_f := 0;
        ELSIF x =- 26687 THEN
            exp_f := 0;
        ELSIF x =- 26686 THEN
            exp_f := 0;
        ELSIF x =- 26685 THEN
            exp_f := 0;
        ELSIF x =- 26684 THEN
            exp_f := 0;
        ELSIF x =- 26683 THEN
            exp_f := 0;
        ELSIF x =- 26682 THEN
            exp_f := 0;
        ELSIF x =- 26681 THEN
            exp_f := 0;
        ELSIF x =- 26680 THEN
            exp_f := 0;
        ELSIF x =- 26679 THEN
            exp_f := 0;
        ELSIF x =- 26678 THEN
            exp_f := 0;
        ELSIF x =- 26677 THEN
            exp_f := 0;
        ELSIF x =- 26676 THEN
            exp_f := 0;
        ELSIF x =- 26675 THEN
            exp_f := 0;
        ELSIF x =- 26674 THEN
            exp_f := 0;
        ELSIF x =- 26673 THEN
            exp_f := 0;
        ELSIF x =- 26672 THEN
            exp_f := 0;
        ELSIF x =- 26671 THEN
            exp_f := 0;
        ELSIF x =- 26670 THEN
            exp_f := 0;
        ELSIF x =- 26669 THEN
            exp_f := 0;
        ELSIF x =- 26668 THEN
            exp_f := 0;
        ELSIF x =- 26667 THEN
            exp_f := 0;
        ELSIF x =- 26666 THEN
            exp_f := 0;
        ELSIF x =- 26665 THEN
            exp_f := 0;
        ELSIF x =- 26664 THEN
            exp_f := 0;
        ELSIF x =- 26663 THEN
            exp_f := 0;
        ELSIF x =- 26662 THEN
            exp_f := 0;
        ELSIF x =- 26661 THEN
            exp_f := 0;
        ELSIF x =- 26660 THEN
            exp_f := 0;
        ELSIF x =- 26659 THEN
            exp_f := 0;
        ELSIF x =- 26658 THEN
            exp_f := 0;
        ELSIF x =- 26657 THEN
            exp_f := 0;
        ELSIF x =- 26656 THEN
            exp_f := 0;
        ELSIF x =- 26655 THEN
            exp_f := 0;
        ELSIF x =- 26654 THEN
            exp_f := 0;
        ELSIF x =- 26653 THEN
            exp_f := 0;
        ELSIF x =- 26652 THEN
            exp_f := 0;
        ELSIF x =- 26651 THEN
            exp_f := 0;
        ELSIF x =- 26650 THEN
            exp_f := 0;
        ELSIF x =- 26649 THEN
            exp_f := 0;
        ELSIF x =- 26648 THEN
            exp_f := 0;
        ELSIF x =- 26647 THEN
            exp_f := 0;
        ELSIF x =- 26646 THEN
            exp_f := 0;
        ELSIF x =- 26645 THEN
            exp_f := 0;
        ELSIF x =- 26644 THEN
            exp_f := 0;
        ELSIF x =- 26643 THEN
            exp_f := 0;
        ELSIF x =- 26642 THEN
            exp_f := 0;
        ELSIF x =- 26641 THEN
            exp_f := 0;
        ELSIF x =- 26640 THEN
            exp_f := 0;
        ELSIF x =- 26639 THEN
            exp_f := 0;
        ELSIF x =- 26638 THEN
            exp_f := 0;
        ELSIF x =- 26637 THEN
            exp_f := 0;
        ELSIF x =- 26636 THEN
            exp_f := 0;
        ELSIF x =- 26635 THEN
            exp_f := 0;
        ELSIF x =- 26634 THEN
            exp_f := 0;
        ELSIF x =- 26633 THEN
            exp_f := 0;
        ELSIF x =- 26632 THEN
            exp_f := 0;
        ELSIF x =- 26631 THEN
            exp_f := 0;
        ELSIF x =- 26630 THEN
            exp_f := 0;
        ELSIF x =- 26629 THEN
            exp_f := 0;
        ELSIF x =- 26628 THEN
            exp_f := 0;
        ELSIF x =- 26627 THEN
            exp_f := 0;
        ELSIF x =- 26626 THEN
            exp_f := 0;
        ELSIF x =- 26625 THEN
            exp_f := 0;
        ELSIF x =- 26624 THEN
            exp_f := 0;
        ELSIF x =- 26623 THEN
            exp_f := 0;
        ELSIF x =- 26622 THEN
            exp_f := 0;
        ELSIF x =- 26621 THEN
            exp_f := 0;
        ELSIF x =- 26620 THEN
            exp_f := 0;
        ELSIF x =- 26619 THEN
            exp_f := 0;
        ELSIF x =- 26618 THEN
            exp_f := 0;
        ELSIF x =- 26617 THEN
            exp_f := 0;
        ELSIF x =- 26616 THEN
            exp_f := 0;
        ELSIF x =- 26615 THEN
            exp_f := 0;
        ELSIF x =- 26614 THEN
            exp_f := 0;
        ELSIF x =- 26613 THEN
            exp_f := 0;
        ELSIF x =- 26612 THEN
            exp_f := 0;
        ELSIF x =- 26611 THEN
            exp_f := 0;
        ELSIF x =- 26610 THEN
            exp_f := 0;
        ELSIF x =- 26609 THEN
            exp_f := 0;
        ELSIF x =- 26608 THEN
            exp_f := 0;
        ELSIF x =- 26607 THEN
            exp_f := 0;
        ELSIF x =- 26606 THEN
            exp_f := 0;
        ELSIF x =- 26605 THEN
            exp_f := 0;
        ELSIF x =- 26604 THEN
            exp_f := 0;
        ELSIF x =- 26603 THEN
            exp_f := 0;
        ELSIF x =- 26602 THEN
            exp_f := 0;
        ELSIF x =- 26601 THEN
            exp_f := 0;
        ELSIF x =- 26600 THEN
            exp_f := 0;
        ELSIF x =- 26599 THEN
            exp_f := 0;
        ELSIF x =- 26598 THEN
            exp_f := 0;
        ELSIF x =- 26597 THEN
            exp_f := 0;
        ELSIF x =- 26596 THEN
            exp_f := 0;
        ELSIF x =- 26595 THEN
            exp_f := 0;
        ELSIF x =- 26594 THEN
            exp_f := 0;
        ELSIF x =- 26593 THEN
            exp_f := 0;
        ELSIF x =- 26592 THEN
            exp_f := 0;
        ELSIF x =- 26591 THEN
            exp_f := 0;
        ELSIF x =- 26590 THEN
            exp_f := 0;
        ELSIF x =- 26589 THEN
            exp_f := 0;
        ELSIF x =- 26588 THEN
            exp_f := 0;
        ELSIF x =- 26587 THEN
            exp_f := 0;
        ELSIF x =- 26586 THEN
            exp_f := 0;
        ELSIF x =- 26585 THEN
            exp_f := 0;
        ELSIF x =- 26584 THEN
            exp_f := 0;
        ELSIF x =- 26583 THEN
            exp_f := 0;
        ELSIF x =- 26582 THEN
            exp_f := 0;
        ELSIF x =- 26581 THEN
            exp_f := 0;
        ELSIF x =- 26580 THEN
            exp_f := 0;
        ELSIF x =- 26579 THEN
            exp_f := 0;
        ELSIF x =- 26578 THEN
            exp_f := 0;
        ELSIF x =- 26577 THEN
            exp_f := 0;
        ELSIF x =- 26576 THEN
            exp_f := 0;
        ELSIF x =- 26575 THEN
            exp_f := 0;
        ELSIF x =- 26574 THEN
            exp_f := 0;
        ELSIF x =- 26573 THEN
            exp_f := 0;
        ELSIF x =- 26572 THEN
            exp_f := 0;
        ELSIF x =- 26571 THEN
            exp_f := 0;
        ELSIF x =- 26570 THEN
            exp_f := 0;
        ELSIF x =- 26569 THEN
            exp_f := 0;
        ELSIF x =- 26568 THEN
            exp_f := 0;
        ELSIF x =- 26567 THEN
            exp_f := 0;
        ELSIF x =- 26566 THEN
            exp_f := 0;
        ELSIF x =- 26565 THEN
            exp_f := 0;
        ELSIF x =- 26564 THEN
            exp_f := 0;
        ELSIF x =- 26563 THEN
            exp_f := 0;
        ELSIF x =- 26562 THEN
            exp_f := 0;
        ELSIF x =- 26561 THEN
            exp_f := 0;
        ELSIF x =- 26560 THEN
            exp_f := 0;
        ELSIF x =- 26559 THEN
            exp_f := 0;
        ELSIF x =- 26558 THEN
            exp_f := 0;
        ELSIF x =- 26557 THEN
            exp_f := 0;
        ELSIF x =- 26556 THEN
            exp_f := 0;
        ELSIF x =- 26555 THEN
            exp_f := 0;
        ELSIF x =- 26554 THEN
            exp_f := 0;
        ELSIF x =- 26553 THEN
            exp_f := 0;
        ELSIF x =- 26552 THEN
            exp_f := 0;
        ELSIF x =- 26551 THEN
            exp_f := 0;
        ELSIF x =- 26550 THEN
            exp_f := 0;
        ELSIF x =- 26549 THEN
            exp_f := 0;
        ELSIF x =- 26548 THEN
            exp_f := 0;
        ELSIF x =- 26547 THEN
            exp_f := 0;
        ELSIF x =- 26546 THEN
            exp_f := 0;
        ELSIF x =- 26545 THEN
            exp_f := 0;
        ELSIF x =- 26544 THEN
            exp_f := 0;
        ELSIF x =- 26543 THEN
            exp_f := 0;
        ELSIF x =- 26542 THEN
            exp_f := 0;
        ELSIF x =- 26541 THEN
            exp_f := 0;
        ELSIF x =- 26540 THEN
            exp_f := 0;
        ELSIF x =- 26539 THEN
            exp_f := 0;
        ELSIF x =- 26538 THEN
            exp_f := 0;
        ELSIF x =- 26537 THEN
            exp_f := 0;
        ELSIF x =- 26536 THEN
            exp_f := 0;
        ELSIF x =- 26535 THEN
            exp_f := 0;
        ELSIF x =- 26534 THEN
            exp_f := 0;
        ELSIF x =- 26533 THEN
            exp_f := 0;
        ELSIF x =- 26532 THEN
            exp_f := 0;
        ELSIF x =- 26531 THEN
            exp_f := 0;
        ELSIF x =- 26530 THEN
            exp_f := 0;
        ELSIF x =- 26529 THEN
            exp_f := 0;
        ELSIF x =- 26528 THEN
            exp_f := 0;
        ELSIF x =- 26527 THEN
            exp_f := 0;
        ELSIF x =- 26526 THEN
            exp_f := 0;
        ELSIF x =- 26525 THEN
            exp_f := 0;
        ELSIF x =- 26524 THEN
            exp_f := 0;
        ELSIF x =- 26523 THEN
            exp_f := 0;
        ELSIF x =- 26522 THEN
            exp_f := 0;
        ELSIF x =- 26521 THEN
            exp_f := 0;
        ELSIF x =- 26520 THEN
            exp_f := 0;
        ELSIF x =- 26519 THEN
            exp_f := 0;
        ELSIF x =- 26518 THEN
            exp_f := 0;
        ELSIF x =- 26517 THEN
            exp_f := 0;
        ELSIF x =- 26516 THEN
            exp_f := 0;
        ELSIF x =- 26515 THEN
            exp_f := 0;
        ELSIF x =- 26514 THEN
            exp_f := 0;
        ELSIF x =- 26513 THEN
            exp_f := 0;
        ELSIF x =- 26512 THEN
            exp_f := 0;
        ELSIF x =- 26511 THEN
            exp_f := 0;
        ELSIF x =- 26510 THEN
            exp_f := 0;
        ELSIF x =- 26509 THEN
            exp_f := 0;
        ELSIF x =- 26508 THEN
            exp_f := 0;
        ELSIF x =- 26507 THEN
            exp_f := 0;
        ELSIF x =- 26506 THEN
            exp_f := 0;
        ELSIF x =- 26505 THEN
            exp_f := 0;
        ELSIF x =- 26504 THEN
            exp_f := 0;
        ELSIF x =- 26503 THEN
            exp_f := 0;
        ELSIF x =- 26502 THEN
            exp_f := 0;
        ELSIF x =- 26501 THEN
            exp_f := 0;
        ELSIF x =- 26500 THEN
            exp_f := 0;
        ELSIF x =- 26499 THEN
            exp_f := 0;
        ELSIF x =- 26498 THEN
            exp_f := 0;
        ELSIF x =- 26497 THEN
            exp_f := 0;
        ELSIF x =- 26496 THEN
            exp_f := 0;
        ELSIF x =- 26495 THEN
            exp_f := 0;
        ELSIF x =- 26494 THEN
            exp_f := 0;
        ELSIF x =- 26493 THEN
            exp_f := 0;
        ELSIF x =- 26492 THEN
            exp_f := 0;
        ELSIF x =- 26491 THEN
            exp_f := 0;
        ELSIF x =- 26490 THEN
            exp_f := 0;
        ELSIF x =- 26489 THEN
            exp_f := 0;
        ELSIF x =- 26488 THEN
            exp_f := 0;
        ELSIF x =- 26487 THEN
            exp_f := 0;
        ELSIF x =- 26486 THEN
            exp_f := 0;
        ELSIF x =- 26485 THEN
            exp_f := 0;
        ELSIF x =- 26484 THEN
            exp_f := 0;
        ELSIF x =- 26483 THEN
            exp_f := 0;
        ELSIF x =- 26482 THEN
            exp_f := 0;
        ELSIF x =- 26481 THEN
            exp_f := 0;
        ELSIF x =- 26480 THEN
            exp_f := 0;
        ELSIF x =- 26479 THEN
            exp_f := 0;
        ELSIF x =- 26478 THEN
            exp_f := 0;
        ELSIF x =- 26477 THEN
            exp_f := 0;
        ELSIF x =- 26476 THEN
            exp_f := 0;
        ELSIF x =- 26475 THEN
            exp_f := 0;
        ELSIF x =- 26474 THEN
            exp_f := 0;
        ELSIF x =- 26473 THEN
            exp_f := 0;
        ELSIF x =- 26472 THEN
            exp_f := 0;
        ELSIF x =- 26471 THEN
            exp_f := 0;
        ELSIF x =- 26470 THEN
            exp_f := 0;
        ELSIF x =- 26469 THEN
            exp_f := 0;
        ELSIF x =- 26468 THEN
            exp_f := 0;
        ELSIF x =- 26467 THEN
            exp_f := 0;
        ELSIF x =- 26466 THEN
            exp_f := 0;
        ELSIF x =- 26465 THEN
            exp_f := 0;
        ELSIF x =- 26464 THEN
            exp_f := 0;
        ELSIF x =- 26463 THEN
            exp_f := 0;
        ELSIF x =- 26462 THEN
            exp_f := 0;
        ELSIF x =- 26461 THEN
            exp_f := 0;
        ELSIF x =- 26460 THEN
            exp_f := 0;
        ELSIF x =- 26459 THEN
            exp_f := 0;
        ELSIF x =- 26458 THEN
            exp_f := 0;
        ELSIF x =- 26457 THEN
            exp_f := 0;
        ELSIF x =- 26456 THEN
            exp_f := 0;
        ELSIF x =- 26455 THEN
            exp_f := 0;
        ELSIF x =- 26454 THEN
            exp_f := 0;
        ELSIF x =- 26453 THEN
            exp_f := 0;
        ELSIF x =- 26452 THEN
            exp_f := 0;
        ELSIF x =- 26451 THEN
            exp_f := 0;
        ELSIF x =- 26450 THEN
            exp_f := 0;
        ELSIF x =- 26449 THEN
            exp_f := 0;
        ELSIF x =- 26448 THEN
            exp_f := 0;
        ELSIF x =- 26447 THEN
            exp_f := 0;
        ELSIF x =- 26446 THEN
            exp_f := 0;
        ELSIF x =- 26445 THEN
            exp_f := 0;
        ELSIF x =- 26444 THEN
            exp_f := 0;
        ELSIF x =- 26443 THEN
            exp_f := 0;
        ELSIF x =- 26442 THEN
            exp_f := 0;
        ELSIF x =- 26441 THEN
            exp_f := 0;
        ELSIF x =- 26440 THEN
            exp_f := 0;
        ELSIF x =- 26439 THEN
            exp_f := 0;
        ELSIF x =- 26438 THEN
            exp_f := 0;
        ELSIF x =- 26437 THEN
            exp_f := 0;
        ELSIF x =- 26436 THEN
            exp_f := 0;
        ELSIF x =- 26435 THEN
            exp_f := 0;
        ELSIF x =- 26434 THEN
            exp_f := 0;
        ELSIF x =- 26433 THEN
            exp_f := 0;
        ELSIF x =- 26432 THEN
            exp_f := 0;
        ELSIF x =- 26431 THEN
            exp_f := 0;
        ELSIF x =- 26430 THEN
            exp_f := 0;
        ELSIF x =- 26429 THEN
            exp_f := 0;
        ELSIF x =- 26428 THEN
            exp_f := 0;
        ELSIF x =- 26427 THEN
            exp_f := 0;
        ELSIF x =- 26426 THEN
            exp_f := 0;
        ELSIF x =- 26425 THEN
            exp_f := 0;
        ELSIF x =- 26424 THEN
            exp_f := 0;
        ELSIF x =- 26423 THEN
            exp_f := 0;
        ELSIF x =- 26422 THEN
            exp_f := 0;
        ELSIF x =- 26421 THEN
            exp_f := 0;
        ELSIF x =- 26420 THEN
            exp_f := 0;
        ELSIF x =- 26419 THEN
            exp_f := 0;
        ELSIF x =- 26418 THEN
            exp_f := 0;
        ELSIF x =- 26417 THEN
            exp_f := 0;
        ELSIF x =- 26416 THEN
            exp_f := 0;
        ELSIF x =- 26415 THEN
            exp_f := 0;
        ELSIF x =- 26414 THEN
            exp_f := 0;
        ELSIF x =- 26413 THEN
            exp_f := 0;
        ELSIF x =- 26412 THEN
            exp_f := 0;
        ELSIF x =- 26411 THEN
            exp_f := 0;
        ELSIF x =- 26410 THEN
            exp_f := 0;
        ELSIF x =- 26409 THEN
            exp_f := 0;
        ELSIF x =- 26408 THEN
            exp_f := 0;
        ELSIF x =- 26407 THEN
            exp_f := 0;
        ELSIF x =- 26406 THEN
            exp_f := 0;
        ELSIF x =- 26405 THEN
            exp_f := 0;
        ELSIF x =- 26404 THEN
            exp_f := 0;
        ELSIF x =- 26403 THEN
            exp_f := 0;
        ELSIF x =- 26402 THEN
            exp_f := 0;
        ELSIF x =- 26401 THEN
            exp_f := 0;
        ELSIF x =- 26400 THEN
            exp_f := 0;
        ELSIF x =- 26399 THEN
            exp_f := 0;
        ELSIF x =- 26398 THEN
            exp_f := 0;
        ELSIF x =- 26397 THEN
            exp_f := 0;
        ELSIF x =- 26396 THEN
            exp_f := 0;
        ELSIF x =- 26395 THEN
            exp_f := 0;
        ELSIF x =- 26394 THEN
            exp_f := 0;
        ELSIF x =- 26393 THEN
            exp_f := 0;
        ELSIF x =- 26392 THEN
            exp_f := 0;
        ELSIF x =- 26391 THEN
            exp_f := 0;
        ELSIF x =- 26390 THEN
            exp_f := 0;
        ELSIF x =- 26389 THEN
            exp_f := 0;
        ELSIF x =- 26388 THEN
            exp_f := 0;
        ELSIF x =- 26387 THEN
            exp_f := 0;
        ELSIF x =- 26386 THEN
            exp_f := 0;
        ELSIF x =- 26385 THEN
            exp_f := 0;
        ELSIF x =- 26384 THEN
            exp_f := 0;
        ELSIF x =- 26383 THEN
            exp_f := 0;
        ELSIF x =- 26382 THEN
            exp_f := 0;
        ELSIF x =- 26381 THEN
            exp_f := 0;
        ELSIF x =- 26380 THEN
            exp_f := 0;
        ELSIF x =- 26379 THEN
            exp_f := 0;
        ELSIF x =- 26378 THEN
            exp_f := 0;
        ELSIF x =- 26377 THEN
            exp_f := 0;
        ELSIF x =- 26376 THEN
            exp_f := 0;
        ELSIF x =- 26375 THEN
            exp_f := 0;
        ELSIF x =- 26374 THEN
            exp_f := 0;
        ELSIF x =- 26373 THEN
            exp_f := 0;
        ELSIF x =- 26372 THEN
            exp_f := 0;
        ELSIF x =- 26371 THEN
            exp_f := 0;
        ELSIF x =- 26370 THEN
            exp_f := 0;
        ELSIF x =- 26369 THEN
            exp_f := 0;
        ELSIF x =- 26368 THEN
            exp_f := 0;
        ELSIF x =- 26367 THEN
            exp_f := 0;
        ELSIF x =- 26366 THEN
            exp_f := 0;
        ELSIF x =- 26365 THEN
            exp_f := 0;
        ELSIF x =- 26364 THEN
            exp_f := 0;
        ELSIF x =- 26363 THEN
            exp_f := 0;
        ELSIF x =- 26362 THEN
            exp_f := 0;
        ELSIF x =- 26361 THEN
            exp_f := 0;
        ELSIF x =- 26360 THEN
            exp_f := 0;
        ELSIF x =- 26359 THEN
            exp_f := 0;
        ELSIF x =- 26358 THEN
            exp_f := 0;
        ELSIF x =- 26357 THEN
            exp_f := 0;
        ELSIF x =- 26356 THEN
            exp_f := 0;
        ELSIF x =- 26355 THEN
            exp_f := 0;
        ELSIF x =- 26354 THEN
            exp_f := 0;
        ELSIF x =- 26353 THEN
            exp_f := 0;
        ELSIF x =- 26352 THEN
            exp_f := 0;
        ELSIF x =- 26351 THEN
            exp_f := 0;
        ELSIF x =- 26350 THEN
            exp_f := 0;
        ELSIF x =- 26349 THEN
            exp_f := 0;
        ELSIF x =- 26348 THEN
            exp_f := 0;
        ELSIF x =- 26347 THEN
            exp_f := 0;
        ELSIF x =- 26346 THEN
            exp_f := 0;
        ELSIF x =- 26345 THEN
            exp_f := 0;
        ELSIF x =- 26344 THEN
            exp_f := 0;
        ELSIF x =- 26343 THEN
            exp_f := 0;
        ELSIF x =- 26342 THEN
            exp_f := 0;
        ELSIF x =- 26341 THEN
            exp_f := 0;
        ELSIF x =- 26340 THEN
            exp_f := 0;
        ELSIF x =- 26339 THEN
            exp_f := 0;
        ELSIF x =- 26338 THEN
            exp_f := 0;
        ELSIF x =- 26337 THEN
            exp_f := 0;
        ELSIF x =- 26336 THEN
            exp_f := 0;
        ELSIF x =- 26335 THEN
            exp_f := 0;
        ELSIF x =- 26334 THEN
            exp_f := 0;
        ELSIF x =- 26333 THEN
            exp_f := 0;
        ELSIF x =- 26332 THEN
            exp_f := 0;
        ELSIF x =- 26331 THEN
            exp_f := 0;
        ELSIF x =- 26330 THEN
            exp_f := 0;
        ELSIF x =- 26329 THEN
            exp_f := 0;
        ELSIF x =- 26328 THEN
            exp_f := 0;
        ELSIF x =- 26327 THEN
            exp_f := 0;
        ELSIF x =- 26326 THEN
            exp_f := 0;
        ELSIF x =- 26325 THEN
            exp_f := 0;
        ELSIF x =- 26324 THEN
            exp_f := 0;
        ELSIF x =- 26323 THEN
            exp_f := 0;
        ELSIF x =- 26322 THEN
            exp_f := 0;
        ELSIF x =- 26321 THEN
            exp_f := 0;
        ELSIF x =- 26320 THEN
            exp_f := 0;
        ELSIF x =- 26319 THEN
            exp_f := 0;
        ELSIF x =- 26318 THEN
            exp_f := 0;
        ELSIF x =- 26317 THEN
            exp_f := 0;
        ELSIF x =- 26316 THEN
            exp_f := 0;
        ELSIF x =- 26315 THEN
            exp_f := 0;
        ELSIF x =- 26314 THEN
            exp_f := 0;
        ELSIF x =- 26313 THEN
            exp_f := 0;
        ELSIF x =- 26312 THEN
            exp_f := 0;
        ELSIF x =- 26311 THEN
            exp_f := 0;
        ELSIF x =- 26310 THEN
            exp_f := 0;
        ELSIF x =- 26309 THEN
            exp_f := 0;
        ELSIF x =- 26308 THEN
            exp_f := 0;
        ELSIF x =- 26307 THEN
            exp_f := 0;
        ELSIF x =- 26306 THEN
            exp_f := 0;
        ELSIF x =- 26305 THEN
            exp_f := 0;
        ELSIF x =- 26304 THEN
            exp_f := 0;
        ELSIF x =- 26303 THEN
            exp_f := 0;
        ELSIF x =- 26302 THEN
            exp_f := 0;
        ELSIF x =- 26301 THEN
            exp_f := 0;
        ELSIF x =- 26300 THEN
            exp_f := 0;
        ELSIF x =- 26299 THEN
            exp_f := 0;
        ELSIF x =- 26298 THEN
            exp_f := 0;
        ELSIF x =- 26297 THEN
            exp_f := 0;
        ELSIF x =- 26296 THEN
            exp_f := 0;
        ELSIF x =- 26295 THEN
            exp_f := 0;
        ELSIF x =- 26294 THEN
            exp_f := 0;
        ELSIF x =- 26293 THEN
            exp_f := 0;
        ELSIF x =- 26292 THEN
            exp_f := 0;
        ELSIF x =- 26291 THEN
            exp_f := 0;
        ELSIF x =- 26290 THEN
            exp_f := 0;
        ELSIF x =- 26289 THEN
            exp_f := 0;
        ELSIF x =- 26288 THEN
            exp_f := 0;
        ELSIF x =- 26287 THEN
            exp_f := 0;
        ELSIF x =- 26286 THEN
            exp_f := 0;
        ELSIF x =- 26285 THEN
            exp_f := 0;
        ELSIF x =- 26284 THEN
            exp_f := 0;
        ELSIF x =- 26283 THEN
            exp_f := 0;
        ELSIF x =- 26282 THEN
            exp_f := 0;
        ELSIF x =- 26281 THEN
            exp_f := 0;
        ELSIF x =- 26280 THEN
            exp_f := 0;
        ELSIF x =- 26279 THEN
            exp_f := 0;
        ELSIF x =- 26278 THEN
            exp_f := 0;
        ELSIF x =- 26277 THEN
            exp_f := 0;
        ELSIF x =- 26276 THEN
            exp_f := 0;
        ELSIF x =- 26275 THEN
            exp_f := 0;
        ELSIF x =- 26274 THEN
            exp_f := 0;
        ELSIF x =- 26273 THEN
            exp_f := 0;
        ELSIF x =- 26272 THEN
            exp_f := 0;
        ELSIF x =- 26271 THEN
            exp_f := 0;
        ELSIF x =- 26270 THEN
            exp_f := 0;
        ELSIF x =- 26269 THEN
            exp_f := 0;
        ELSIF x =- 26268 THEN
            exp_f := 0;
        ELSIF x =- 26267 THEN
            exp_f := 0;
        ELSIF x =- 26266 THEN
            exp_f := 0;
        ELSIF x =- 26265 THEN
            exp_f := 0;
        ELSIF x =- 26264 THEN
            exp_f := 0;
        ELSIF x =- 26263 THEN
            exp_f := 0;
        ELSIF x =- 26262 THEN
            exp_f := 0;
        ELSIF x =- 26261 THEN
            exp_f := 0;
        ELSIF x =- 26260 THEN
            exp_f := 0;
        ELSIF x =- 26259 THEN
            exp_f := 0;
        ELSIF x =- 26258 THEN
            exp_f := 0;
        ELSIF x =- 26257 THEN
            exp_f := 0;
        ELSIF x =- 26256 THEN
            exp_f := 0;
        ELSIF x =- 26255 THEN
            exp_f := 0;
        ELSIF x =- 26254 THEN
            exp_f := 0;
        ELSIF x =- 26253 THEN
            exp_f := 0;
        ELSIF x =- 26252 THEN
            exp_f := 0;
        ELSIF x =- 26251 THEN
            exp_f := 0;
        ELSIF x =- 26250 THEN
            exp_f := 0;
        ELSIF x =- 26249 THEN
            exp_f := 0;
        ELSIF x =- 26248 THEN
            exp_f := 0;
        ELSIF x =- 26247 THEN
            exp_f := 0;
        ELSIF x =- 26246 THEN
            exp_f := 0;
        ELSIF x =- 26245 THEN
            exp_f := 0;
        ELSIF x =- 26244 THEN
            exp_f := 0;
        ELSIF x =- 26243 THEN
            exp_f := 0;
        ELSIF x =- 26242 THEN
            exp_f := 0;
        ELSIF x =- 26241 THEN
            exp_f := 0;
        ELSIF x =- 26240 THEN
            exp_f := 0;
        ELSIF x =- 26239 THEN
            exp_f := 0;
        ELSIF x =- 26238 THEN
            exp_f := 0;
        ELSIF x =- 26237 THEN
            exp_f := 0;
        ELSIF x =- 26236 THEN
            exp_f := 0;
        ELSIF x =- 26235 THEN
            exp_f := 0;
        ELSIF x =- 26234 THEN
            exp_f := 0;
        ELSIF x =- 26233 THEN
            exp_f := 0;
        ELSIF x =- 26232 THEN
            exp_f := 0;
        ELSIF x =- 26231 THEN
            exp_f := 0;
        ELSIF x =- 26230 THEN
            exp_f := 0;
        ELSIF x =- 26229 THEN
            exp_f := 0;
        ELSIF x =- 26228 THEN
            exp_f := 0;
        ELSIF x =- 26227 THEN
            exp_f := 0;
        ELSIF x =- 26226 THEN
            exp_f := 0;
        ELSIF x =- 26225 THEN
            exp_f := 0;
        ELSIF x =- 26224 THEN
            exp_f := 0;
        ELSIF x =- 26223 THEN
            exp_f := 0;
        ELSIF x =- 26222 THEN
            exp_f := 0;
        ELSIF x =- 26221 THEN
            exp_f := 0;
        ELSIF x =- 26220 THEN
            exp_f := 0;
        ELSIF x =- 26219 THEN
            exp_f := 0;
        ELSIF x =- 26218 THEN
            exp_f := 0;
        ELSIF x =- 26217 THEN
            exp_f := 0;
        ELSIF x =- 26216 THEN
            exp_f := 0;
        ELSIF x =- 26215 THEN
            exp_f := 0;
        ELSIF x =- 26214 THEN
            exp_f := 0;
        ELSIF x =- 26213 THEN
            exp_f := 0;
        ELSIF x =- 26212 THEN
            exp_f := 0;
        ELSIF x =- 26211 THEN
            exp_f := 0;
        ELSIF x =- 26210 THEN
            exp_f := 0;
        ELSIF x =- 26209 THEN
            exp_f := 0;
        ELSIF x =- 26208 THEN
            exp_f := 0;
        ELSIF x =- 26207 THEN
            exp_f := 0;
        ELSIF x =- 26206 THEN
            exp_f := 0;
        ELSIF x =- 26205 THEN
            exp_f := 0;
        ELSIF x =- 26204 THEN
            exp_f := 0;
        ELSIF x =- 26203 THEN
            exp_f := 0;
        ELSIF x =- 26202 THEN
            exp_f := 0;
        ELSIF x =- 26201 THEN
            exp_f := 0;
        ELSIF x =- 26200 THEN
            exp_f := 0;
        ELSIF x =- 26199 THEN
            exp_f := 0;
        ELSIF x =- 26198 THEN
            exp_f := 0;
        ELSIF x =- 26197 THEN
            exp_f := 0;
        ELSIF x =- 26196 THEN
            exp_f := 0;
        ELSIF x =- 26195 THEN
            exp_f := 0;
        ELSIF x =- 26194 THEN
            exp_f := 0;
        ELSIF x =- 26193 THEN
            exp_f := 0;
        ELSIF x =- 26192 THEN
            exp_f := 0;
        ELSIF x =- 26191 THEN
            exp_f := 0;
        ELSIF x =- 26190 THEN
            exp_f := 0;
        ELSIF x =- 26189 THEN
            exp_f := 0;
        ELSIF x =- 26188 THEN
            exp_f := 0;
        ELSIF x =- 26187 THEN
            exp_f := 0;
        ELSIF x =- 26186 THEN
            exp_f := 0;
        ELSIF x =- 26185 THEN
            exp_f := 0;
        ELSIF x =- 26184 THEN
            exp_f := 0;
        ELSIF x =- 26183 THEN
            exp_f := 0;
        ELSIF x =- 26182 THEN
            exp_f := 0;
        ELSIF x =- 26181 THEN
            exp_f := 0;
        ELSIF x =- 26180 THEN
            exp_f := 0;
        ELSIF x =- 26179 THEN
            exp_f := 0;
        ELSIF x =- 26178 THEN
            exp_f := 0;
        ELSIF x =- 26177 THEN
            exp_f := 0;
        ELSIF x =- 26176 THEN
            exp_f := 0;
        ELSIF x =- 26175 THEN
            exp_f := 0;
        ELSIF x =- 26174 THEN
            exp_f := 0;
        ELSIF x =- 26173 THEN
            exp_f := 0;
        ELSIF x =- 26172 THEN
            exp_f := 0;
        ELSIF x =- 26171 THEN
            exp_f := 0;
        ELSIF x =- 26170 THEN
            exp_f := 0;
        ELSIF x =- 26169 THEN
            exp_f := 0;
        ELSIF x =- 26168 THEN
            exp_f := 0;
        ELSIF x =- 26167 THEN
            exp_f := 0;
        ELSIF x =- 26166 THEN
            exp_f := 0;
        ELSIF x =- 26165 THEN
            exp_f := 0;
        ELSIF x =- 26164 THEN
            exp_f := 0;
        ELSIF x =- 26163 THEN
            exp_f := 0;
        ELSIF x =- 26162 THEN
            exp_f := 0;
        ELSIF x =- 26161 THEN
            exp_f := 0;
        ELSIF x =- 26160 THEN
            exp_f := 0;
        ELSIF x =- 26159 THEN
            exp_f := 0;
        ELSIF x =- 26158 THEN
            exp_f := 0;
        ELSIF x =- 26157 THEN
            exp_f := 0;
        ELSIF x =- 26156 THEN
            exp_f := 0;
        ELSIF x =- 26155 THEN
            exp_f := 0;
        ELSIF x =- 26154 THEN
            exp_f := 0;
        ELSIF x =- 26153 THEN
            exp_f := 0;
        ELSIF x =- 26152 THEN
            exp_f := 0;
        ELSIF x =- 26151 THEN
            exp_f := 0;
        ELSIF x =- 26150 THEN
            exp_f := 0;
        ELSIF x =- 26149 THEN
            exp_f := 0;
        ELSIF x =- 26148 THEN
            exp_f := 0;
        ELSIF x =- 26147 THEN
            exp_f := 0;
        ELSIF x =- 26146 THEN
            exp_f := 0;
        ELSIF x =- 26145 THEN
            exp_f := 0;
        ELSIF x =- 26144 THEN
            exp_f := 0;
        ELSIF x =- 26143 THEN
            exp_f := 0;
        ELSIF x =- 26142 THEN
            exp_f := 0;
        ELSIF x =- 26141 THEN
            exp_f := 0;
        ELSIF x =- 26140 THEN
            exp_f := 0;
        ELSIF x =- 26139 THEN
            exp_f := 0;
        ELSIF x =- 26138 THEN
            exp_f := 0;
        ELSIF x =- 26137 THEN
            exp_f := 0;
        ELSIF x =- 26136 THEN
            exp_f := 0;
        ELSIF x =- 26135 THEN
            exp_f := 0;
        ELSIF x =- 26134 THEN
            exp_f := 0;
        ELSIF x =- 26133 THEN
            exp_f := 0;
        ELSIF x =- 26132 THEN
            exp_f := 0;
        ELSIF x =- 26131 THEN
            exp_f := 0;
        ELSIF x =- 26130 THEN
            exp_f := 0;
        ELSIF x =- 26129 THEN
            exp_f := 0;
        ELSIF x =- 26128 THEN
            exp_f := 0;
        ELSIF x =- 26127 THEN
            exp_f := 0;
        ELSIF x =- 26126 THEN
            exp_f := 0;
        ELSIF x =- 26125 THEN
            exp_f := 0;
        ELSIF x =- 26124 THEN
            exp_f := 0;
        ELSIF x =- 26123 THEN
            exp_f := 0;
        ELSIF x =- 26122 THEN
            exp_f := 0;
        ELSIF x =- 26121 THEN
            exp_f := 0;
        ELSIF x =- 26120 THEN
            exp_f := 0;
        ELSIF x =- 26119 THEN
            exp_f := 0;
        ELSIF x =- 26118 THEN
            exp_f := 0;
        ELSIF x =- 26117 THEN
            exp_f := 0;
        ELSIF x =- 26116 THEN
            exp_f := 0;
        ELSIF x =- 26115 THEN
            exp_f := 0;
        ELSIF x =- 26114 THEN
            exp_f := 0;
        ELSIF x =- 26113 THEN
            exp_f := 0;
        ELSIF x =- 26112 THEN
            exp_f := 0;
        ELSIF x =- 26111 THEN
            exp_f := 0;
        ELSIF x =- 26110 THEN
            exp_f := 0;
        ELSIF x =- 26109 THEN
            exp_f := 0;
        ELSIF x =- 26108 THEN
            exp_f := 0;
        ELSIF x =- 26107 THEN
            exp_f := 0;
        ELSIF x =- 26106 THEN
            exp_f := 0;
        ELSIF x =- 26105 THEN
            exp_f := 0;
        ELSIF x =- 26104 THEN
            exp_f := 0;
        ELSIF x =- 26103 THEN
            exp_f := 0;
        ELSIF x =- 26102 THEN
            exp_f := 0;
        ELSIF x =- 26101 THEN
            exp_f := 0;
        ELSIF x =- 26100 THEN
            exp_f := 0;
        ELSIF x =- 26099 THEN
            exp_f := 0;
        ELSIF x =- 26098 THEN
            exp_f := 0;
        ELSIF x =- 26097 THEN
            exp_f := 0;
        ELSIF x =- 26096 THEN
            exp_f := 0;
        ELSIF x =- 26095 THEN
            exp_f := 0;
        ELSIF x =- 26094 THEN
            exp_f := 0;
        ELSIF x =- 26093 THEN
            exp_f := 0;
        ELSIF x =- 26092 THEN
            exp_f := 0;
        ELSIF x =- 26091 THEN
            exp_f := 0;
        ELSIF x =- 26090 THEN
            exp_f := 0;
        ELSIF x =- 26089 THEN
            exp_f := 0;
        ELSIF x =- 26088 THEN
            exp_f := 0;
        ELSIF x =- 26087 THEN
            exp_f := 0;
        ELSIF x =- 26086 THEN
            exp_f := 0;
        ELSIF x =- 26085 THEN
            exp_f := 0;
        ELSIF x =- 26084 THEN
            exp_f := 0;
        ELSIF x =- 26083 THEN
            exp_f := 0;
        ELSIF x =- 26082 THEN
            exp_f := 0;
        ELSIF x =- 26081 THEN
            exp_f := 0;
        ELSIF x =- 26080 THEN
            exp_f := 0;
        ELSIF x =- 26079 THEN
            exp_f := 0;
        ELSIF x =- 26078 THEN
            exp_f := 0;
        ELSIF x =- 26077 THEN
            exp_f := 0;
        ELSIF x =- 26076 THEN
            exp_f := 0;
        ELSIF x =- 26075 THEN
            exp_f := 0;
        ELSIF x =- 26074 THEN
            exp_f := 0;
        ELSIF x =- 26073 THEN
            exp_f := 0;
        ELSIF x =- 26072 THEN
            exp_f := 0;
        ELSIF x =- 26071 THEN
            exp_f := 0;
        ELSIF x =- 26070 THEN
            exp_f := 0;
        ELSIF x =- 26069 THEN
            exp_f := 0;
        ELSIF x =- 26068 THEN
            exp_f := 0;
        ELSIF x =- 26067 THEN
            exp_f := 0;
        ELSIF x =- 26066 THEN
            exp_f := 0;
        ELSIF x =- 26065 THEN
            exp_f := 0;
        ELSIF x =- 26064 THEN
            exp_f := 0;
        ELSIF x =- 26063 THEN
            exp_f := 0;
        ELSIF x =- 26062 THEN
            exp_f := 0;
        ELSIF x =- 26061 THEN
            exp_f := 0;
        ELSIF x =- 26060 THEN
            exp_f := 0;
        ELSIF x =- 26059 THEN
            exp_f := 0;
        ELSIF x =- 26058 THEN
            exp_f := 0;
        ELSIF x =- 26057 THEN
            exp_f := 0;
        ELSIF x =- 26056 THEN
            exp_f := 0;
        ELSIF x =- 26055 THEN
            exp_f := 0;
        ELSIF x =- 26054 THEN
            exp_f := 0;
        ELSIF x =- 26053 THEN
            exp_f := 0;
        ELSIF x =- 26052 THEN
            exp_f := 0;
        ELSIF x =- 26051 THEN
            exp_f := 0;
        ELSIF x =- 26050 THEN
            exp_f := 0;
        ELSIF x =- 26049 THEN
            exp_f := 0;
        ELSIF x =- 26048 THEN
            exp_f := 0;
        ELSIF x =- 26047 THEN
            exp_f := 0;
        ELSIF x =- 26046 THEN
            exp_f := 0;
        ELSIF x =- 26045 THEN
            exp_f := 0;
        ELSIF x =- 26044 THEN
            exp_f := 0;
        ELSIF x =- 26043 THEN
            exp_f := 0;
        ELSIF x =- 26042 THEN
            exp_f := 0;
        ELSIF x =- 26041 THEN
            exp_f := 0;
        ELSIF x =- 26040 THEN
            exp_f := 0;
        ELSIF x =- 26039 THEN
            exp_f := 0;
        ELSIF x =- 26038 THEN
            exp_f := 0;
        ELSIF x =- 26037 THEN
            exp_f := 0;
        ELSIF x =- 26036 THEN
            exp_f := 0;
        ELSIF x =- 26035 THEN
            exp_f := 0;
        ELSIF x =- 26034 THEN
            exp_f := 0;
        ELSIF x =- 26033 THEN
            exp_f := 0;
        ELSIF x =- 26032 THEN
            exp_f := 0;
        ELSIF x =- 26031 THEN
            exp_f := 0;
        ELSIF x =- 26030 THEN
            exp_f := 0;
        ELSIF x =- 26029 THEN
            exp_f := 0;
        ELSIF x =- 26028 THEN
            exp_f := 0;
        ELSIF x =- 26027 THEN
            exp_f := 0;
        ELSIF x =- 26026 THEN
            exp_f := 0;
        ELSIF x =- 26025 THEN
            exp_f := 0;
        ELSIF x =- 26024 THEN
            exp_f := 0;
        ELSIF x =- 26023 THEN
            exp_f := 0;
        ELSIF x =- 26022 THEN
            exp_f := 0;
        ELSIF x =- 26021 THEN
            exp_f := 0;
        ELSIF x =- 26020 THEN
            exp_f := 0;
        ELSIF x =- 26019 THEN
            exp_f := 0;
        ELSIF x =- 26018 THEN
            exp_f := 0;
        ELSIF x =- 26017 THEN
            exp_f := 0;
        ELSIF x =- 26016 THEN
            exp_f := 0;
        ELSIF x =- 26015 THEN
            exp_f := 0;
        ELSIF x =- 26014 THEN
            exp_f := 0;
        ELSIF x =- 26013 THEN
            exp_f := 0;
        ELSIF x =- 26012 THEN
            exp_f := 0;
        ELSIF x =- 26011 THEN
            exp_f := 0;
        ELSIF x =- 26010 THEN
            exp_f := 0;
        ELSIF x =- 26009 THEN
            exp_f := 0;
        ELSIF x =- 26008 THEN
            exp_f := 0;
        ELSIF x =- 26007 THEN
            exp_f := 0;
        ELSIF x =- 26006 THEN
            exp_f := 0;
        ELSIF x =- 26005 THEN
            exp_f := 0;
        ELSIF x =- 26004 THEN
            exp_f := 0;
        ELSIF x =- 26003 THEN
            exp_f := 0;
        ELSIF x =- 26002 THEN
            exp_f := 0;
        ELSIF x =- 26001 THEN
            exp_f := 0;
        ELSIF x =- 26000 THEN
            exp_f := 0;
        ELSIF x =- 25999 THEN
            exp_f := 0;
        ELSIF x =- 25998 THEN
            exp_f := 0;
        ELSIF x =- 25997 THEN
            exp_f := 0;
        ELSIF x =- 25996 THEN
            exp_f := 0;
        ELSIF x =- 25995 THEN
            exp_f := 0;
        ELSIF x =- 25994 THEN
            exp_f := 0;
        ELSIF x =- 25993 THEN
            exp_f := 0;
        ELSIF x =- 25992 THEN
            exp_f := 0;
        ELSIF x =- 25991 THEN
            exp_f := 0;
        ELSIF x =- 25990 THEN
            exp_f := 0;
        ELSIF x =- 25989 THEN
            exp_f := 0;
        ELSIF x =- 25988 THEN
            exp_f := 0;
        ELSIF x =- 25987 THEN
            exp_f := 0;
        ELSIF x =- 25986 THEN
            exp_f := 0;
        ELSIF x =- 25985 THEN
            exp_f := 0;
        ELSIF x =- 25984 THEN
            exp_f := 0;
        ELSIF x =- 25983 THEN
            exp_f := 0;
        ELSIF x =- 25982 THEN
            exp_f := 0;
        ELSIF x =- 25981 THEN
            exp_f := 0;
        ELSIF x =- 25980 THEN
            exp_f := 0;
        ELSIF x =- 25979 THEN
            exp_f := 0;
        ELSIF x =- 25978 THEN
            exp_f := 0;
        ELSIF x =- 25977 THEN
            exp_f := 0;
        ELSIF x =- 25976 THEN
            exp_f := 0;
        ELSIF x =- 25975 THEN
            exp_f := 0;
        ELSIF x =- 25974 THEN
            exp_f := 0;
        ELSIF x =- 25973 THEN
            exp_f := 0;
        ELSIF x =- 25972 THEN
            exp_f := 0;
        ELSIF x =- 25971 THEN
            exp_f := 0;
        ELSIF x =- 25970 THEN
            exp_f := 0;
        ELSIF x =- 25969 THEN
            exp_f := 0;
        ELSIF x =- 25968 THEN
            exp_f := 0;
        ELSIF x =- 25967 THEN
            exp_f := 0;
        ELSIF x =- 25966 THEN
            exp_f := 0;
        ELSIF x =- 25965 THEN
            exp_f := 0;
        ELSIF x =- 25964 THEN
            exp_f := 0;
        ELSIF x =- 25963 THEN
            exp_f := 0;
        ELSIF x =- 25962 THEN
            exp_f := 0;
        ELSIF x =- 25961 THEN
            exp_f := 0;
        ELSIF x =- 25960 THEN
            exp_f := 0;
        ELSIF x =- 25959 THEN
            exp_f := 0;
        ELSIF x =- 25958 THEN
            exp_f := 0;
        ELSIF x =- 25957 THEN
            exp_f := 0;
        ELSIF x =- 25956 THEN
            exp_f := 0;
        ELSIF x =- 25955 THEN
            exp_f := 0;
        ELSIF x =- 25954 THEN
            exp_f := 0;
        ELSIF x =- 25953 THEN
            exp_f := 0;
        ELSIF x =- 25952 THEN
            exp_f := 0;
        ELSIF x =- 25951 THEN
            exp_f := 0;
        ELSIF x =- 25950 THEN
            exp_f := 0;
        ELSIF x =- 25949 THEN
            exp_f := 0;
        ELSIF x =- 25948 THEN
            exp_f := 0;
        ELSIF x =- 25947 THEN
            exp_f := 0;
        ELSIF x =- 25946 THEN
            exp_f := 0;
        ELSIF x =- 25945 THEN
            exp_f := 0;
        ELSIF x =- 25944 THEN
            exp_f := 0;
        ELSIF x =- 25943 THEN
            exp_f := 0;
        ELSIF x =- 25942 THEN
            exp_f := 0;
        ELSIF x =- 25941 THEN
            exp_f := 0;
        ELSIF x =- 25940 THEN
            exp_f := 0;
        ELSIF x =- 25939 THEN
            exp_f := 0;
        ELSIF x =- 25938 THEN
            exp_f := 0;
        ELSIF x =- 25937 THEN
            exp_f := 0;
        ELSIF x =- 25936 THEN
            exp_f := 0;
        ELSIF x =- 25935 THEN
            exp_f := 0;
        ELSIF x =- 25934 THEN
            exp_f := 0;
        ELSIF x =- 25933 THEN
            exp_f := 0;
        ELSIF x =- 25932 THEN
            exp_f := 0;
        ELSIF x =- 25931 THEN
            exp_f := 0;
        ELSIF x =- 25930 THEN
            exp_f := 0;
        ELSIF x =- 25929 THEN
            exp_f := 0;
        ELSIF x =- 25928 THEN
            exp_f := 0;
        ELSIF x =- 25927 THEN
            exp_f := 0;
        ELSIF x =- 25926 THEN
            exp_f := 0;
        ELSIF x =- 25925 THEN
            exp_f := 0;
        ELSIF x =- 25924 THEN
            exp_f := 0;
        ELSIF x =- 25923 THEN
            exp_f := 0;
        ELSIF x =- 25922 THEN
            exp_f := 0;
        ELSIF x =- 25921 THEN
            exp_f := 0;
        ELSIF x =- 25920 THEN
            exp_f := 0;
        ELSIF x =- 25919 THEN
            exp_f := 0;
        ELSIF x =- 25918 THEN
            exp_f := 0;
        ELSIF x =- 25917 THEN
            exp_f := 0;
        ELSIF x =- 25916 THEN
            exp_f := 0;
        ELSIF x =- 25915 THEN
            exp_f := 0;
        ELSIF x =- 25914 THEN
            exp_f := 0;
        ELSIF x =- 25913 THEN
            exp_f := 0;
        ELSIF x =- 25912 THEN
            exp_f := 0;
        ELSIF x =- 25911 THEN
            exp_f := 0;
        ELSIF x =- 25910 THEN
            exp_f := 0;
        ELSIF x =- 25909 THEN
            exp_f := 0;
        ELSIF x =- 25908 THEN
            exp_f := 0;
        ELSIF x =- 25907 THEN
            exp_f := 0;
        ELSIF x =- 25906 THEN
            exp_f := 0;
        ELSIF x =- 25905 THEN
            exp_f := 0;
        ELSIF x =- 25904 THEN
            exp_f := 0;
        ELSIF x =- 25903 THEN
            exp_f := 0;
        ELSIF x =- 25902 THEN
            exp_f := 0;
        ELSIF x =- 25901 THEN
            exp_f := 0;
        ELSIF x =- 25900 THEN
            exp_f := 0;
        ELSIF x =- 25899 THEN
            exp_f := 0;
        ELSIF x =- 25898 THEN
            exp_f := 0;
        ELSIF x =- 25897 THEN
            exp_f := 0;
        ELSIF x =- 25896 THEN
            exp_f := 0;
        ELSIF x =- 25895 THEN
            exp_f := 0;
        ELSIF x =- 25894 THEN
            exp_f := 0;
        ELSIF x =- 25893 THEN
            exp_f := 0;
        ELSIF x =- 25892 THEN
            exp_f := 0;
        ELSIF x =- 25891 THEN
            exp_f := 0;
        ELSIF x =- 25890 THEN
            exp_f := 0;
        ELSIF x =- 25889 THEN
            exp_f := 0;
        ELSIF x =- 25888 THEN
            exp_f := 0;
        ELSIF x =- 25887 THEN
            exp_f := 0;
        ELSIF x =- 25886 THEN
            exp_f := 0;
        ELSIF x =- 25885 THEN
            exp_f := 0;
        ELSIF x =- 25884 THEN
            exp_f := 0;
        ELSIF x =- 25883 THEN
            exp_f := 0;
        ELSIF x =- 25882 THEN
            exp_f := 0;
        ELSIF x =- 25881 THEN
            exp_f := 0;
        ELSIF x =- 25880 THEN
            exp_f := 0;
        ELSIF x =- 25879 THEN
            exp_f := 0;
        ELSIF x =- 25878 THEN
            exp_f := 0;
        ELSIF x =- 25877 THEN
            exp_f := 0;
        ELSIF x =- 25876 THEN
            exp_f := 0;
        ELSIF x =- 25875 THEN
            exp_f := 0;
        ELSIF x =- 25874 THEN
            exp_f := 0;
        ELSIF x =- 25873 THEN
            exp_f := 0;
        ELSIF x =- 25872 THEN
            exp_f := 0;
        ELSIF x =- 25871 THEN
            exp_f := 0;
        ELSIF x =- 25870 THEN
            exp_f := 0;
        ELSIF x =- 25869 THEN
            exp_f := 0;
        ELSIF x =- 25868 THEN
            exp_f := 0;
        ELSIF x =- 25867 THEN
            exp_f := 0;
        ELSIF x =- 25866 THEN
            exp_f := 0;
        ELSIF x =- 25865 THEN
            exp_f := 0;
        ELSIF x =- 25864 THEN
            exp_f := 0;
        ELSIF x =- 25863 THEN
            exp_f := 0;
        ELSIF x =- 25862 THEN
            exp_f := 0;
        ELSIF x =- 25861 THEN
            exp_f := 0;
        ELSIF x =- 25860 THEN
            exp_f := 0;
        ELSIF x =- 25859 THEN
            exp_f := 0;
        ELSIF x =- 25858 THEN
            exp_f := 0;
        ELSIF x =- 25857 THEN
            exp_f := 0;
        ELSIF x =- 25856 THEN
            exp_f := 0;
        ELSIF x =- 25855 THEN
            exp_f := 0;
        ELSIF x =- 25854 THEN
            exp_f := 0;
        ELSIF x =- 25853 THEN
            exp_f := 0;
        ELSIF x =- 25852 THEN
            exp_f := 0;
        ELSIF x =- 25851 THEN
            exp_f := 0;
        ELSIF x =- 25850 THEN
            exp_f := 0;
        ELSIF x =- 25849 THEN
            exp_f := 0;
        ELSIF x =- 25848 THEN
            exp_f := 0;
        ELSIF x =- 25847 THEN
            exp_f := 0;
        ELSIF x =- 25846 THEN
            exp_f := 0;
        ELSIF x =- 25845 THEN
            exp_f := 0;
        ELSIF x =- 25844 THEN
            exp_f := 0;
        ELSIF x =- 25843 THEN
            exp_f := 0;
        ELSIF x =- 25842 THEN
            exp_f := 0;
        ELSIF x =- 25841 THEN
            exp_f := 0;
        ELSIF x =- 25840 THEN
            exp_f := 0;
        ELSIF x =- 25839 THEN
            exp_f := 0;
        ELSIF x =- 25838 THEN
            exp_f := 0;
        ELSIF x =- 25837 THEN
            exp_f := 0;
        ELSIF x =- 25836 THEN
            exp_f := 0;
        ELSIF x =- 25835 THEN
            exp_f := 0;
        ELSIF x =- 25834 THEN
            exp_f := 0;
        ELSIF x =- 25833 THEN
            exp_f := 0;
        ELSIF x =- 25832 THEN
            exp_f := 0;
        ELSIF x =- 25831 THEN
            exp_f := 0;
        ELSIF x =- 25830 THEN
            exp_f := 0;
        ELSIF x =- 25829 THEN
            exp_f := 0;
        ELSIF x =- 25828 THEN
            exp_f := 0;
        ELSIF x =- 25827 THEN
            exp_f := 0;
        ELSIF x =- 25826 THEN
            exp_f := 0;
        ELSIF x =- 25825 THEN
            exp_f := 0;
        ELSIF x =- 25824 THEN
            exp_f := 0;
        ELSIF x =- 25823 THEN
            exp_f := 0;
        ELSIF x =- 25822 THEN
            exp_f := 0;
        ELSIF x =- 25821 THEN
            exp_f := 0;
        ELSIF x =- 25820 THEN
            exp_f := 0;
        ELSIF x =- 25819 THEN
            exp_f := 0;
        ELSIF x =- 25818 THEN
            exp_f := 0;
        ELSIF x =- 25817 THEN
            exp_f := 0;
        ELSIF x =- 25816 THEN
            exp_f := 0;
        ELSIF x =- 25815 THEN
            exp_f := 0;
        ELSIF x =- 25814 THEN
            exp_f := 0;
        ELSIF x =- 25813 THEN
            exp_f := 0;
        ELSIF x =- 25812 THEN
            exp_f := 0;
        ELSIF x =- 25811 THEN
            exp_f := 0;
        ELSIF x =- 25810 THEN
            exp_f := 0;
        ELSIF x =- 25809 THEN
            exp_f := 0;
        ELSIF x =- 25808 THEN
            exp_f := 0;
        ELSIF x =- 25807 THEN
            exp_f := 0;
        ELSIF x =- 25806 THEN
            exp_f := 0;
        ELSIF x =- 25805 THEN
            exp_f := 0;
        ELSIF x =- 25804 THEN
            exp_f := 0;
        ELSIF x =- 25803 THEN
            exp_f := 0;
        ELSIF x =- 25802 THEN
            exp_f := 0;
        ELSIF x =- 25801 THEN
            exp_f := 0;
        ELSIF x =- 25800 THEN
            exp_f := 0;
        ELSIF x =- 25799 THEN
            exp_f := 0;
        ELSIF x =- 25798 THEN
            exp_f := 0;
        ELSIF x =- 25797 THEN
            exp_f := 0;
        ELSIF x =- 25796 THEN
            exp_f := 0;
        ELSIF x =- 25795 THEN
            exp_f := 0;
        ELSIF x =- 25794 THEN
            exp_f := 0;
        ELSIF x =- 25793 THEN
            exp_f := 0;
        ELSIF x =- 25792 THEN
            exp_f := 0;
        ELSIF x =- 25791 THEN
            exp_f := 0;
        ELSIF x =- 25790 THEN
            exp_f := 0;
        ELSIF x =- 25789 THEN
            exp_f := 0;
        ELSIF x =- 25788 THEN
            exp_f := 0;
        ELSIF x =- 25787 THEN
            exp_f := 0;
        ELSIF x =- 25786 THEN
            exp_f := 0;
        ELSIF x =- 25785 THEN
            exp_f := 0;
        ELSIF x =- 25784 THEN
            exp_f := 0;
        ELSIF x =- 25783 THEN
            exp_f := 0;
        ELSIF x =- 25782 THEN
            exp_f := 0;
        ELSIF x =- 25781 THEN
            exp_f := 0;
        ELSIF x =- 25780 THEN
            exp_f := 0;
        ELSIF x =- 25779 THEN
            exp_f := 0;
        ELSIF x =- 25778 THEN
            exp_f := 0;
        ELSIF x =- 25777 THEN
            exp_f := 0;
        ELSIF x =- 25776 THEN
            exp_f := 0;
        ELSIF x =- 25775 THEN
            exp_f := 0;
        ELSIF x =- 25774 THEN
            exp_f := 0;
        ELSIF x =- 25773 THEN
            exp_f := 0;
        ELSIF x =- 25772 THEN
            exp_f := 0;
        ELSIF x =- 25771 THEN
            exp_f := 0;
        ELSIF x =- 25770 THEN
            exp_f := 0;
        ELSIF x =- 25769 THEN
            exp_f := 0;
        ELSIF x =- 25768 THEN
            exp_f := 0;
        ELSIF x =- 25767 THEN
            exp_f := 0;
        ELSIF x =- 25766 THEN
            exp_f := 0;
        ELSIF x =- 25765 THEN
            exp_f := 0;
        ELSIF x =- 25764 THEN
            exp_f := 0;
        ELSIF x =- 25763 THEN
            exp_f := 0;
        ELSIF x =- 25762 THEN
            exp_f := 0;
        ELSIF x =- 25761 THEN
            exp_f := 0;
        ELSIF x =- 25760 THEN
            exp_f := 0;
        ELSIF x =- 25759 THEN
            exp_f := 0;
        ELSIF x =- 25758 THEN
            exp_f := 0;
        ELSIF x =- 25757 THEN
            exp_f := 0;
        ELSIF x =- 25756 THEN
            exp_f := 0;
        ELSIF x =- 25755 THEN
            exp_f := 0;
        ELSIF x =- 25754 THEN
            exp_f := 0;
        ELSIF x =- 25753 THEN
            exp_f := 0;
        ELSIF x =- 25752 THEN
            exp_f := 0;
        ELSIF x =- 25751 THEN
            exp_f := 0;
        ELSIF x =- 25750 THEN
            exp_f := 0;
        ELSIF x =- 25749 THEN
            exp_f := 0;
        ELSIF x =- 25748 THEN
            exp_f := 0;
        ELSIF x =- 25747 THEN
            exp_f := 0;
        ELSIF x =- 25746 THEN
            exp_f := 0;
        ELSIF x =- 25745 THEN
            exp_f := 0;
        ELSIF x =- 25744 THEN
            exp_f := 0;
        ELSIF x =- 25743 THEN
            exp_f := 0;
        ELSIF x =- 25742 THEN
            exp_f := 0;
        ELSIF x =- 25741 THEN
            exp_f := 0;
        ELSIF x =- 25740 THEN
            exp_f := 0;
        ELSIF x =- 25739 THEN
            exp_f := 0;
        ELSIF x =- 25738 THEN
            exp_f := 0;
        ELSIF x =- 25737 THEN
            exp_f := 0;
        ELSIF x =- 25736 THEN
            exp_f := 0;
        ELSIF x =- 25735 THEN
            exp_f := 0;
        ELSIF x =- 25734 THEN
            exp_f := 0;
        ELSIF x =- 25733 THEN
            exp_f := 0;
        ELSIF x =- 25732 THEN
            exp_f := 0;
        ELSIF x =- 25731 THEN
            exp_f := 0;
        ELSIF x =- 25730 THEN
            exp_f := 0;
        ELSIF x =- 25729 THEN
            exp_f := 0;
        ELSIF x =- 25728 THEN
            exp_f := 0;
        ELSIF x =- 25727 THEN
            exp_f := 0;
        ELSIF x =- 25726 THEN
            exp_f := 0;
        ELSIF x =- 25725 THEN
            exp_f := 0;
        ELSIF x =- 25724 THEN
            exp_f := 0;
        ELSIF x =- 25723 THEN
            exp_f := 0;
        ELSIF x =- 25722 THEN
            exp_f := 0;
        ELSIF x =- 25721 THEN
            exp_f := 0;
        ELSIF x =- 25720 THEN
            exp_f := 0;
        ELSIF x =- 25719 THEN
            exp_f := 0;
        ELSIF x =- 25718 THEN
            exp_f := 0;
        ELSIF x =- 25717 THEN
            exp_f := 0;
        ELSIF x =- 25716 THEN
            exp_f := 0;
        ELSIF x =- 25715 THEN
            exp_f := 0;
        ELSIF x =- 25714 THEN
            exp_f := 0;
        ELSIF x =- 25713 THEN
            exp_f := 0;
        ELSIF x =- 25712 THEN
            exp_f := 0;
        ELSIF x =- 25711 THEN
            exp_f := 0;
        ELSIF x =- 25710 THEN
            exp_f := 0;
        ELSIF x =- 25709 THEN
            exp_f := 0;
        ELSIF x =- 25708 THEN
            exp_f := 0;
        ELSIF x =- 25707 THEN
            exp_f := 0;
        ELSIF x =- 25706 THEN
            exp_f := 0;
        ELSIF x =- 25705 THEN
            exp_f := 0;
        ELSIF x =- 25704 THEN
            exp_f := 0;
        ELSIF x =- 25703 THEN
            exp_f := 0;
        ELSIF x =- 25702 THEN
            exp_f := 0;
        ELSIF x =- 25701 THEN
            exp_f := 0;
        ELSIF x =- 25700 THEN
            exp_f := 0;
        ELSIF x =- 25699 THEN
            exp_f := 0;
        ELSIF x =- 25698 THEN
            exp_f := 0;
        ELSIF x =- 25697 THEN
            exp_f := 0;
        ELSIF x =- 25696 THEN
            exp_f := 0;
        ELSIF x =- 25695 THEN
            exp_f := 0;
        ELSIF x =- 25694 THEN
            exp_f := 0;
        ELSIF x =- 25693 THEN
            exp_f := 0;
        ELSIF x =- 25692 THEN
            exp_f := 0;
        ELSIF x =- 25691 THEN
            exp_f := 0;
        ELSIF x =- 25690 THEN
            exp_f := 0;
        ELSIF x =- 25689 THEN
            exp_f := 0;
        ELSIF x =- 25688 THEN
            exp_f := 0;
        ELSIF x =- 25687 THEN
            exp_f := 0;
        ELSIF x =- 25686 THEN
            exp_f := 0;
        ELSIF x =- 25685 THEN
            exp_f := 0;
        ELSIF x =- 25684 THEN
            exp_f := 0;
        ELSIF x =- 25683 THEN
            exp_f := 0;
        ELSIF x =- 25682 THEN
            exp_f := 0;
        ELSIF x =- 25681 THEN
            exp_f := 0;
        ELSIF x =- 25680 THEN
            exp_f := 0;
        ELSIF x =- 25679 THEN
            exp_f := 0;
        ELSIF x =- 25678 THEN
            exp_f := 0;
        ELSIF x =- 25677 THEN
            exp_f := 0;
        ELSIF x =- 25676 THEN
            exp_f := 0;
        ELSIF x =- 25675 THEN
            exp_f := 0;
        ELSIF x =- 25674 THEN
            exp_f := 0;
        ELSIF x =- 25673 THEN
            exp_f := 0;
        ELSIF x =- 25672 THEN
            exp_f := 0;
        ELSIF x =- 25671 THEN
            exp_f := 0;
        ELSIF x =- 25670 THEN
            exp_f := 0;
        ELSIF x =- 25669 THEN
            exp_f := 0;
        ELSIF x =- 25668 THEN
            exp_f := 0;
        ELSIF x =- 25667 THEN
            exp_f := 0;
        ELSIF x =- 25666 THEN
            exp_f := 0;
        ELSIF x =- 25665 THEN
            exp_f := 0;
        ELSIF x =- 25664 THEN
            exp_f := 0;
        ELSIF x =- 25663 THEN
            exp_f := 0;
        ELSIF x =- 25662 THEN
            exp_f := 0;
        ELSIF x =- 25661 THEN
            exp_f := 0;
        ELSIF x =- 25660 THEN
            exp_f := 0;
        ELSIF x =- 25659 THEN
            exp_f := 0;
        ELSIF x =- 25658 THEN
            exp_f := 0;
        ELSIF x =- 25657 THEN
            exp_f := 0;
        ELSIF x =- 25656 THEN
            exp_f := 0;
        ELSIF x =- 25655 THEN
            exp_f := 0;
        ELSIF x =- 25654 THEN
            exp_f := 0;
        ELSIF x =- 25653 THEN
            exp_f := 0;
        ELSIF x =- 25652 THEN
            exp_f := 0;
        ELSIF x =- 25651 THEN
            exp_f := 0;
        ELSIF x =- 25650 THEN
            exp_f := 0;
        ELSIF x =- 25649 THEN
            exp_f := 0;
        ELSIF x =- 25648 THEN
            exp_f := 0;
        ELSIF x =- 25647 THEN
            exp_f := 0;
        ELSIF x =- 25646 THEN
            exp_f := 0;
        ELSIF x =- 25645 THEN
            exp_f := 0;
        ELSIF x =- 25644 THEN
            exp_f := 0;
        ELSIF x =- 25643 THEN
            exp_f := 0;
        ELSIF x =- 25642 THEN
            exp_f := 0;
        ELSIF x =- 25641 THEN
            exp_f := 0;
        ELSIF x =- 25640 THEN
            exp_f := 0;
        ELSIF x =- 25639 THEN
            exp_f := 0;
        ELSIF x =- 25638 THEN
            exp_f := 0;
        ELSIF x =- 25637 THEN
            exp_f := 0;
        ELSIF x =- 25636 THEN
            exp_f := 0;
        ELSIF x =- 25635 THEN
            exp_f := 0;
        ELSIF x =- 25634 THEN
            exp_f := 0;
        ELSIF x =- 25633 THEN
            exp_f := 0;
        ELSIF x =- 25632 THEN
            exp_f := 0;
        ELSIF x =- 25631 THEN
            exp_f := 0;
        ELSIF x =- 25630 THEN
            exp_f := 0;
        ELSIF x =- 25629 THEN
            exp_f := 0;
        ELSIF x =- 25628 THEN
            exp_f := 0;
        ELSIF x =- 25627 THEN
            exp_f := 0;
        ELSIF x =- 25626 THEN
            exp_f := 0;
        ELSIF x =- 25625 THEN
            exp_f := 0;
        ELSIF x =- 25624 THEN
            exp_f := 0;
        ELSIF x =- 25623 THEN
            exp_f := 0;
        ELSIF x =- 25622 THEN
            exp_f := 0;
        ELSIF x =- 25621 THEN
            exp_f := 0;
        ELSIF x =- 25620 THEN
            exp_f := 0;
        ELSIF x =- 25619 THEN
            exp_f := 0;
        ELSIF x =- 25618 THEN
            exp_f := 0;
        ELSIF x =- 25617 THEN
            exp_f := 0;
        ELSIF x =- 25616 THEN
            exp_f := 0;
        ELSIF x =- 25615 THEN
            exp_f := 0;
        ELSIF x =- 25614 THEN
            exp_f := 0;
        ELSIF x =- 25613 THEN
            exp_f := 0;
        ELSIF x =- 25612 THEN
            exp_f := 0;
        ELSIF x =- 25611 THEN
            exp_f := 0;
        ELSIF x =- 25610 THEN
            exp_f := 0;
        ELSIF x =- 25609 THEN
            exp_f := 0;
        ELSIF x =- 25608 THEN
            exp_f := 0;
        ELSIF x =- 25607 THEN
            exp_f := 0;
        ELSIF x =- 25606 THEN
            exp_f := 0;
        ELSIF x =- 25605 THEN
            exp_f := 0;
        ELSIF x =- 25604 THEN
            exp_f := 0;
        ELSIF x =- 25603 THEN
            exp_f := 0;
        ELSIF x =- 25602 THEN
            exp_f := 0;
        ELSIF x =- 25601 THEN
            exp_f := 0;
        ELSIF x =- 25600 THEN
            exp_f := 0;
        ELSIF x =- 25599 THEN
            exp_f := 0;
        ELSIF x =- 25598 THEN
            exp_f := 0;
        ELSIF x =- 25597 THEN
            exp_f := 0;
        ELSIF x =- 25596 THEN
            exp_f := 0;
        ELSIF x =- 25595 THEN
            exp_f := 0;
        ELSIF x =- 25594 THEN
            exp_f := 0;
        ELSIF x =- 25593 THEN
            exp_f := 0;
        ELSIF x =- 25592 THEN
            exp_f := 0;
        ELSIF x =- 25591 THEN
            exp_f := 0;
        ELSIF x =- 25590 THEN
            exp_f := 0;
        ELSIF x =- 25589 THEN
            exp_f := 0;
        ELSIF x =- 25588 THEN
            exp_f := 0;
        ELSIF x =- 25587 THEN
            exp_f := 0;
        ELSIF x =- 25586 THEN
            exp_f := 0;
        ELSIF x =- 25585 THEN
            exp_f := 0;
        ELSIF x =- 25584 THEN
            exp_f := 0;
        ELSIF x =- 25583 THEN
            exp_f := 0;
        ELSIF x =- 25582 THEN
            exp_f := 0;
        ELSIF x =- 25581 THEN
            exp_f := 0;
        ELSIF x =- 25580 THEN
            exp_f := 0;
        ELSIF x =- 25579 THEN
            exp_f := 0;
        ELSIF x =- 25578 THEN
            exp_f := 0;
        ELSIF x =- 25577 THEN
            exp_f := 0;
        ELSIF x =- 25576 THEN
            exp_f := 0;
        ELSIF x =- 25575 THEN
            exp_f := 0;
        ELSIF x =- 25574 THEN
            exp_f := 0;
        ELSIF x =- 25573 THEN
            exp_f := 0;
        ELSIF x =- 25572 THEN
            exp_f := 0;
        ELSIF x =- 25571 THEN
            exp_f := 0;
        ELSIF x =- 25570 THEN
            exp_f := 0;
        ELSIF x =- 25569 THEN
            exp_f := 0;
        ELSIF x =- 25568 THEN
            exp_f := 0;
        ELSIF x =- 25567 THEN
            exp_f := 0;
        ELSIF x =- 25566 THEN
            exp_f := 0;
        ELSIF x =- 25565 THEN
            exp_f := 0;
        ELSIF x =- 25564 THEN
            exp_f := 0;
        ELSIF x =- 25563 THEN
            exp_f := 0;
        ELSIF x =- 25562 THEN
            exp_f := 0;
        ELSIF x =- 25561 THEN
            exp_f := 0;
        ELSIF x =- 25560 THEN
            exp_f := 0;
        ELSIF x =- 25559 THEN
            exp_f := 0;
        ELSIF x =- 25558 THEN
            exp_f := 0;
        ELSIF x =- 25557 THEN
            exp_f := 0;
        ELSIF x =- 25556 THEN
            exp_f := 0;
        ELSIF x =- 25555 THEN
            exp_f := 0;
        ELSIF x =- 25554 THEN
            exp_f := 0;
        ELSIF x =- 25553 THEN
            exp_f := 0;
        ELSIF x =- 25552 THEN
            exp_f := 0;
        ELSIF x =- 25551 THEN
            exp_f := 0;
        ELSIF x =- 25550 THEN
            exp_f := 0;
        ELSIF x =- 25549 THEN
            exp_f := 0;
        ELSIF x =- 25548 THEN
            exp_f := 0;
        ELSIF x =- 25547 THEN
            exp_f := 0;
        ELSIF x =- 25546 THEN
            exp_f := 0;
        ELSIF x =- 25545 THEN
            exp_f := 0;
        ELSIF x =- 25544 THEN
            exp_f := 0;
        ELSIF x =- 25543 THEN
            exp_f := 0;
        ELSIF x =- 25542 THEN
            exp_f := 0;
        ELSIF x =- 25541 THEN
            exp_f := 0;
        ELSIF x =- 25540 THEN
            exp_f := 0;
        ELSIF x =- 25539 THEN
            exp_f := 0;
        ELSIF x =- 25538 THEN
            exp_f := 0;
        ELSIF x =- 25537 THEN
            exp_f := 0;
        ELSIF x =- 25536 THEN
            exp_f := 0;
        ELSIF x =- 25535 THEN
            exp_f := 0;
        ELSIF x =- 25534 THEN
            exp_f := 0;
        ELSIF x =- 25533 THEN
            exp_f := 0;
        ELSIF x =- 25532 THEN
            exp_f := 0;
        ELSIF x =- 25531 THEN
            exp_f := 0;
        ELSIF x =- 25530 THEN
            exp_f := 0;
        ELSIF x =- 25529 THEN
            exp_f := 0;
        ELSIF x =- 25528 THEN
            exp_f := 0;
        ELSIF x =- 25527 THEN
            exp_f := 0;
        ELSIF x =- 25526 THEN
            exp_f := 0;
        ELSIF x =- 25525 THEN
            exp_f := 0;
        ELSIF x =- 25524 THEN
            exp_f := 0;
        ELSIF x =- 25523 THEN
            exp_f := 0;
        ELSIF x =- 25522 THEN
            exp_f := 0;
        ELSIF x =- 25521 THEN
            exp_f := 0;
        ELSIF x =- 25520 THEN
            exp_f := 0;
        ELSIF x =- 25519 THEN
            exp_f := 0;
        ELSIF x =- 25518 THEN
            exp_f := 0;
        ELSIF x =- 25517 THEN
            exp_f := 0;
        ELSIF x =- 25516 THEN
            exp_f := 0;
        ELSIF x =- 25515 THEN
            exp_f := 0;
        ELSIF x =- 25514 THEN
            exp_f := 0;
        ELSIF x =- 25513 THEN
            exp_f := 0;
        ELSIF x =- 25512 THEN
            exp_f := 0;
        ELSIF x =- 25511 THEN
            exp_f := 0;
        ELSIF x =- 25510 THEN
            exp_f := 0;
        ELSIF x =- 25509 THEN
            exp_f := 0;
        ELSIF x =- 25508 THEN
            exp_f := 0;
        ELSIF x =- 25507 THEN
            exp_f := 0;
        ELSIF x =- 25506 THEN
            exp_f := 0;
        ELSIF x =- 25505 THEN
            exp_f := 0;
        ELSIF x =- 25504 THEN
            exp_f := 0;
        ELSIF x =- 25503 THEN
            exp_f := 0;
        ELSIF x =- 25502 THEN
            exp_f := 0;
        ELSIF x =- 25501 THEN
            exp_f := 0;
        ELSIF x =- 25500 THEN
            exp_f := 0;
        ELSIF x =- 25499 THEN
            exp_f := 0;
        ELSIF x =- 25498 THEN
            exp_f := 0;
        ELSIF x =- 25497 THEN
            exp_f := 0;
        ELSIF x =- 25496 THEN
            exp_f := 0;
        ELSIF x =- 25495 THEN
            exp_f := 0;
        ELSIF x =- 25494 THEN
            exp_f := 0;
        ELSIF x =- 25493 THEN
            exp_f := 0;
        ELSIF x =- 25492 THEN
            exp_f := 0;
        ELSIF x =- 25491 THEN
            exp_f := 0;
        ELSIF x =- 25490 THEN
            exp_f := 0;
        ELSIF x =- 25489 THEN
            exp_f := 0;
        ELSIF x =- 25488 THEN
            exp_f := 0;
        ELSIF x =- 25487 THEN
            exp_f := 0;
        ELSIF x =- 25486 THEN
            exp_f := 0;
        ELSIF x =- 25485 THEN
            exp_f := 0;
        ELSIF x =- 25484 THEN
            exp_f := 0;
        ELSIF x =- 25483 THEN
            exp_f := 0;
        ELSIF x =- 25482 THEN
            exp_f := 0;
        ELSIF x =- 25481 THEN
            exp_f := 0;
        ELSIF x =- 25480 THEN
            exp_f := 0;
        ELSIF x =- 25479 THEN
            exp_f := 0;
        ELSIF x =- 25478 THEN
            exp_f := 0;
        ELSIF x =- 25477 THEN
            exp_f := 0;
        ELSIF x =- 25476 THEN
            exp_f := 0;
        ELSIF x =- 25475 THEN
            exp_f := 0;
        ELSIF x =- 25474 THEN
            exp_f := 0;
        ELSIF x =- 25473 THEN
            exp_f := 0;
        ELSIF x =- 25472 THEN
            exp_f := 0;
        ELSIF x =- 25471 THEN
            exp_f := 0;
        ELSIF x =- 25470 THEN
            exp_f := 0;
        ELSIF x =- 25469 THEN
            exp_f := 0;
        ELSIF x =- 25468 THEN
            exp_f := 0;
        ELSIF x =- 25467 THEN
            exp_f := 0;
        ELSIF x =- 25466 THEN
            exp_f := 0;
        ELSIF x =- 25465 THEN
            exp_f := 0;
        ELSIF x =- 25464 THEN
            exp_f := 0;
        ELSIF x =- 25463 THEN
            exp_f := 0;
        ELSIF x =- 25462 THEN
            exp_f := 0;
        ELSIF x =- 25461 THEN
            exp_f := 0;
        ELSIF x =- 25460 THEN
            exp_f := 0;
        ELSIF x =- 25459 THEN
            exp_f := 0;
        ELSIF x =- 25458 THEN
            exp_f := 0;
        ELSIF x =- 25457 THEN
            exp_f := 0;
        ELSIF x =- 25456 THEN
            exp_f := 0;
        ELSIF x =- 25455 THEN
            exp_f := 0;
        ELSIF x =- 25454 THEN
            exp_f := 0;
        ELSIF x =- 25453 THEN
            exp_f := 0;
        ELSIF x =- 25452 THEN
            exp_f := 0;
        ELSIF x =- 25451 THEN
            exp_f := 0;
        ELSIF x =- 25450 THEN
            exp_f := 0;
        ELSIF x =- 25449 THEN
            exp_f := 0;
        ELSIF x =- 25448 THEN
            exp_f := 0;
        ELSIF x =- 25447 THEN
            exp_f := 0;
        ELSIF x =- 25446 THEN
            exp_f := 0;
        ELSIF x =- 25445 THEN
            exp_f := 0;
        ELSIF x =- 25444 THEN
            exp_f := 0;
        ELSIF x =- 25443 THEN
            exp_f := 0;
        ELSIF x =- 25442 THEN
            exp_f := 0;
        ELSIF x =- 25441 THEN
            exp_f := 0;
        ELSIF x =- 25440 THEN
            exp_f := 0;
        ELSIF x =- 25439 THEN
            exp_f := 0;
        ELSIF x =- 25438 THEN
            exp_f := 0;
        ELSIF x =- 25437 THEN
            exp_f := 0;
        ELSIF x =- 25436 THEN
            exp_f := 0;
        ELSIF x =- 25435 THEN
            exp_f := 0;
        ELSIF x =- 25434 THEN
            exp_f := 0;
        ELSIF x =- 25433 THEN
            exp_f := 0;
        ELSIF x =- 25432 THEN
            exp_f := 0;
        ELSIF x =- 25431 THEN
            exp_f := 0;
        ELSIF x =- 25430 THEN
            exp_f := 0;
        ELSIF x =- 25429 THEN
            exp_f := 0;
        ELSIF x =- 25428 THEN
            exp_f := 0;
        ELSIF x =- 25427 THEN
            exp_f := 0;
        ELSIF x =- 25426 THEN
            exp_f := 0;
        ELSIF x =- 25425 THEN
            exp_f := 0;
        ELSIF x =- 25424 THEN
            exp_f := 0;
        ELSIF x =- 25423 THEN
            exp_f := 0;
        ELSIF x =- 25422 THEN
            exp_f := 0;
        ELSIF x =- 25421 THEN
            exp_f := 0;
        ELSIF x =- 25420 THEN
            exp_f := 0;
        ELSIF x =- 25419 THEN
            exp_f := 0;
        ELSIF x =- 25418 THEN
            exp_f := 0;
        ELSIF x =- 25417 THEN
            exp_f := 0;
        ELSIF x =- 25416 THEN
            exp_f := 0;
        ELSIF x =- 25415 THEN
            exp_f := 0;
        ELSIF x =- 25414 THEN
            exp_f := 0;
        ELSIF x =- 25413 THEN
            exp_f := 0;
        ELSIF x =- 25412 THEN
            exp_f := 0;
        ELSIF x =- 25411 THEN
            exp_f := 0;
        ELSIF x =- 25410 THEN
            exp_f := 0;
        ELSIF x =- 25409 THEN
            exp_f := 0;
        ELSIF x =- 25408 THEN
            exp_f := 0;
        ELSIF x =- 25407 THEN
            exp_f := 0;
        ELSIF x =- 25406 THEN
            exp_f := 0;
        ELSIF x =- 25405 THEN
            exp_f := 0;
        ELSIF x =- 25404 THEN
            exp_f := 0;
        ELSIF x =- 25403 THEN
            exp_f := 0;
        ELSIF x =- 25402 THEN
            exp_f := 0;
        ELSIF x =- 25401 THEN
            exp_f := 0;
        ELSIF x =- 25400 THEN
            exp_f := 0;
        ELSIF x =- 25399 THEN
            exp_f := 0;
        ELSIF x =- 25398 THEN
            exp_f := 0;
        ELSIF x =- 25397 THEN
            exp_f := 0;
        ELSIF x =- 25396 THEN
            exp_f := 0;
        ELSIF x =- 25395 THEN
            exp_f := 0;
        ELSIF x =- 25394 THEN
            exp_f := 0;
        ELSIF x =- 25393 THEN
            exp_f := 0;
        ELSIF x =- 25392 THEN
            exp_f := 0;
        ELSIF x =- 25391 THEN
            exp_f := 0;
        ELSIF x =- 25390 THEN
            exp_f := 0;
        ELSIF x =- 25389 THEN
            exp_f := 0;
        ELSIF x =- 25388 THEN
            exp_f := 0;
        ELSIF x =- 25387 THEN
            exp_f := 0;
        ELSIF x =- 25386 THEN
            exp_f := 0;
        ELSIF x =- 25385 THEN
            exp_f := 0;
        ELSIF x =- 25384 THEN
            exp_f := 0;
        ELSIF x =- 25383 THEN
            exp_f := 0;
        ELSIF x =- 25382 THEN
            exp_f := 0;
        ELSIF x =- 25381 THEN
            exp_f := 0;
        ELSIF x =- 25380 THEN
            exp_f := 0;
        ELSIF x =- 25379 THEN
            exp_f := 0;
        ELSIF x =- 25378 THEN
            exp_f := 0;
        ELSIF x =- 25377 THEN
            exp_f := 0;
        ELSIF x =- 25376 THEN
            exp_f := 0;
        ELSIF x =- 25375 THEN
            exp_f := 0;
        ELSIF x =- 25374 THEN
            exp_f := 0;
        ELSIF x =- 25373 THEN
            exp_f := 0;
        ELSIF x =- 25372 THEN
            exp_f := 0;
        ELSIF x =- 25371 THEN
            exp_f := 0;
        ELSIF x =- 25370 THEN
            exp_f := 0;
        ELSIF x =- 25369 THEN
            exp_f := 0;
        ELSIF x =- 25368 THEN
            exp_f := 0;
        ELSIF x =- 25367 THEN
            exp_f := 0;
        ELSIF x =- 25366 THEN
            exp_f := 0;
        ELSIF x =- 25365 THEN
            exp_f := 0;
        ELSIF x =- 25364 THEN
            exp_f := 0;
        ELSIF x =- 25363 THEN
            exp_f := 0;
        ELSIF x =- 25362 THEN
            exp_f := 0;
        ELSIF x =- 25361 THEN
            exp_f := 0;
        ELSIF x =- 25360 THEN
            exp_f := 0;
        ELSIF x =- 25359 THEN
            exp_f := 0;
        ELSIF x =- 25358 THEN
            exp_f := 0;
        ELSIF x =- 25357 THEN
            exp_f := 0;
        ELSIF x =- 25356 THEN
            exp_f := 0;
        ELSIF x =- 25355 THEN
            exp_f := 0;
        ELSIF x =- 25354 THEN
            exp_f := 0;
        ELSIF x =- 25353 THEN
            exp_f := 0;
        ELSIF x =- 25352 THEN
            exp_f := 0;
        ELSIF x =- 25351 THEN
            exp_f := 0;
        ELSIF x =- 25350 THEN
            exp_f := 0;
        ELSIF x =- 25349 THEN
            exp_f := 0;
        ELSIF x =- 25348 THEN
            exp_f := 0;
        ELSIF x =- 25347 THEN
            exp_f := 0;
        ELSIF x =- 25346 THEN
            exp_f := 0;
        ELSIF x =- 25345 THEN
            exp_f := 0;
        ELSIF x =- 25344 THEN
            exp_f := 0;
        ELSIF x =- 25343 THEN
            exp_f := 0;
        ELSIF x =- 25342 THEN
            exp_f := 0;
        ELSIF x =- 25341 THEN
            exp_f := 0;
        ELSIF x =- 25340 THEN
            exp_f := 0;
        ELSIF x =- 25339 THEN
            exp_f := 0;
        ELSIF x =- 25338 THEN
            exp_f := 0;
        ELSIF x =- 25337 THEN
            exp_f := 0;
        ELSIF x =- 25336 THEN
            exp_f := 0;
        ELSIF x =- 25335 THEN
            exp_f := 0;
        ELSIF x =- 25334 THEN
            exp_f := 0;
        ELSIF x =- 25333 THEN
            exp_f := 0;
        ELSIF x =- 25332 THEN
            exp_f := 0;
        ELSIF x =- 25331 THEN
            exp_f := 0;
        ELSIF x =- 25330 THEN
            exp_f := 0;
        ELSIF x =- 25329 THEN
            exp_f := 0;
        ELSIF x =- 25328 THEN
            exp_f := 0;
        ELSIF x =- 25327 THEN
            exp_f := 0;
        ELSIF x =- 25326 THEN
            exp_f := 0;
        ELSIF x =- 25325 THEN
            exp_f := 0;
        ELSIF x =- 25324 THEN
            exp_f := 0;
        ELSIF x =- 25323 THEN
            exp_f := 0;
        ELSIF x =- 25322 THEN
            exp_f := 0;
        ELSIF x =- 25321 THEN
            exp_f := 0;
        ELSIF x =- 25320 THEN
            exp_f := 0;
        ELSIF x =- 25319 THEN
            exp_f := 0;
        ELSIF x =- 25318 THEN
            exp_f := 0;
        ELSIF x =- 25317 THEN
            exp_f := 0;
        ELSIF x =- 25316 THEN
            exp_f := 0;
        ELSIF x =- 25315 THEN
            exp_f := 0;
        ELSIF x =- 25314 THEN
            exp_f := 0;
        ELSIF x =- 25313 THEN
            exp_f := 0;
        ELSIF x =- 25312 THEN
            exp_f := 0;
        ELSIF x =- 25311 THEN
            exp_f := 0;
        ELSIF x =- 25310 THEN
            exp_f := 0;
        ELSIF x =- 25309 THEN
            exp_f := 0;
        ELSIF x =- 25308 THEN
            exp_f := 0;
        ELSIF x =- 25307 THEN
            exp_f := 0;
        ELSIF x =- 25306 THEN
            exp_f := 0;
        ELSIF x =- 25305 THEN
            exp_f := 0;
        ELSIF x =- 25304 THEN
            exp_f := 0;
        ELSIF x =- 25303 THEN
            exp_f := 0;
        ELSIF x =- 25302 THEN
            exp_f := 0;
        ELSIF x =- 25301 THEN
            exp_f := 0;
        ELSIF x =- 25300 THEN
            exp_f := 0;
        ELSIF x =- 25299 THEN
            exp_f := 0;
        ELSIF x =- 25298 THEN
            exp_f := 0;
        ELSIF x =- 25297 THEN
            exp_f := 0;
        ELSIF x =- 25296 THEN
            exp_f := 0;
        ELSIF x =- 25295 THEN
            exp_f := 0;
        ELSIF x =- 25294 THEN
            exp_f := 0;
        ELSIF x =- 25293 THEN
            exp_f := 0;
        ELSIF x =- 25292 THEN
            exp_f := 0;
        ELSIF x =- 25291 THEN
            exp_f := 0;
        ELSIF x =- 25290 THEN
            exp_f := 0;
        ELSIF x =- 25289 THEN
            exp_f := 0;
        ELSIF x =- 25288 THEN
            exp_f := 0;
        ELSIF x =- 25287 THEN
            exp_f := 0;
        ELSIF x =- 25286 THEN
            exp_f := 0;
        ELSIF x =- 25285 THEN
            exp_f := 0;
        ELSIF x =- 25284 THEN
            exp_f := 0;
        ELSIF x =- 25283 THEN
            exp_f := 0;
        ELSIF x =- 25282 THEN
            exp_f := 0;
        ELSIF x =- 25281 THEN
            exp_f := 0;
        ELSIF x =- 25280 THEN
            exp_f := 0;
        ELSIF x =- 25279 THEN
            exp_f := 0;
        ELSIF x =- 25278 THEN
            exp_f := 0;
        ELSIF x =- 25277 THEN
            exp_f := 0;
        ELSIF x =- 25276 THEN
            exp_f := 0;
        ELSIF x =- 25275 THEN
            exp_f := 0;
        ELSIF x =- 25274 THEN
            exp_f := 0;
        ELSIF x =- 25273 THEN
            exp_f := 0;
        ELSIF x =- 25272 THEN
            exp_f := 0;
        ELSIF x =- 25271 THEN
            exp_f := 0;
        ELSIF x =- 25270 THEN
            exp_f := 0;
        ELSIF x =- 25269 THEN
            exp_f := 0;
        ELSIF x =- 25268 THEN
            exp_f := 0;
        ELSIF x =- 25267 THEN
            exp_f := 0;
        ELSIF x =- 25266 THEN
            exp_f := 0;
        ELSIF x =- 25265 THEN
            exp_f := 0;
        ELSIF x =- 25264 THEN
            exp_f := 0;
        ELSIF x =- 25263 THEN
            exp_f := 0;
        ELSIF x =- 25262 THEN
            exp_f := 0;
        ELSIF x =- 25261 THEN
            exp_f := 0;
        ELSIF x =- 25260 THEN
            exp_f := 0;
        ELSIF x =- 25259 THEN
            exp_f := 0;
        ELSIF x =- 25258 THEN
            exp_f := 0;
        ELSIF x =- 25257 THEN
            exp_f := 0;
        ELSIF x =- 25256 THEN
            exp_f := 0;
        ELSIF x =- 25255 THEN
            exp_f := 0;
        ELSIF x =- 25254 THEN
            exp_f := 0;
        ELSIF x =- 25253 THEN
            exp_f := 0;
        ELSIF x =- 25252 THEN
            exp_f := 0;
        ELSIF x =- 25251 THEN
            exp_f := 0;
        ELSIF x =- 25250 THEN
            exp_f := 0;
        ELSIF x =- 25249 THEN
            exp_f := 0;
        ELSIF x =- 25248 THEN
            exp_f := 0;
        ELSIF x =- 25247 THEN
            exp_f := 0;
        ELSIF x =- 25246 THEN
            exp_f := 0;
        ELSIF x =- 25245 THEN
            exp_f := 0;
        ELSIF x =- 25244 THEN
            exp_f := 0;
        ELSIF x =- 25243 THEN
            exp_f := 0;
        ELSIF x =- 25242 THEN
            exp_f := 0;
        ELSIF x =- 25241 THEN
            exp_f := 0;
        ELSIF x =- 25240 THEN
            exp_f := 0;
        ELSIF x =- 25239 THEN
            exp_f := 0;
        ELSIF x =- 25238 THEN
            exp_f := 0;
        ELSIF x =- 25237 THEN
            exp_f := 0;
        ELSIF x =- 25236 THEN
            exp_f := 0;
        ELSIF x =- 25235 THEN
            exp_f := 0;
        ELSIF x =- 25234 THEN
            exp_f := 0;
        ELSIF x =- 25233 THEN
            exp_f := 0;
        ELSIF x =- 25232 THEN
            exp_f := 0;
        ELSIF x =- 25231 THEN
            exp_f := 0;
        ELSIF x =- 25230 THEN
            exp_f := 0;
        ELSIF x =- 25229 THEN
            exp_f := 0;
        ELSIF x =- 25228 THEN
            exp_f := 0;
        ELSIF x =- 25227 THEN
            exp_f := 0;
        ELSIF x =- 25226 THEN
            exp_f := 0;
        ELSIF x =- 25225 THEN
            exp_f := 0;
        ELSIF x =- 25224 THEN
            exp_f := 0;
        ELSIF x =- 25223 THEN
            exp_f := 0;
        ELSIF x =- 25222 THEN
            exp_f := 0;
        ELSIF x =- 25221 THEN
            exp_f := 0;
        ELSIF x =- 25220 THEN
            exp_f := 0;
        ELSIF x =- 25219 THEN
            exp_f := 0;
        ELSIF x =- 25218 THEN
            exp_f := 0;
        ELSIF x =- 25217 THEN
            exp_f := 0;
        ELSIF x =- 25216 THEN
            exp_f := 0;
        ELSIF x =- 25215 THEN
            exp_f := 0;
        ELSIF x =- 25214 THEN
            exp_f := 0;
        ELSIF x =- 25213 THEN
            exp_f := 0;
        ELSIF x =- 25212 THEN
            exp_f := 0;
        ELSIF x =- 25211 THEN
            exp_f := 0;
        ELSIF x =- 25210 THEN
            exp_f := 0;
        ELSIF x =- 25209 THEN
            exp_f := 0;
        ELSIF x =- 25208 THEN
            exp_f := 0;
        ELSIF x =- 25207 THEN
            exp_f := 0;
        ELSIF x =- 25206 THEN
            exp_f := 0;
        ELSIF x =- 25205 THEN
            exp_f := 0;
        ELSIF x =- 25204 THEN
            exp_f := 0;
        ELSIF x =- 25203 THEN
            exp_f := 0;
        ELSIF x =- 25202 THEN
            exp_f := 0;
        ELSIF x =- 25201 THEN
            exp_f := 0;
        ELSIF x =- 25200 THEN
            exp_f := 0;
        ELSIF x =- 25199 THEN
            exp_f := 0;
        ELSIF x =- 25198 THEN
            exp_f := 0;
        ELSIF x =- 25197 THEN
            exp_f := 0;
        ELSIF x =- 25196 THEN
            exp_f := 0;
        ELSIF x =- 25195 THEN
            exp_f := 0;
        ELSIF x =- 25194 THEN
            exp_f := 0;
        ELSIF x =- 25193 THEN
            exp_f := 0;
        ELSIF x =- 25192 THEN
            exp_f := 0;
        ELSIF x =- 25191 THEN
            exp_f := 0;
        ELSIF x =- 25190 THEN
            exp_f := 0;
        ELSIF x =- 25189 THEN
            exp_f := 0;
        ELSIF x =- 25188 THEN
            exp_f := 0;
        ELSIF x =- 25187 THEN
            exp_f := 0;
        ELSIF x =- 25186 THEN
            exp_f := 0;
        ELSIF x =- 25185 THEN
            exp_f := 0;
        ELSIF x =- 25184 THEN
            exp_f := 0;
        ELSIF x =- 25183 THEN
            exp_f := 0;
        ELSIF x =- 25182 THEN
            exp_f := 0;
        ELSIF x =- 25181 THEN
            exp_f := 0;
        ELSIF x =- 25180 THEN
            exp_f := 0;
        ELSIF x =- 25179 THEN
            exp_f := 0;
        ELSIF x =- 25178 THEN
            exp_f := 0;
        ELSIF x =- 25177 THEN
            exp_f := 0;
        ELSIF x =- 25176 THEN
            exp_f := 0;
        ELSIF x =- 25175 THEN
            exp_f := 0;
        ELSIF x =- 25174 THEN
            exp_f := 0;
        ELSIF x =- 25173 THEN
            exp_f := 0;
        ELSIF x =- 25172 THEN
            exp_f := 0;
        ELSIF x =- 25171 THEN
            exp_f := 0;
        ELSIF x =- 25170 THEN
            exp_f := 0;
        ELSIF x =- 25169 THEN
            exp_f := 0;
        ELSIF x =- 25168 THEN
            exp_f := 0;
        ELSIF x =- 25167 THEN
            exp_f := 0;
        ELSIF x =- 25166 THEN
            exp_f := 0;
        ELSIF x =- 25165 THEN
            exp_f := 0;
        ELSIF x =- 25164 THEN
            exp_f := 0;
        ELSIF x =- 25163 THEN
            exp_f := 0;
        ELSIF x =- 25162 THEN
            exp_f := 0;
        ELSIF x =- 25161 THEN
            exp_f := 0;
        ELSIF x =- 25160 THEN
            exp_f := 0;
        ELSIF x =- 25159 THEN
            exp_f := 0;
        ELSIF x =- 25158 THEN
            exp_f := 0;
        ELSIF x =- 25157 THEN
            exp_f := 0;
        ELSIF x =- 25156 THEN
            exp_f := 0;
        ELSIF x =- 25155 THEN
            exp_f := 0;
        ELSIF x =- 25154 THEN
            exp_f := 0;
        ELSIF x =- 25153 THEN
            exp_f := 0;
        ELSIF x =- 25152 THEN
            exp_f := 0;
        ELSIF x =- 25151 THEN
            exp_f := 0;
        ELSIF x =- 25150 THEN
            exp_f := 0;
        ELSIF x =- 25149 THEN
            exp_f := 0;
        ELSIF x =- 25148 THEN
            exp_f := 0;
        ELSIF x =- 25147 THEN
            exp_f := 0;
        ELSIF x =- 25146 THEN
            exp_f := 0;
        ELSIF x =- 25145 THEN
            exp_f := 0;
        ELSIF x =- 25144 THEN
            exp_f := 0;
        ELSIF x =- 25143 THEN
            exp_f := 0;
        ELSIF x =- 25142 THEN
            exp_f := 0;
        ELSIF x =- 25141 THEN
            exp_f := 0;
        ELSIF x =- 25140 THEN
            exp_f := 0;
        ELSIF x =- 25139 THEN
            exp_f := 0;
        ELSIF x =- 25138 THEN
            exp_f := 0;
        ELSIF x =- 25137 THEN
            exp_f := 0;
        ELSIF x =- 25136 THEN
            exp_f := 0;
        ELSIF x =- 25135 THEN
            exp_f := 0;
        ELSIF x =- 25134 THEN
            exp_f := 0;
        ELSIF x =- 25133 THEN
            exp_f := 0;
        ELSIF x =- 25132 THEN
            exp_f := 0;
        ELSIF x =- 25131 THEN
            exp_f := 0;
        ELSIF x =- 25130 THEN
            exp_f := 0;
        ELSIF x =- 25129 THEN
            exp_f := 0;
        ELSIF x =- 25128 THEN
            exp_f := 0;
        ELSIF x =- 25127 THEN
            exp_f := 0;
        ELSIF x =- 25126 THEN
            exp_f := 0;
        ELSIF x =- 25125 THEN
            exp_f := 0;
        ELSIF x =- 25124 THEN
            exp_f := 0;
        ELSIF x =- 25123 THEN
            exp_f := 0;
        ELSIF x =- 25122 THEN
            exp_f := 0;
        ELSIF x =- 25121 THEN
            exp_f := 0;
        ELSIF x =- 25120 THEN
            exp_f := 0;
        ELSIF x =- 25119 THEN
            exp_f := 0;
        ELSIF x =- 25118 THEN
            exp_f := 0;
        ELSIF x =- 25117 THEN
            exp_f := 0;
        ELSIF x =- 25116 THEN
            exp_f := 0;
        ELSIF x =- 25115 THEN
            exp_f := 0;
        ELSIF x =- 25114 THEN
            exp_f := 0;
        ELSIF x =- 25113 THEN
            exp_f := 0;
        ELSIF x =- 25112 THEN
            exp_f := 0;
        ELSIF x =- 25111 THEN
            exp_f := 0;
        ELSIF x =- 25110 THEN
            exp_f := 0;
        ELSIF x =- 25109 THEN
            exp_f := 0;
        ELSIF x =- 25108 THEN
            exp_f := 0;
        ELSIF x =- 25107 THEN
            exp_f := 0;
        ELSIF x =- 25106 THEN
            exp_f := 0;
        ELSIF x =- 25105 THEN
            exp_f := 0;
        ELSIF x =- 25104 THEN
            exp_f := 0;
        ELSIF x =- 25103 THEN
            exp_f := 0;
        ELSIF x =- 25102 THEN
            exp_f := 0;
        ELSIF x =- 25101 THEN
            exp_f := 0;
        ELSIF x =- 25100 THEN
            exp_f := 0;
        ELSIF x =- 25099 THEN
            exp_f := 0;
        ELSIF x =- 25098 THEN
            exp_f := 0;
        ELSIF x =- 25097 THEN
            exp_f := 0;
        ELSIF x =- 25096 THEN
            exp_f := 0;
        ELSIF x =- 25095 THEN
            exp_f := 0;
        ELSIF x =- 25094 THEN
            exp_f := 0;
        ELSIF x =- 25093 THEN
            exp_f := 0;
        ELSIF x =- 25092 THEN
            exp_f := 0;
        ELSIF x =- 25091 THEN
            exp_f := 0;
        ELSIF x =- 25090 THEN
            exp_f := 0;
        ELSIF x =- 25089 THEN
            exp_f := 0;
        ELSIF x =- 25088 THEN
            exp_f := 0;
        ELSIF x =- 25087 THEN
            exp_f := 0;
        ELSIF x =- 25086 THEN
            exp_f := 0;
        ELSIF x =- 25085 THEN
            exp_f := 0;
        ELSIF x =- 25084 THEN
            exp_f := 0;
        ELSIF x =- 25083 THEN
            exp_f := 0;
        ELSIF x =- 25082 THEN
            exp_f := 0;
        ELSIF x =- 25081 THEN
            exp_f := 0;
        ELSIF x =- 25080 THEN
            exp_f := 0;
        ELSIF x =- 25079 THEN
            exp_f := 0;
        ELSIF x =- 25078 THEN
            exp_f := 0;
        ELSIF x =- 25077 THEN
            exp_f := 0;
        ELSIF x =- 25076 THEN
            exp_f := 0;
        ELSIF x =- 25075 THEN
            exp_f := 0;
        ELSIF x =- 25074 THEN
            exp_f := 0;
        ELSIF x =- 25073 THEN
            exp_f := 0;
        ELSIF x =- 25072 THEN
            exp_f := 0;
        ELSIF x =- 25071 THEN
            exp_f := 0;
        ELSIF x =- 25070 THEN
            exp_f := 0;
        ELSIF x =- 25069 THEN
            exp_f := 0;
        ELSIF x =- 25068 THEN
            exp_f := 0;
        ELSIF x =- 25067 THEN
            exp_f := 0;
        ELSIF x =- 25066 THEN
            exp_f := 0;
        ELSIF x =- 25065 THEN
            exp_f := 0;
        ELSIF x =- 25064 THEN
            exp_f := 0;
        ELSIF x =- 25063 THEN
            exp_f := 0;
        ELSIF x =- 25062 THEN
            exp_f := 0;
        ELSIF x =- 25061 THEN
            exp_f := 0;
        ELSIF x =- 25060 THEN
            exp_f := 0;
        ELSIF x =- 25059 THEN
            exp_f := 0;
        ELSIF x =- 25058 THEN
            exp_f := 0;
        ELSIF x =- 25057 THEN
            exp_f := 0;
        ELSIF x =- 25056 THEN
            exp_f := 0;
        ELSIF x =- 25055 THEN
            exp_f := 0;
        ELSIF x =- 25054 THEN
            exp_f := 0;
        ELSIF x =- 25053 THEN
            exp_f := 0;
        ELSIF x =- 25052 THEN
            exp_f := 0;
        ELSIF x =- 25051 THEN
            exp_f := 0;
        ELSIF x =- 25050 THEN
            exp_f := 0;
        ELSIF x =- 25049 THEN
            exp_f := 0;
        ELSIF x =- 25048 THEN
            exp_f := 0;
        ELSIF x =- 25047 THEN
            exp_f := 0;
        ELSIF x =- 25046 THEN
            exp_f := 0;
        ELSIF x =- 25045 THEN
            exp_f := 0;
        ELSIF x =- 25044 THEN
            exp_f := 0;
        ELSIF x =- 25043 THEN
            exp_f := 0;
        ELSIF x =- 25042 THEN
            exp_f := 0;
        ELSIF x =- 25041 THEN
            exp_f := 0;
        ELSIF x =- 25040 THEN
            exp_f := 0;
        ELSIF x =- 25039 THEN
            exp_f := 0;
        ELSIF x =- 25038 THEN
            exp_f := 0;
        ELSIF x =- 25037 THEN
            exp_f := 0;
        ELSIF x =- 25036 THEN
            exp_f := 0;
        ELSIF x =- 25035 THEN
            exp_f := 0;
        ELSIF x =- 25034 THEN
            exp_f := 0;
        ELSIF x =- 25033 THEN
            exp_f := 0;
        ELSIF x =- 25032 THEN
            exp_f := 0;
        ELSIF x =- 25031 THEN
            exp_f := 0;
        ELSIF x =- 25030 THEN
            exp_f := 0;
        ELSIF x =- 25029 THEN
            exp_f := 0;
        ELSIF x =- 25028 THEN
            exp_f := 0;
        ELSIF x =- 25027 THEN
            exp_f := 0;
        ELSIF x =- 25026 THEN
            exp_f := 0;
        ELSIF x =- 25025 THEN
            exp_f := 0;
        ELSIF x =- 25024 THEN
            exp_f := 0;
        ELSIF x =- 25023 THEN
            exp_f := 0;
        ELSIF x =- 25022 THEN
            exp_f := 0;
        ELSIF x =- 25021 THEN
            exp_f := 0;
        ELSIF x =- 25020 THEN
            exp_f := 0;
        ELSIF x =- 25019 THEN
            exp_f := 0;
        ELSIF x =- 25018 THEN
            exp_f := 0;
        ELSIF x =- 25017 THEN
            exp_f := 0;
        ELSIF x =- 25016 THEN
            exp_f := 0;
        ELSIF x =- 25015 THEN
            exp_f := 0;
        ELSIF x =- 25014 THEN
            exp_f := 0;
        ELSIF x =- 25013 THEN
            exp_f := 0;
        ELSIF x =- 25012 THEN
            exp_f := 0;
        ELSIF x =- 25011 THEN
            exp_f := 0;
        ELSIF x =- 25010 THEN
            exp_f := 0;
        ELSIF x =- 25009 THEN
            exp_f := 0;
        ELSIF x =- 25008 THEN
            exp_f := 0;
        ELSIF x =- 25007 THEN
            exp_f := 0;
        ELSIF x =- 25006 THEN
            exp_f := 0;
        ELSIF x =- 25005 THEN
            exp_f := 0;
        ELSIF x =- 25004 THEN
            exp_f := 0;
        ELSIF x =- 25003 THEN
            exp_f := 0;
        ELSIF x =- 25002 THEN
            exp_f := 0;
        ELSIF x =- 25001 THEN
            exp_f := 0;
        ELSIF x =- 25000 THEN
            exp_f := 0;
        ELSIF x =- 24999 THEN
            exp_f := 0;
        ELSIF x =- 24998 THEN
            exp_f := 0;
        ELSIF x =- 24997 THEN
            exp_f := 0;
        ELSIF x =- 24996 THEN
            exp_f := 0;
        ELSIF x =- 24995 THEN
            exp_f := 0;
        ELSIF x =- 24994 THEN
            exp_f := 0;
        ELSIF x =- 24993 THEN
            exp_f := 0;
        ELSIF x =- 24992 THEN
            exp_f := 0;
        ELSIF x =- 24991 THEN
            exp_f := 0;
        ELSIF x =- 24990 THEN
            exp_f := 0;
        ELSIF x =- 24989 THEN
            exp_f := 0;
        ELSIF x =- 24988 THEN
            exp_f := 0;
        ELSIF x =- 24987 THEN
            exp_f := 0;
        ELSIF x =- 24986 THEN
            exp_f := 0;
        ELSIF x =- 24985 THEN
            exp_f := 0;
        ELSIF x =- 24984 THEN
            exp_f := 0;
        ELSIF x =- 24983 THEN
            exp_f := 0;
        ELSIF x =- 24982 THEN
            exp_f := 0;
        ELSIF x =- 24981 THEN
            exp_f := 0;
        ELSIF x =- 24980 THEN
            exp_f := 0;
        ELSIF x =- 24979 THEN
            exp_f := 0;
        ELSIF x =- 24978 THEN
            exp_f := 0;
        ELSIF x =- 24977 THEN
            exp_f := 0;
        ELSIF x =- 24976 THEN
            exp_f := 0;
        ELSIF x =- 24975 THEN
            exp_f := 0;
        ELSIF x =- 24974 THEN
            exp_f := 0;
        ELSIF x =- 24973 THEN
            exp_f := 0;
        ELSIF x =- 24972 THEN
            exp_f := 0;
        ELSIF x =- 24971 THEN
            exp_f := 0;
        ELSIF x =- 24970 THEN
            exp_f := 0;
        ELSIF x =- 24969 THEN
            exp_f := 0;
        ELSIF x =- 24968 THEN
            exp_f := 0;
        ELSIF x =- 24967 THEN
            exp_f := 0;
        ELSIF x =- 24966 THEN
            exp_f := 0;
        ELSIF x =- 24965 THEN
            exp_f := 0;
        ELSIF x =- 24964 THEN
            exp_f := 0;
        ELSIF x =- 24963 THEN
            exp_f := 0;
        ELSIF x =- 24962 THEN
            exp_f := 0;
        ELSIF x =- 24961 THEN
            exp_f := 0;
        ELSIF x =- 24960 THEN
            exp_f := 0;
        ELSIF x =- 24959 THEN
            exp_f := 0;
        ELSIF x =- 24958 THEN
            exp_f := 0;
        ELSIF x =- 24957 THEN
            exp_f := 0;
        ELSIF x =- 24956 THEN
            exp_f := 0;
        ELSIF x =- 24955 THEN
            exp_f := 0;
        ELSIF x =- 24954 THEN
            exp_f := 0;
        ELSIF x =- 24953 THEN
            exp_f := 0;
        ELSIF x =- 24952 THEN
            exp_f := 0;
        ELSIF x =- 24951 THEN
            exp_f := 0;
        ELSIF x =- 24950 THEN
            exp_f := 0;
        ELSIF x =- 24949 THEN
            exp_f := 0;
        ELSIF x =- 24948 THEN
            exp_f := 0;
        ELSIF x =- 24947 THEN
            exp_f := 0;
        ELSIF x =- 24946 THEN
            exp_f := 0;
        ELSIF x =- 24945 THEN
            exp_f := 0;
        ELSIF x =- 24944 THEN
            exp_f := 0;
        ELSIF x =- 24943 THEN
            exp_f := 0;
        ELSIF x =- 24942 THEN
            exp_f := 0;
        ELSIF x =- 24941 THEN
            exp_f := 0;
        ELSIF x =- 24940 THEN
            exp_f := 0;
        ELSIF x =- 24939 THEN
            exp_f := 0;
        ELSIF x =- 24938 THEN
            exp_f := 0;
        ELSIF x =- 24937 THEN
            exp_f := 0;
        ELSIF x =- 24936 THEN
            exp_f := 0;
        ELSIF x =- 24935 THEN
            exp_f := 0;
        ELSIF x =- 24934 THEN
            exp_f := 0;
        ELSIF x =- 24933 THEN
            exp_f := 0;
        ELSIF x =- 24932 THEN
            exp_f := 0;
        ELSIF x =- 24931 THEN
            exp_f := 0;
        ELSIF x =- 24930 THEN
            exp_f := 0;
        ELSIF x =- 24929 THEN
            exp_f := 0;
        ELSIF x =- 24928 THEN
            exp_f := 0;
        ELSIF x =- 24927 THEN
            exp_f := 0;
        ELSIF x =- 24926 THEN
            exp_f := 0;
        ELSIF x =- 24925 THEN
            exp_f := 0;
        ELSIF x =- 24924 THEN
            exp_f := 0;
        ELSIF x =- 24923 THEN
            exp_f := 0;
        ELSIF x =- 24922 THEN
            exp_f := 0;
        ELSIF x =- 24921 THEN
            exp_f := 0;
        ELSIF x =- 24920 THEN
            exp_f := 0;
        ELSIF x =- 24919 THEN
            exp_f := 0;
        ELSIF x =- 24918 THEN
            exp_f := 0;
        ELSIF x =- 24917 THEN
            exp_f := 0;
        ELSIF x =- 24916 THEN
            exp_f := 0;
        ELSIF x =- 24915 THEN
            exp_f := 0;
        ELSIF x =- 24914 THEN
            exp_f := 0;
        ELSIF x =- 24913 THEN
            exp_f := 0;
        ELSIF x =- 24912 THEN
            exp_f := 0;
        ELSIF x =- 24911 THEN
            exp_f := 0;
        ELSIF x =- 24910 THEN
            exp_f := 0;
        ELSIF x =- 24909 THEN
            exp_f := 0;
        ELSIF x =- 24908 THEN
            exp_f := 0;
        ELSIF x =- 24907 THEN
            exp_f := 0;
        ELSIF x =- 24906 THEN
            exp_f := 0;
        ELSIF x =- 24905 THEN
            exp_f := 0;
        ELSIF x =- 24904 THEN
            exp_f := 0;
        ELSIF x =- 24903 THEN
            exp_f := 0;
        ELSIF x =- 24902 THEN
            exp_f := 0;
        ELSIF x =- 24901 THEN
            exp_f := 0;
        ELSIF x =- 24900 THEN
            exp_f := 0;
        ELSIF x =- 24899 THEN
            exp_f := 0;
        ELSIF x =- 24898 THEN
            exp_f := 0;
        ELSIF x =- 24897 THEN
            exp_f := 0;
        ELSIF x =- 24896 THEN
            exp_f := 0;
        ELSIF x =- 24895 THEN
            exp_f := 0;
        ELSIF x =- 24894 THEN
            exp_f := 0;
        ELSIF x =- 24893 THEN
            exp_f := 0;
        ELSIF x =- 24892 THEN
            exp_f := 0;
        ELSIF x =- 24891 THEN
            exp_f := 0;
        ELSIF x =- 24890 THEN
            exp_f := 0;
        ELSIF x =- 24889 THEN
            exp_f := 0;
        ELSIF x =- 24888 THEN
            exp_f := 0;
        ELSIF x =- 24887 THEN
            exp_f := 0;
        ELSIF x =- 24886 THEN
            exp_f := 0;
        ELSIF x =- 24885 THEN
            exp_f := 0;
        ELSIF x =- 24884 THEN
            exp_f := 0;
        ELSIF x =- 24883 THEN
            exp_f := 0;
        ELSIF x =- 24882 THEN
            exp_f := 0;
        ELSIF x =- 24881 THEN
            exp_f := 0;
        ELSIF x =- 24880 THEN
            exp_f := 0;
        ELSIF x =- 24879 THEN
            exp_f := 0;
        ELSIF x =- 24878 THEN
            exp_f := 0;
        ELSIF x =- 24877 THEN
            exp_f := 0;
        ELSIF x =- 24876 THEN
            exp_f := 0;
        ELSIF x =- 24875 THEN
            exp_f := 0;
        ELSIF x =- 24874 THEN
            exp_f := 0;
        ELSIF x =- 24873 THEN
            exp_f := 0;
        ELSIF x =- 24872 THEN
            exp_f := 0;
        ELSIF x =- 24871 THEN
            exp_f := 0;
        ELSIF x =- 24870 THEN
            exp_f := 0;
        ELSIF x =- 24869 THEN
            exp_f := 0;
        ELSIF x =- 24868 THEN
            exp_f := 0;
        ELSIF x =- 24867 THEN
            exp_f := 0;
        ELSIF x =- 24866 THEN
            exp_f := 0;
        ELSIF x =- 24865 THEN
            exp_f := 0;
        ELSIF x =- 24864 THEN
            exp_f := 0;
        ELSIF x =- 24863 THEN
            exp_f := 0;
        ELSIF x =- 24862 THEN
            exp_f := 0;
        ELSIF x =- 24861 THEN
            exp_f := 0;
        ELSIF x =- 24860 THEN
            exp_f := 0;
        ELSIF x =- 24859 THEN
            exp_f := 0;
        ELSIF x =- 24858 THEN
            exp_f := 0;
        ELSIF x =- 24857 THEN
            exp_f := 0;
        ELSIF x =- 24856 THEN
            exp_f := 0;
        ELSIF x =- 24855 THEN
            exp_f := 0;
        ELSIF x =- 24854 THEN
            exp_f := 0;
        ELSIF x =- 24853 THEN
            exp_f := 0;
        ELSIF x =- 24852 THEN
            exp_f := 0;
        ELSIF x =- 24851 THEN
            exp_f := 0;
        ELSIF x =- 24850 THEN
            exp_f := 0;
        ELSIF x =- 24849 THEN
            exp_f := 0;
        ELSIF x =- 24848 THEN
            exp_f := 0;
        ELSIF x =- 24847 THEN
            exp_f := 0;
        ELSIF x =- 24846 THEN
            exp_f := 0;
        ELSIF x =- 24845 THEN
            exp_f := 0;
        ELSIF x =- 24844 THEN
            exp_f := 0;
        ELSIF x =- 24843 THEN
            exp_f := 0;
        ELSIF x =- 24842 THEN
            exp_f := 0;
        ELSIF x =- 24841 THEN
            exp_f := 0;
        ELSIF x =- 24840 THEN
            exp_f := 0;
        ELSIF x =- 24839 THEN
            exp_f := 0;
        ELSIF x =- 24838 THEN
            exp_f := 0;
        ELSIF x =- 24837 THEN
            exp_f := 0;
        ELSIF x =- 24836 THEN
            exp_f := 0;
        ELSIF x =- 24835 THEN
            exp_f := 0;
        ELSIF x =- 24834 THEN
            exp_f := 0;
        ELSIF x =- 24833 THEN
            exp_f := 0;
        ELSIF x =- 24832 THEN
            exp_f := 0;
        ELSIF x =- 24831 THEN
            exp_f := 0;
        ELSIF x =- 24830 THEN
            exp_f := 0;
        ELSIF x =- 24829 THEN
            exp_f := 0;
        ELSIF x =- 24828 THEN
            exp_f := 0;
        ELSIF x =- 24827 THEN
            exp_f := 0;
        ELSIF x =- 24826 THEN
            exp_f := 0;
        ELSIF x =- 24825 THEN
            exp_f := 0;
        ELSIF x =- 24824 THEN
            exp_f := 0;
        ELSIF x =- 24823 THEN
            exp_f := 0;
        ELSIF x =- 24822 THEN
            exp_f := 0;
        ELSIF x =- 24821 THEN
            exp_f := 0;
        ELSIF x =- 24820 THEN
            exp_f := 0;
        ELSIF x =- 24819 THEN
            exp_f := 0;
        ELSIF x =- 24818 THEN
            exp_f := 0;
        ELSIF x =- 24817 THEN
            exp_f := 0;
        ELSIF x =- 24816 THEN
            exp_f := 0;
        ELSIF x =- 24815 THEN
            exp_f := 0;
        ELSIF x =- 24814 THEN
            exp_f := 0;
        ELSIF x =- 24813 THEN
            exp_f := 0;
        ELSIF x =- 24812 THEN
            exp_f := 0;
        ELSIF x =- 24811 THEN
            exp_f := 0;
        ELSIF x =- 24810 THEN
            exp_f := 0;
        ELSIF x =- 24809 THEN
            exp_f := 0;
        ELSIF x =- 24808 THEN
            exp_f := 0;
        ELSIF x =- 24807 THEN
            exp_f := 0;
        ELSIF x =- 24806 THEN
            exp_f := 0;
        ELSIF x =- 24805 THEN
            exp_f := 0;
        ELSIF x =- 24804 THEN
            exp_f := 0;
        ELSIF x =- 24803 THEN
            exp_f := 0;
        ELSIF x =- 24802 THEN
            exp_f := 0;
        ELSIF x =- 24801 THEN
            exp_f := 0;
        ELSIF x =- 24800 THEN
            exp_f := 0;
        ELSIF x =- 24799 THEN
            exp_f := 0;
        ELSIF x =- 24798 THEN
            exp_f := 0;
        ELSIF x =- 24797 THEN
            exp_f := 0;
        ELSIF x =- 24796 THEN
            exp_f := 0;
        ELSIF x =- 24795 THEN
            exp_f := 0;
        ELSIF x =- 24794 THEN
            exp_f := 0;
        ELSIF x =- 24793 THEN
            exp_f := 0;
        ELSIF x =- 24792 THEN
            exp_f := 0;
        ELSIF x =- 24791 THEN
            exp_f := 0;
        ELSIF x =- 24790 THEN
            exp_f := 0;
        ELSIF x =- 24789 THEN
            exp_f := 0;
        ELSIF x =- 24788 THEN
            exp_f := 0;
        ELSIF x =- 24787 THEN
            exp_f := 0;
        ELSIF x =- 24786 THEN
            exp_f := 0;
        ELSIF x =- 24785 THEN
            exp_f := 0;
        ELSIF x =- 24784 THEN
            exp_f := 0;
        ELSIF x =- 24783 THEN
            exp_f := 0;
        ELSIF x =- 24782 THEN
            exp_f := 0;
        ELSIF x =- 24781 THEN
            exp_f := 0;
        ELSIF x =- 24780 THEN
            exp_f := 0;
        ELSIF x =- 24779 THEN
            exp_f := 0;
        ELSIF x =- 24778 THEN
            exp_f := 0;
        ELSIF x =- 24777 THEN
            exp_f := 0;
        ELSIF x =- 24776 THEN
            exp_f := 0;
        ELSIF x =- 24775 THEN
            exp_f := 0;
        ELSIF x =- 24774 THEN
            exp_f := 0;
        ELSIF x =- 24773 THEN
            exp_f := 0;
        ELSIF x =- 24772 THEN
            exp_f := 0;
        ELSIF x =- 24771 THEN
            exp_f := 0;
        ELSIF x =- 24770 THEN
            exp_f := 0;
        ELSIF x =- 24769 THEN
            exp_f := 0;
        ELSIF x =- 24768 THEN
            exp_f := 0;
        ELSIF x =- 24767 THEN
            exp_f := 0;
        ELSIF x =- 24766 THEN
            exp_f := 0;
        ELSIF x =- 24765 THEN
            exp_f := 0;
        ELSIF x =- 24764 THEN
            exp_f := 0;
        ELSIF x =- 24763 THEN
            exp_f := 0;
        ELSIF x =- 24762 THEN
            exp_f := 0;
        ELSIF x =- 24761 THEN
            exp_f := 0;
        ELSIF x =- 24760 THEN
            exp_f := 0;
        ELSIF x =- 24759 THEN
            exp_f := 0;
        ELSIF x =- 24758 THEN
            exp_f := 0;
        ELSIF x =- 24757 THEN
            exp_f := 0;
        ELSIF x =- 24756 THEN
            exp_f := 0;
        ELSIF x =- 24755 THEN
            exp_f := 0;
        ELSIF x =- 24754 THEN
            exp_f := 0;
        ELSIF x =- 24753 THEN
            exp_f := 0;
        ELSIF x =- 24752 THEN
            exp_f := 0;
        ELSIF x =- 24751 THEN
            exp_f := 0;
        ELSIF x =- 24750 THEN
            exp_f := 0;
        ELSIF x =- 24749 THEN
            exp_f := 0;
        ELSIF x =- 24748 THEN
            exp_f := 0;
        ELSIF x =- 24747 THEN
            exp_f := 0;
        ELSIF x =- 24746 THEN
            exp_f := 0;
        ELSIF x =- 24745 THEN
            exp_f := 0;
        ELSIF x =- 24744 THEN
            exp_f := 0;
        ELSIF x =- 24743 THEN
            exp_f := 0;
        ELSIF x =- 24742 THEN
            exp_f := 0;
        ELSIF x =- 24741 THEN
            exp_f := 0;
        ELSIF x =- 24740 THEN
            exp_f := 0;
        ELSIF x =- 24739 THEN
            exp_f := 0;
        ELSIF x =- 24738 THEN
            exp_f := 0;
        ELSIF x =- 24737 THEN
            exp_f := 0;
        ELSIF x =- 24736 THEN
            exp_f := 0;
        ELSIF x =- 24735 THEN
            exp_f := 0;
        ELSIF x =- 24734 THEN
            exp_f := 0;
        ELSIF x =- 24733 THEN
            exp_f := 0;
        ELSIF x =- 24732 THEN
            exp_f := 0;
        ELSIF x =- 24731 THEN
            exp_f := 0;
        ELSIF x =- 24730 THEN
            exp_f := 0;
        ELSIF x =- 24729 THEN
            exp_f := 0;
        ELSIF x =- 24728 THEN
            exp_f := 0;
        ELSIF x =- 24727 THEN
            exp_f := 0;
        ELSIF x =- 24726 THEN
            exp_f := 0;
        ELSIF x =- 24725 THEN
            exp_f := 0;
        ELSIF x =- 24724 THEN
            exp_f := 0;
        ELSIF x =- 24723 THEN
            exp_f := 0;
        ELSIF x =- 24722 THEN
            exp_f := 0;
        ELSIF x =- 24721 THEN
            exp_f := 0;
        ELSIF x =- 24720 THEN
            exp_f := 0;
        ELSIF x =- 24719 THEN
            exp_f := 0;
        ELSIF x =- 24718 THEN
            exp_f := 0;
        ELSIF x =- 24717 THEN
            exp_f := 0;
        ELSIF x =- 24716 THEN
            exp_f := 0;
        ELSIF x =- 24715 THEN
            exp_f := 0;
        ELSIF x =- 24714 THEN
            exp_f := 0;
        ELSIF x =- 24713 THEN
            exp_f := 0;
        ELSIF x =- 24712 THEN
            exp_f := 0;
        ELSIF x =- 24711 THEN
            exp_f := 0;
        ELSIF x =- 24710 THEN
            exp_f := 0;
        ELSIF x =- 24709 THEN
            exp_f := 0;
        ELSIF x =- 24708 THEN
            exp_f := 0;
        ELSIF x =- 24707 THEN
            exp_f := 0;
        ELSIF x =- 24706 THEN
            exp_f := 0;
        ELSIF x =- 24705 THEN
            exp_f := 0;
        ELSIF x =- 24704 THEN
            exp_f := 0;
        ELSIF x =- 24703 THEN
            exp_f := 0;
        ELSIF x =- 24702 THEN
            exp_f := 0;
        ELSIF x =- 24701 THEN
            exp_f := 0;
        ELSIF x =- 24700 THEN
            exp_f := 0;
        ELSIF x =- 24699 THEN
            exp_f := 0;
        ELSIF x =- 24698 THEN
            exp_f := 0;
        ELSIF x =- 24697 THEN
            exp_f := 0;
        ELSIF x =- 24696 THEN
            exp_f := 0;
        ELSIF x =- 24695 THEN
            exp_f := 0;
        ELSIF x =- 24694 THEN
            exp_f := 0;
        ELSIF x =- 24693 THEN
            exp_f := 0;
        ELSIF x =- 24692 THEN
            exp_f := 0;
        ELSIF x =- 24691 THEN
            exp_f := 0;
        ELSIF x =- 24690 THEN
            exp_f := 0;
        ELSIF x =- 24689 THEN
            exp_f := 0;
        ELSIF x =- 24688 THEN
            exp_f := 0;
        ELSIF x =- 24687 THEN
            exp_f := 0;
        ELSIF x =- 24686 THEN
            exp_f := 0;
        ELSIF x =- 24685 THEN
            exp_f := 0;
        ELSIF x =- 24684 THEN
            exp_f := 0;
        ELSIF x =- 24683 THEN
            exp_f := 0;
        ELSIF x =- 24682 THEN
            exp_f := 0;
        ELSIF x =- 24681 THEN
            exp_f := 0;
        ELSIF x =- 24680 THEN
            exp_f := 0;
        ELSIF x =- 24679 THEN
            exp_f := 0;
        ELSIF x =- 24678 THEN
            exp_f := 0;
        ELSIF x =- 24677 THEN
            exp_f := 0;
        ELSIF x =- 24676 THEN
            exp_f := 0;
        ELSIF x =- 24675 THEN
            exp_f := 0;
        ELSIF x =- 24674 THEN
            exp_f := 0;
        ELSIF x =- 24673 THEN
            exp_f := 0;
        ELSIF x =- 24672 THEN
            exp_f := 0;
        ELSIF x =- 24671 THEN
            exp_f := 0;
        ELSIF x =- 24670 THEN
            exp_f := 0;
        ELSIF x =- 24669 THEN
            exp_f := 0;
        ELSIF x =- 24668 THEN
            exp_f := 0;
        ELSIF x =- 24667 THEN
            exp_f := 0;
        ELSIF x =- 24666 THEN
            exp_f := 0;
        ELSIF x =- 24665 THEN
            exp_f := 0;
        ELSIF x =- 24664 THEN
            exp_f := 0;
        ELSIF x =- 24663 THEN
            exp_f := 0;
        ELSIF x =- 24662 THEN
            exp_f := 0;
        ELSIF x =- 24661 THEN
            exp_f := 0;
        ELSIF x =- 24660 THEN
            exp_f := 0;
        ELSIF x =- 24659 THEN
            exp_f := 0;
        ELSIF x =- 24658 THEN
            exp_f := 0;
        ELSIF x =- 24657 THEN
            exp_f := 0;
        ELSIF x =- 24656 THEN
            exp_f := 0;
        ELSIF x =- 24655 THEN
            exp_f := 0;
        ELSIF x =- 24654 THEN
            exp_f := 0;
        ELSIF x =- 24653 THEN
            exp_f := 0;
        ELSIF x =- 24652 THEN
            exp_f := 0;
        ELSIF x =- 24651 THEN
            exp_f := 0;
        ELSIF x =- 24650 THEN
            exp_f := 0;
        ELSIF x =- 24649 THEN
            exp_f := 0;
        ELSIF x =- 24648 THEN
            exp_f := 0;
        ELSIF x =- 24647 THEN
            exp_f := 0;
        ELSIF x =- 24646 THEN
            exp_f := 0;
        ELSIF x =- 24645 THEN
            exp_f := 0;
        ELSIF x =- 24644 THEN
            exp_f := 0;
        ELSIF x =- 24643 THEN
            exp_f := 0;
        ELSIF x =- 24642 THEN
            exp_f := 0;
        ELSIF x =- 24641 THEN
            exp_f := 0;
        ELSIF x =- 24640 THEN
            exp_f := 0;
        ELSIF x =- 24639 THEN
            exp_f := 0;
        ELSIF x =- 24638 THEN
            exp_f := 0;
        ELSIF x =- 24637 THEN
            exp_f := 0;
        ELSIF x =- 24636 THEN
            exp_f := 0;
        ELSIF x =- 24635 THEN
            exp_f := 0;
        ELSIF x =- 24634 THEN
            exp_f := 0;
        ELSIF x =- 24633 THEN
            exp_f := 0;
        ELSIF x =- 24632 THEN
            exp_f := 0;
        ELSIF x =- 24631 THEN
            exp_f := 0;
        ELSIF x =- 24630 THEN
            exp_f := 0;
        ELSIF x =- 24629 THEN
            exp_f := 0;
        ELSIF x =- 24628 THEN
            exp_f := 0;
        ELSIF x =- 24627 THEN
            exp_f := 0;
        ELSIF x =- 24626 THEN
            exp_f := 0;
        ELSIF x =- 24625 THEN
            exp_f := 0;
        ELSIF x =- 24624 THEN
            exp_f := 0;
        ELSIF x =- 24623 THEN
            exp_f := 0;
        ELSIF x =- 24622 THEN
            exp_f := 0;
        ELSIF x =- 24621 THEN
            exp_f := 0;
        ELSIF x =- 24620 THEN
            exp_f := 0;
        ELSIF x =- 24619 THEN
            exp_f := 0;
        ELSIF x =- 24618 THEN
            exp_f := 0;
        ELSIF x =- 24617 THEN
            exp_f := 0;
        ELSIF x =- 24616 THEN
            exp_f := 0;
        ELSIF x =- 24615 THEN
            exp_f := 0;
        ELSIF x =- 24614 THEN
            exp_f := 0;
        ELSIF x =- 24613 THEN
            exp_f := 0;
        ELSIF x =- 24612 THEN
            exp_f := 0;
        ELSIF x =- 24611 THEN
            exp_f := 0;
        ELSIF x =- 24610 THEN
            exp_f := 0;
        ELSIF x =- 24609 THEN
            exp_f := 0;
        ELSIF x =- 24608 THEN
            exp_f := 0;
        ELSIF x =- 24607 THEN
            exp_f := 0;
        ELSIF x =- 24606 THEN
            exp_f := 0;
        ELSIF x =- 24605 THEN
            exp_f := 0;
        ELSIF x =- 24604 THEN
            exp_f := 0;
        ELSIF x =- 24603 THEN
            exp_f := 0;
        ELSIF x =- 24602 THEN
            exp_f := 0;
        ELSIF x =- 24601 THEN
            exp_f := 0;
        ELSIF x =- 24600 THEN
            exp_f := 0;
        ELSIF x =- 24599 THEN
            exp_f := 0;
        ELSIF x =- 24598 THEN
            exp_f := 0;
        ELSIF x =- 24597 THEN
            exp_f := 0;
        ELSIF x =- 24596 THEN
            exp_f := 0;
        ELSIF x =- 24595 THEN
            exp_f := 0;
        ELSIF x =- 24594 THEN
            exp_f := 0;
        ELSIF x =- 24593 THEN
            exp_f := 0;
        ELSIF x =- 24592 THEN
            exp_f := 0;
        ELSIF x =- 24591 THEN
            exp_f := 0;
        ELSIF x =- 24590 THEN
            exp_f := 0;
        ELSIF x =- 24589 THEN
            exp_f := 0;
        ELSIF x =- 24588 THEN
            exp_f := 0;
        ELSIF x =- 24587 THEN
            exp_f := 0;
        ELSIF x =- 24586 THEN
            exp_f := 0;
        ELSIF x =- 24585 THEN
            exp_f := 0;
        ELSIF x =- 24584 THEN
            exp_f := 0;
        ELSIF x =- 24583 THEN
            exp_f := 0;
        ELSIF x =- 24582 THEN
            exp_f := 0;
        ELSIF x =- 24581 THEN
            exp_f := 0;
        ELSIF x =- 24580 THEN
            exp_f := 0;
        ELSIF x =- 24579 THEN
            exp_f := 0;
        ELSIF x =- 24578 THEN
            exp_f := 0;
        ELSIF x =- 24577 THEN
            exp_f := 0;
        ELSIF x =- 24576 THEN
            exp_f := 0;
        ELSIF x =- 24575 THEN
            exp_f := 0;
        ELSIF x =- 24574 THEN
            exp_f := 0;
        ELSIF x =- 24573 THEN
            exp_f := 0;
        ELSIF x =- 24572 THEN
            exp_f := 0;
        ELSIF x =- 24571 THEN
            exp_f := 0;
        ELSIF x =- 24570 THEN
            exp_f := 0;
        ELSIF x =- 24569 THEN
            exp_f := 0;
        ELSIF x =- 24568 THEN
            exp_f := 0;
        ELSIF x =- 24567 THEN
            exp_f := 0;
        ELSIF x =- 24566 THEN
            exp_f := 0;
        ELSIF x =- 24565 THEN
            exp_f := 0;
        ELSIF x =- 24564 THEN
            exp_f := 0;
        ELSIF x =- 24563 THEN
            exp_f := 0;
        ELSIF x =- 24562 THEN
            exp_f := 0;
        ELSIF x =- 24561 THEN
            exp_f := 0;
        ELSIF x =- 24560 THEN
            exp_f := 0;
        ELSIF x =- 24559 THEN
            exp_f := 0;
        ELSIF x =- 24558 THEN
            exp_f := 0;
        ELSIF x =- 24557 THEN
            exp_f := 0;
        ELSIF x =- 24556 THEN
            exp_f := 0;
        ELSIF x =- 24555 THEN
            exp_f := 0;
        ELSIF x =- 24554 THEN
            exp_f := 0;
        ELSIF x =- 24553 THEN
            exp_f := 0;
        ELSIF x =- 24552 THEN
            exp_f := 0;
        ELSIF x =- 24551 THEN
            exp_f := 0;
        ELSIF x =- 24550 THEN
            exp_f := 0;
        ELSIF x =- 24549 THEN
            exp_f := 0;
        ELSIF x =- 24548 THEN
            exp_f := 0;
        ELSIF x =- 24547 THEN
            exp_f := 0;
        ELSIF x =- 24546 THEN
            exp_f := 0;
        ELSIF x =- 24545 THEN
            exp_f := 0;
        ELSIF x =- 24544 THEN
            exp_f := 0;
        ELSIF x =- 24543 THEN
            exp_f := 0;
        ELSIF x =- 24542 THEN
            exp_f := 0;
        ELSIF x =- 24541 THEN
            exp_f := 0;
        ELSIF x =- 24540 THEN
            exp_f := 0;
        ELSIF x =- 24539 THEN
            exp_f := 0;
        ELSIF x =- 24538 THEN
            exp_f := 0;
        ELSIF x =- 24537 THEN
            exp_f := 0;
        ELSIF x =- 24536 THEN
            exp_f := 0;
        ELSIF x =- 24535 THEN
            exp_f := 0;
        ELSIF x =- 24534 THEN
            exp_f := 0;
        ELSIF x =- 24533 THEN
            exp_f := 0;
        ELSIF x =- 24532 THEN
            exp_f := 0;
        ELSIF x =- 24531 THEN
            exp_f := 0;
        ELSIF x =- 24530 THEN
            exp_f := 0;
        ELSIF x =- 24529 THEN
            exp_f := 0;
        ELSIF x =- 24528 THEN
            exp_f := 0;
        ELSIF x =- 24527 THEN
            exp_f := 0;
        ELSIF x =- 24526 THEN
            exp_f := 0;
        ELSIF x =- 24525 THEN
            exp_f := 0;
        ELSIF x =- 24524 THEN
            exp_f := 0;
        ELSIF x =- 24523 THEN
            exp_f := 0;
        ELSIF x =- 24522 THEN
            exp_f := 0;
        ELSIF x =- 24521 THEN
            exp_f := 0;
        ELSIF x =- 24520 THEN
            exp_f := 0;
        ELSIF x =- 24519 THEN
            exp_f := 0;
        ELSIF x =- 24518 THEN
            exp_f := 0;
        ELSIF x =- 24517 THEN
            exp_f := 0;
        ELSIF x =- 24516 THEN
            exp_f := 0;
        ELSIF x =- 24515 THEN
            exp_f := 0;
        ELSIF x =- 24514 THEN
            exp_f := 0;
        ELSIF x =- 24513 THEN
            exp_f := 0;
        ELSIF x =- 24512 THEN
            exp_f := 0;
        ELSIF x =- 24511 THEN
            exp_f := 0;
        ELSIF x =- 24510 THEN
            exp_f := 0;
        ELSIF x =- 24509 THEN
            exp_f := 0;
        ELSIF x =- 24508 THEN
            exp_f := 0;
        ELSIF x =- 24507 THEN
            exp_f := 0;
        ELSIF x =- 24506 THEN
            exp_f := 0;
        ELSIF x =- 24505 THEN
            exp_f := 0;
        ELSIF x =- 24504 THEN
            exp_f := 0;
        ELSIF x =- 24503 THEN
            exp_f := 0;
        ELSIF x =- 24502 THEN
            exp_f := 0;
        ELSIF x =- 24501 THEN
            exp_f := 0;
        ELSIF x =- 24500 THEN
            exp_f := 0;
        ELSIF x =- 24499 THEN
            exp_f := 0;
        ELSIF x =- 24498 THEN
            exp_f := 0;
        ELSIF x =- 24497 THEN
            exp_f := 0;
        ELSIF x =- 24496 THEN
            exp_f := 0;
        ELSIF x =- 24495 THEN
            exp_f := 0;
        ELSIF x =- 24494 THEN
            exp_f := 0;
        ELSIF x =- 24493 THEN
            exp_f := 0;
        ELSIF x =- 24492 THEN
            exp_f := 0;
        ELSIF x =- 24491 THEN
            exp_f := 0;
        ELSIF x =- 24490 THEN
            exp_f := 0;
        ELSIF x =- 24489 THEN
            exp_f := 0;
        ELSIF x =- 24488 THEN
            exp_f := 0;
        ELSIF x =- 24487 THEN
            exp_f := 0;
        ELSIF x =- 24486 THEN
            exp_f := 0;
        ELSIF x =- 24485 THEN
            exp_f := 0;
        ELSIF x =- 24484 THEN
            exp_f := 0;
        ELSIF x =- 24483 THEN
            exp_f := 0;
        ELSIF x =- 24482 THEN
            exp_f := 0;
        ELSIF x =- 24481 THEN
            exp_f := 0;
        ELSIF x =- 24480 THEN
            exp_f := 0;
        ELSIF x =- 24479 THEN
            exp_f := 0;
        ELSIF x =- 24478 THEN
            exp_f := 0;
        ELSIF x =- 24477 THEN
            exp_f := 0;
        ELSIF x =- 24476 THEN
            exp_f := 0;
        ELSIF x =- 24475 THEN
            exp_f := 0;
        ELSIF x =- 24474 THEN
            exp_f := 0;
        ELSIF x =- 24473 THEN
            exp_f := 0;
        ELSIF x =- 24472 THEN
            exp_f := 0;
        ELSIF x =- 24471 THEN
            exp_f := 0;
        ELSIF x =- 24470 THEN
            exp_f := 0;
        ELSIF x =- 24469 THEN
            exp_f := 0;
        ELSIF x =- 24468 THEN
            exp_f := 0;
        ELSIF x =- 24467 THEN
            exp_f := 0;
        ELSIF x =- 24466 THEN
            exp_f := 0;
        ELSIF x =- 24465 THEN
            exp_f := 0;
        ELSIF x =- 24464 THEN
            exp_f := 0;
        ELSIF x =- 24463 THEN
            exp_f := 0;
        ELSIF x =- 24462 THEN
            exp_f := 0;
        ELSIF x =- 24461 THEN
            exp_f := 0;
        ELSIF x =- 24460 THEN
            exp_f := 0;
        ELSIF x =- 24459 THEN
            exp_f := 0;
        ELSIF x =- 24458 THEN
            exp_f := 0;
        ELSIF x =- 24457 THEN
            exp_f := 0;
        ELSIF x =- 24456 THEN
            exp_f := 0;
        ELSIF x =- 24455 THEN
            exp_f := 0;
        ELSIF x =- 24454 THEN
            exp_f := 0;
        ELSIF x =- 24453 THEN
            exp_f := 0;
        ELSIF x =- 24452 THEN
            exp_f := 0;
        ELSIF x =- 24451 THEN
            exp_f := 0;
        ELSIF x =- 24450 THEN
            exp_f := 0;
        ELSIF x =- 24449 THEN
            exp_f := 0;
        ELSIF x =- 24448 THEN
            exp_f := 0;
        ELSIF x =- 24447 THEN
            exp_f := 0;
        ELSIF x =- 24446 THEN
            exp_f := 0;
        ELSIF x =- 24445 THEN
            exp_f := 0;
        ELSIF x =- 24444 THEN
            exp_f := 0;
        ELSIF x =- 24443 THEN
            exp_f := 0;
        ELSIF x =- 24442 THEN
            exp_f := 0;
        ELSIF x =- 24441 THEN
            exp_f := 0;
        ELSIF x =- 24440 THEN
            exp_f := 0;
        ELSIF x =- 24439 THEN
            exp_f := 0;
        ELSIF x =- 24438 THEN
            exp_f := 0;
        ELSIF x =- 24437 THEN
            exp_f := 0;
        ELSIF x =- 24436 THEN
            exp_f := 0;
        ELSIF x =- 24435 THEN
            exp_f := 0;
        ELSIF x =- 24434 THEN
            exp_f := 0;
        ELSIF x =- 24433 THEN
            exp_f := 0;
        ELSIF x =- 24432 THEN
            exp_f := 0;
        ELSIF x =- 24431 THEN
            exp_f := 0;
        ELSIF x =- 24430 THEN
            exp_f := 0;
        ELSIF x =- 24429 THEN
            exp_f := 0;
        ELSIF x =- 24428 THEN
            exp_f := 0;
        ELSIF x =- 24427 THEN
            exp_f := 0;
        ELSIF x =- 24426 THEN
            exp_f := 0;
        ELSIF x =- 24425 THEN
            exp_f := 0;
        ELSIF x =- 24424 THEN
            exp_f := 0;
        ELSIF x =- 24423 THEN
            exp_f := 0;
        ELSIF x =- 24422 THEN
            exp_f := 0;
        ELSIF x =- 24421 THEN
            exp_f := 0;
        ELSIF x =- 24420 THEN
            exp_f := 0;
        ELSIF x =- 24419 THEN
            exp_f := 0;
        ELSIF x =- 24418 THEN
            exp_f := 0;
        ELSIF x =- 24417 THEN
            exp_f := 0;
        ELSIF x =- 24416 THEN
            exp_f := 0;
        ELSIF x =- 24415 THEN
            exp_f := 0;
        ELSIF x =- 24414 THEN
            exp_f := 0;
        ELSIF x =- 24413 THEN
            exp_f := 0;
        ELSIF x =- 24412 THEN
            exp_f := 0;
        ELSIF x =- 24411 THEN
            exp_f := 0;
        ELSIF x =- 24410 THEN
            exp_f := 0;
        ELSIF x =- 24409 THEN
            exp_f := 0;
        ELSIF x =- 24408 THEN
            exp_f := 0;
        ELSIF x =- 24407 THEN
            exp_f := 0;
        ELSIF x =- 24406 THEN
            exp_f := 0;
        ELSIF x =- 24405 THEN
            exp_f := 0;
        ELSIF x =- 24404 THEN
            exp_f := 0;
        ELSIF x =- 24403 THEN
            exp_f := 0;
        ELSIF x =- 24402 THEN
            exp_f := 0;
        ELSIF x =- 24401 THEN
            exp_f := 0;
        ELSIF x =- 24400 THEN
            exp_f := 0;
        ELSIF x =- 24399 THEN
            exp_f := 0;
        ELSIF x =- 24398 THEN
            exp_f := 0;
        ELSIF x =- 24397 THEN
            exp_f := 0;
        ELSIF x =- 24396 THEN
            exp_f := 0;
        ELSIF x =- 24395 THEN
            exp_f := 0;
        ELSIF x =- 24394 THEN
            exp_f := 0;
        ELSIF x =- 24393 THEN
            exp_f := 0;
        ELSIF x =- 24392 THEN
            exp_f := 0;
        ELSIF x =- 24391 THEN
            exp_f := 0;
        ELSIF x =- 24390 THEN
            exp_f := 0;
        ELSIF x =- 24389 THEN
            exp_f := 0;
        ELSIF x =- 24388 THEN
            exp_f := 0;
        ELSIF x =- 24387 THEN
            exp_f := 0;
        ELSIF x =- 24386 THEN
            exp_f := 0;
        ELSIF x =- 24385 THEN
            exp_f := 0;
        ELSIF x =- 24384 THEN
            exp_f := 0;
        ELSIF x =- 24383 THEN
            exp_f := 0;
        ELSIF x =- 24382 THEN
            exp_f := 0;
        ELSIF x =- 24381 THEN
            exp_f := 0;
        ELSIF x =- 24380 THEN
            exp_f := 0;
        ELSIF x =- 24379 THEN
            exp_f := 0;
        ELSIF x =- 24378 THEN
            exp_f := 0;
        ELSIF x =- 24377 THEN
            exp_f := 0;
        ELSIF x =- 24376 THEN
            exp_f := 0;
        ELSIF x =- 24375 THEN
            exp_f := 0;
        ELSIF x =- 24374 THEN
            exp_f := 0;
        ELSIF x =- 24373 THEN
            exp_f := 0;
        ELSIF x =- 24372 THEN
            exp_f := 0;
        ELSIF x =- 24371 THEN
            exp_f := 0;
        ELSIF x =- 24370 THEN
            exp_f := 0;
        ELSIF x =- 24369 THEN
            exp_f := 0;
        ELSIF x =- 24368 THEN
            exp_f := 0;
        ELSIF x =- 24367 THEN
            exp_f := 0;
        ELSIF x =- 24366 THEN
            exp_f := 0;
        ELSIF x =- 24365 THEN
            exp_f := 0;
        ELSIF x =- 24364 THEN
            exp_f := 0;
        ELSIF x =- 24363 THEN
            exp_f := 0;
        ELSIF x =- 24362 THEN
            exp_f := 0;
        ELSIF x =- 24361 THEN
            exp_f := 0;
        ELSIF x =- 24360 THEN
            exp_f := 0;
        ELSIF x =- 24359 THEN
            exp_f := 0;
        ELSIF x =- 24358 THEN
            exp_f := 0;
        ELSIF x =- 24357 THEN
            exp_f := 0;
        ELSIF x =- 24356 THEN
            exp_f := 0;
        ELSIF x =- 24355 THEN
            exp_f := 0;
        ELSIF x =- 24354 THEN
            exp_f := 0;
        ELSIF x =- 24353 THEN
            exp_f := 0;
        ELSIF x =- 24352 THEN
            exp_f := 0;
        ELSIF x =- 24351 THEN
            exp_f := 0;
        ELSIF x =- 24350 THEN
            exp_f := 0;
        ELSIF x =- 24349 THEN
            exp_f := 0;
        ELSIF x =- 24348 THEN
            exp_f := 0;
        ELSIF x =- 24347 THEN
            exp_f := 0;
        ELSIF x =- 24346 THEN
            exp_f := 0;
        ELSIF x =- 24345 THEN
            exp_f := 0;
        ELSIF x =- 24344 THEN
            exp_f := 0;
        ELSIF x =- 24343 THEN
            exp_f := 0;
        ELSIF x =- 24342 THEN
            exp_f := 0;
        ELSIF x =- 24341 THEN
            exp_f := 0;
        ELSIF x =- 24340 THEN
            exp_f := 0;
        ELSIF x =- 24339 THEN
            exp_f := 0;
        ELSIF x =- 24338 THEN
            exp_f := 0;
        ELSIF x =- 24337 THEN
            exp_f := 0;
        ELSIF x =- 24336 THEN
            exp_f := 0;
        ELSIF x =- 24335 THEN
            exp_f := 0;
        ELSIF x =- 24334 THEN
            exp_f := 0;
        ELSIF x =- 24333 THEN
            exp_f := 0;
        ELSIF x =- 24332 THEN
            exp_f := 0;
        ELSIF x =- 24331 THEN
            exp_f := 0;
        ELSIF x =- 24330 THEN
            exp_f := 0;
        ELSIF x =- 24329 THEN
            exp_f := 0;
        ELSIF x =- 24328 THEN
            exp_f := 0;
        ELSIF x =- 24327 THEN
            exp_f := 0;
        ELSIF x =- 24326 THEN
            exp_f := 0;
        ELSIF x =- 24325 THEN
            exp_f := 0;
        ELSIF x =- 24324 THEN
            exp_f := 0;
        ELSIF x =- 24323 THEN
            exp_f := 0;
        ELSIF x =- 24322 THEN
            exp_f := 0;
        ELSIF x =- 24321 THEN
            exp_f := 0;
        ELSIF x =- 24320 THEN
            exp_f := 0;
        ELSIF x =- 24319 THEN
            exp_f := 0;
        ELSIF x =- 24318 THEN
            exp_f := 0;
        ELSIF x =- 24317 THEN
            exp_f := 0;
        ELSIF x =- 24316 THEN
            exp_f := 0;
        ELSIF x =- 24315 THEN
            exp_f := 0;
        ELSIF x =- 24314 THEN
            exp_f := 0;
        ELSIF x =- 24313 THEN
            exp_f := 0;
        ELSIF x =- 24312 THEN
            exp_f := 0;
        ELSIF x =- 24311 THEN
            exp_f := 0;
        ELSIF x =- 24310 THEN
            exp_f := 0;
        ELSIF x =- 24309 THEN
            exp_f := 0;
        ELSIF x =- 24308 THEN
            exp_f := 0;
        ELSIF x =- 24307 THEN
            exp_f := 0;
        ELSIF x =- 24306 THEN
            exp_f := 0;
        ELSIF x =- 24305 THEN
            exp_f := 0;
        ELSIF x =- 24304 THEN
            exp_f := 0;
        ELSIF x =- 24303 THEN
            exp_f := 0;
        ELSIF x =- 24302 THEN
            exp_f := 0;
        ELSIF x =- 24301 THEN
            exp_f := 0;
        ELSIF x =- 24300 THEN
            exp_f := 0;
        ELSIF x =- 24299 THEN
            exp_f := 0;
        ELSIF x =- 24298 THEN
            exp_f := 0;
        ELSIF x =- 24297 THEN
            exp_f := 0;
        ELSIF x =- 24296 THEN
            exp_f := 0;
        ELSIF x =- 24295 THEN
            exp_f := 0;
        ELSIF x =- 24294 THEN
            exp_f := 0;
        ELSIF x =- 24293 THEN
            exp_f := 0;
        ELSIF x =- 24292 THEN
            exp_f := 0;
        ELSIF x =- 24291 THEN
            exp_f := 0;
        ELSIF x =- 24290 THEN
            exp_f := 0;
        ELSIF x =- 24289 THEN
            exp_f := 0;
        ELSIF x =- 24288 THEN
            exp_f := 0;
        ELSIF x =- 24287 THEN
            exp_f := 0;
        ELSIF x =- 24286 THEN
            exp_f := 0;
        ELSIF x =- 24285 THEN
            exp_f := 0;
        ELSIF x =- 24284 THEN
            exp_f := 0;
        ELSIF x =- 24283 THEN
            exp_f := 0;
        ELSIF x =- 24282 THEN
            exp_f := 0;
        ELSIF x =- 24281 THEN
            exp_f := 0;
        ELSIF x =- 24280 THEN
            exp_f := 0;
        ELSIF x =- 24279 THEN
            exp_f := 0;
        ELSIF x =- 24278 THEN
            exp_f := 0;
        ELSIF x =- 24277 THEN
            exp_f := 0;
        ELSIF x =- 24276 THEN
            exp_f := 0;
        ELSIF x =- 24275 THEN
            exp_f := 0;
        ELSIF x =- 24274 THEN
            exp_f := 0;
        ELSIF x =- 24273 THEN
            exp_f := 0;
        ELSIF x =- 24272 THEN
            exp_f := 0;
        ELSIF x =- 24271 THEN
            exp_f := 0;
        ELSIF x =- 24270 THEN
            exp_f := 0;
        ELSIF x =- 24269 THEN
            exp_f := 0;
        ELSIF x =- 24268 THEN
            exp_f := 0;
        ELSIF x =- 24267 THEN
            exp_f := 0;
        ELSIF x =- 24266 THEN
            exp_f := 0;
        ELSIF x =- 24265 THEN
            exp_f := 0;
        ELSIF x =- 24264 THEN
            exp_f := 0;
        ELSIF x =- 24263 THEN
            exp_f := 0;
        ELSIF x =- 24262 THEN
            exp_f := 0;
        ELSIF x =- 24261 THEN
            exp_f := 0;
        ELSIF x =- 24260 THEN
            exp_f := 0;
        ELSIF x =- 24259 THEN
            exp_f := 0;
        ELSIF x =- 24258 THEN
            exp_f := 0;
        ELSIF x =- 24257 THEN
            exp_f := 0;
        ELSIF x =- 24256 THEN
            exp_f := 0;
        ELSIF x =- 24255 THEN
            exp_f := 0;
        ELSIF x =- 24254 THEN
            exp_f := 0;
        ELSIF x =- 24253 THEN
            exp_f := 0;
        ELSIF x =- 24252 THEN
            exp_f := 0;
        ELSIF x =- 24251 THEN
            exp_f := 0;
        ELSIF x =- 24250 THEN
            exp_f := 0;
        ELSIF x =- 24249 THEN
            exp_f := 0;
        ELSIF x =- 24248 THEN
            exp_f := 0;
        ELSIF x =- 24247 THEN
            exp_f := 0;
        ELSIF x =- 24246 THEN
            exp_f := 0;
        ELSIF x =- 24245 THEN
            exp_f := 0;
        ELSIF x =- 24244 THEN
            exp_f := 0;
        ELSIF x =- 24243 THEN
            exp_f := 0;
        ELSIF x =- 24242 THEN
            exp_f := 0;
        ELSIF x =- 24241 THEN
            exp_f := 0;
        ELSIF x =- 24240 THEN
            exp_f := 0;
        ELSIF x =- 24239 THEN
            exp_f := 0;
        ELSIF x =- 24238 THEN
            exp_f := 0;
        ELSIF x =- 24237 THEN
            exp_f := 0;
        ELSIF x =- 24236 THEN
            exp_f := 0;
        ELSIF x =- 24235 THEN
            exp_f := 0;
        ELSIF x =- 24234 THEN
            exp_f := 0;
        ELSIF x =- 24233 THEN
            exp_f := 0;
        ELSIF x =- 24232 THEN
            exp_f := 0;
        ELSIF x =- 24231 THEN
            exp_f := 0;
        ELSIF x =- 24230 THEN
            exp_f := 0;
        ELSIF x =- 24229 THEN
            exp_f := 0;
        ELSIF x =- 24228 THEN
            exp_f := 0;
        ELSIF x =- 24227 THEN
            exp_f := 0;
        ELSIF x =- 24226 THEN
            exp_f := 0;
        ELSIF x =- 24225 THEN
            exp_f := 0;
        ELSIF x =- 24224 THEN
            exp_f := 0;
        ELSIF x =- 24223 THEN
            exp_f := 0;
        ELSIF x =- 24222 THEN
            exp_f := 0;
        ELSIF x =- 24221 THEN
            exp_f := 0;
        ELSIF x =- 24220 THEN
            exp_f := 0;
        ELSIF x =- 24219 THEN
            exp_f := 0;
        ELSIF x =- 24218 THEN
            exp_f := 0;
        ELSIF x =- 24217 THEN
            exp_f := 0;
        ELSIF x =- 24216 THEN
            exp_f := 0;
        ELSIF x =- 24215 THEN
            exp_f := 0;
        ELSIF x =- 24214 THEN
            exp_f := 0;
        ELSIF x =- 24213 THEN
            exp_f := 0;
        ELSIF x =- 24212 THEN
            exp_f := 0;
        ELSIF x =- 24211 THEN
            exp_f := 0;
        ELSIF x =- 24210 THEN
            exp_f := 0;
        ELSIF x =- 24209 THEN
            exp_f := 0;
        ELSIF x =- 24208 THEN
            exp_f := 0;
        ELSIF x =- 24207 THEN
            exp_f := 0;
        ELSIF x =- 24206 THEN
            exp_f := 0;
        ELSIF x =- 24205 THEN
            exp_f := 0;
        ELSIF x =- 24204 THEN
            exp_f := 0;
        ELSIF x =- 24203 THEN
            exp_f := 0;
        ELSIF x =- 24202 THEN
            exp_f := 0;
        ELSIF x =- 24201 THEN
            exp_f := 0;
        ELSIF x =- 24200 THEN
            exp_f := 0;
        ELSIF x =- 24199 THEN
            exp_f := 0;
        ELSIF x =- 24198 THEN
            exp_f := 0;
        ELSIF x =- 24197 THEN
            exp_f := 0;
        ELSIF x =- 24196 THEN
            exp_f := 0;
        ELSIF x =- 24195 THEN
            exp_f := 0;
        ELSIF x =- 24194 THEN
            exp_f := 0;
        ELSIF x =- 24193 THEN
            exp_f := 0;
        ELSIF x =- 24192 THEN
            exp_f := 0;
        ELSIF x =- 24191 THEN
            exp_f := 0;
        ELSIF x =- 24190 THEN
            exp_f := 0;
        ELSIF x =- 24189 THEN
            exp_f := 0;
        ELSIF x =- 24188 THEN
            exp_f := 0;
        ELSIF x =- 24187 THEN
            exp_f := 0;
        ELSIF x =- 24186 THEN
            exp_f := 0;
        ELSIF x =- 24185 THEN
            exp_f := 0;
        ELSIF x =- 24184 THEN
            exp_f := 0;
        ELSIF x =- 24183 THEN
            exp_f := 0;
        ELSIF x =- 24182 THEN
            exp_f := 0;
        ELSIF x =- 24181 THEN
            exp_f := 0;
        ELSIF x =- 24180 THEN
            exp_f := 0;
        ELSIF x =- 24179 THEN
            exp_f := 0;
        ELSIF x =- 24178 THEN
            exp_f := 0;
        ELSIF x =- 24177 THEN
            exp_f := 0;
        ELSIF x =- 24176 THEN
            exp_f := 0;
        ELSIF x =- 24175 THEN
            exp_f := 0;
        ELSIF x =- 24174 THEN
            exp_f := 0;
        ELSIF x =- 24173 THEN
            exp_f := 0;
        ELSIF x =- 24172 THEN
            exp_f := 0;
        ELSIF x =- 24171 THEN
            exp_f := 0;
        ELSIF x =- 24170 THEN
            exp_f := 0;
        ELSIF x =- 24169 THEN
            exp_f := 0;
        ELSIF x =- 24168 THEN
            exp_f := 0;
        ELSIF x =- 24167 THEN
            exp_f := 0;
        ELSIF x =- 24166 THEN
            exp_f := 0;
        ELSIF x =- 24165 THEN
            exp_f := 0;
        ELSIF x =- 24164 THEN
            exp_f := 0;
        ELSIF x =- 24163 THEN
            exp_f := 0;
        ELSIF x =- 24162 THEN
            exp_f := 0;
        ELSIF x =- 24161 THEN
            exp_f := 0;
        ELSIF x =- 24160 THEN
            exp_f := 0;
        ELSIF x =- 24159 THEN
            exp_f := 0;
        ELSIF x =- 24158 THEN
            exp_f := 0;
        ELSIF x =- 24157 THEN
            exp_f := 0;
        ELSIF x =- 24156 THEN
            exp_f := 0;
        ELSIF x =- 24155 THEN
            exp_f := 0;
        ELSIF x =- 24154 THEN
            exp_f := 0;
        ELSIF x =- 24153 THEN
            exp_f := 0;
        ELSIF x =- 24152 THEN
            exp_f := 0;
        ELSIF x =- 24151 THEN
            exp_f := 0;
        ELSIF x =- 24150 THEN
            exp_f := 0;
        ELSIF x =- 24149 THEN
            exp_f := 0;
        ELSIF x =- 24148 THEN
            exp_f := 0;
        ELSIF x =- 24147 THEN
            exp_f := 0;
        ELSIF x =- 24146 THEN
            exp_f := 0;
        ELSIF x =- 24145 THEN
            exp_f := 0;
        ELSIF x =- 24144 THEN
            exp_f := 0;
        ELSIF x =- 24143 THEN
            exp_f := 0;
        ELSIF x =- 24142 THEN
            exp_f := 0;
        ELSIF x =- 24141 THEN
            exp_f := 0;
        ELSIF x =- 24140 THEN
            exp_f := 0;
        ELSIF x =- 24139 THEN
            exp_f := 0;
        ELSIF x =- 24138 THEN
            exp_f := 0;
        ELSIF x =- 24137 THEN
            exp_f := 0;
        ELSIF x =- 24136 THEN
            exp_f := 0;
        ELSIF x =- 24135 THEN
            exp_f := 0;
        ELSIF x =- 24134 THEN
            exp_f := 0;
        ELSIF x =- 24133 THEN
            exp_f := 0;
        ELSIF x =- 24132 THEN
            exp_f := 0;
        ELSIF x =- 24131 THEN
            exp_f := 0;
        ELSIF x =- 24130 THEN
            exp_f := 0;
        ELSIF x =- 24129 THEN
            exp_f := 0;
        ELSIF x =- 24128 THEN
            exp_f := 0;
        ELSIF x =- 24127 THEN
            exp_f := 0;
        ELSIF x =- 24126 THEN
            exp_f := 0;
        ELSIF x =- 24125 THEN
            exp_f := 0;
        ELSIF x =- 24124 THEN
            exp_f := 0;
        ELSIF x =- 24123 THEN
            exp_f := 0;
        ELSIF x =- 24122 THEN
            exp_f := 0;
        ELSIF x =- 24121 THEN
            exp_f := 0;
        ELSIF x =- 24120 THEN
            exp_f := 0;
        ELSIF x =- 24119 THEN
            exp_f := 0;
        ELSIF x =- 24118 THEN
            exp_f := 0;
        ELSIF x =- 24117 THEN
            exp_f := 0;
        ELSIF x =- 24116 THEN
            exp_f := 0;
        ELSIF x =- 24115 THEN
            exp_f := 0;
        ELSIF x =- 24114 THEN
            exp_f := 0;
        ELSIF x =- 24113 THEN
            exp_f := 0;
        ELSIF x =- 24112 THEN
            exp_f := 0;
        ELSIF x =- 24111 THEN
            exp_f := 0;
        ELSIF x =- 24110 THEN
            exp_f := 0;
        ELSIF x =- 24109 THEN
            exp_f := 0;
        ELSIF x =- 24108 THEN
            exp_f := 0;
        ELSIF x =- 24107 THEN
            exp_f := 0;
        ELSIF x =- 24106 THEN
            exp_f := 0;
        ELSIF x =- 24105 THEN
            exp_f := 0;
        ELSIF x =- 24104 THEN
            exp_f := 0;
        ELSIF x =- 24103 THEN
            exp_f := 0;
        ELSIF x =- 24102 THEN
            exp_f := 0;
        ELSIF x =- 24101 THEN
            exp_f := 0;
        ELSIF x =- 24100 THEN
            exp_f := 0;
        ELSIF x =- 24099 THEN
            exp_f := 0;
        ELSIF x =- 24098 THEN
            exp_f := 0;
        ELSIF x =- 24097 THEN
            exp_f := 0;
        ELSIF x =- 24096 THEN
            exp_f := 0;
        ELSIF x =- 24095 THEN
            exp_f := 0;
        ELSIF x =- 24094 THEN
            exp_f := 0;
        ELSIF x =- 24093 THEN
            exp_f := 0;
        ELSIF x =- 24092 THEN
            exp_f := 0;
        ELSIF x =- 24091 THEN
            exp_f := 0;
        ELSIF x =- 24090 THEN
            exp_f := 0;
        ELSIF x =- 24089 THEN
            exp_f := 0;
        ELSIF x =- 24088 THEN
            exp_f := 0;
        ELSIF x =- 24087 THEN
            exp_f := 0;
        ELSIF x =- 24086 THEN
            exp_f := 0;
        ELSIF x =- 24085 THEN
            exp_f := 0;
        ELSIF x =- 24084 THEN
            exp_f := 0;
        ELSIF x =- 24083 THEN
            exp_f := 0;
        ELSIF x =- 24082 THEN
            exp_f := 0;
        ELSIF x =- 24081 THEN
            exp_f := 0;
        ELSIF x =- 24080 THEN
            exp_f := 0;
        ELSIF x =- 24079 THEN
            exp_f := 0;
        ELSIF x =- 24078 THEN
            exp_f := 0;
        ELSIF x =- 24077 THEN
            exp_f := 0;
        ELSIF x =- 24076 THEN
            exp_f := 0;
        ELSIF x =- 24075 THEN
            exp_f := 0;
        ELSIF x =- 24074 THEN
            exp_f := 0;
        ELSIF x =- 24073 THEN
            exp_f := 0;
        ELSIF x =- 24072 THEN
            exp_f := 0;
        ELSIF x =- 24071 THEN
            exp_f := 0;
        ELSIF x =- 24070 THEN
            exp_f := 0;
        ELSIF x =- 24069 THEN
            exp_f := 0;
        ELSIF x =- 24068 THEN
            exp_f := 0;
        ELSIF x =- 24067 THEN
            exp_f := 0;
        ELSIF x =- 24066 THEN
            exp_f := 0;
        ELSIF x =- 24065 THEN
            exp_f := 0;
        ELSIF x =- 24064 THEN
            exp_f := 0;
        ELSIF x =- 24063 THEN
            exp_f := 0;
        ELSIF x =- 24062 THEN
            exp_f := 0;
        ELSIF x =- 24061 THEN
            exp_f := 0;
        ELSIF x =- 24060 THEN
            exp_f := 0;
        ELSIF x =- 24059 THEN
            exp_f := 0;
        ELSIF x =- 24058 THEN
            exp_f := 0;
        ELSIF x =- 24057 THEN
            exp_f := 0;
        ELSIF x =- 24056 THEN
            exp_f := 0;
        ELSIF x =- 24055 THEN
            exp_f := 0;
        ELSIF x =- 24054 THEN
            exp_f := 0;
        ELSIF x =- 24053 THEN
            exp_f := 0;
        ELSIF x =- 24052 THEN
            exp_f := 0;
        ELSIF x =- 24051 THEN
            exp_f := 0;
        ELSIF x =- 24050 THEN
            exp_f := 0;
        ELSIF x =- 24049 THEN
            exp_f := 0;
        ELSIF x =- 24048 THEN
            exp_f := 0;
        ELSIF x =- 24047 THEN
            exp_f := 0;
        ELSIF x =- 24046 THEN
            exp_f := 0;
        ELSIF x =- 24045 THEN
            exp_f := 0;
        ELSIF x =- 24044 THEN
            exp_f := 0;
        ELSIF x =- 24043 THEN
            exp_f := 0;
        ELSIF x =- 24042 THEN
            exp_f := 0;
        ELSIF x =- 24041 THEN
            exp_f := 0;
        ELSIF x =- 24040 THEN
            exp_f := 0;
        ELSIF x =- 24039 THEN
            exp_f := 0;
        ELSIF x =- 24038 THEN
            exp_f := 0;
        ELSIF x =- 24037 THEN
            exp_f := 0;
        ELSIF x =- 24036 THEN
            exp_f := 0;
        ELSIF x =- 24035 THEN
            exp_f := 0;
        ELSIF x =- 24034 THEN
            exp_f := 0;
        ELSIF x =- 24033 THEN
            exp_f := 0;
        ELSIF x =- 24032 THEN
            exp_f := 0;
        ELSIF x =- 24031 THEN
            exp_f := 0;
        ELSIF x =- 24030 THEN
            exp_f := 0;
        ELSIF x =- 24029 THEN
            exp_f := 0;
        ELSIF x =- 24028 THEN
            exp_f := 0;
        ELSIF x =- 24027 THEN
            exp_f := 0;
        ELSIF x =- 24026 THEN
            exp_f := 0;
        ELSIF x =- 24025 THEN
            exp_f := 0;
        ELSIF x =- 24024 THEN
            exp_f := 0;
        ELSIF x =- 24023 THEN
            exp_f := 0;
        ELSIF x =- 24022 THEN
            exp_f := 0;
        ELSIF x =- 24021 THEN
            exp_f := 0;
        ELSIF x =- 24020 THEN
            exp_f := 0;
        ELSIF x =- 24019 THEN
            exp_f := 0;
        ELSIF x =- 24018 THEN
            exp_f := 0;
        ELSIF x =- 24017 THEN
            exp_f := 0;
        ELSIF x =- 24016 THEN
            exp_f := 0;
        ELSIF x =- 24015 THEN
            exp_f := 0;
        ELSIF x =- 24014 THEN
            exp_f := 0;
        ELSIF x =- 24013 THEN
            exp_f := 0;
        ELSIF x =- 24012 THEN
            exp_f := 0;
        ELSIF x =- 24011 THEN
            exp_f := 0;
        ELSIF x =- 24010 THEN
            exp_f := 0;
        ELSIF x =- 24009 THEN
            exp_f := 0;
        ELSIF x =- 24008 THEN
            exp_f := 0;
        ELSIF x =- 24007 THEN
            exp_f := 0;
        ELSIF x =- 24006 THEN
            exp_f := 0;
        ELSIF x =- 24005 THEN
            exp_f := 0;
        ELSIF x =- 24004 THEN
            exp_f := 0;
        ELSIF x =- 24003 THEN
            exp_f := 0;
        ELSIF x =- 24002 THEN
            exp_f := 0;
        ELSIF x =- 24001 THEN
            exp_f := 0;
        ELSIF x =- 24000 THEN
            exp_f := 0;
        ELSIF x =- 23999 THEN
            exp_f := 0;
        ELSIF x =- 23998 THEN
            exp_f := 0;
        ELSIF x =- 23997 THEN
            exp_f := 0;
        ELSIF x =- 23996 THEN
            exp_f := 0;
        ELSIF x =- 23995 THEN
            exp_f := 0;
        ELSIF x =- 23994 THEN
            exp_f := 0;
        ELSIF x =- 23993 THEN
            exp_f := 0;
        ELSIF x =- 23992 THEN
            exp_f := 0;
        ELSIF x =- 23991 THEN
            exp_f := 0;
        ELSIF x =- 23990 THEN
            exp_f := 0;
        ELSIF x =- 23989 THEN
            exp_f := 0;
        ELSIF x =- 23988 THEN
            exp_f := 0;
        ELSIF x =- 23987 THEN
            exp_f := 0;
        ELSIF x =- 23986 THEN
            exp_f := 0;
        ELSIF x =- 23985 THEN
            exp_f := 0;
        ELSIF x =- 23984 THEN
            exp_f := 0;
        ELSIF x =- 23983 THEN
            exp_f := 0;
        ELSIF x =- 23982 THEN
            exp_f := 0;
        ELSIF x =- 23981 THEN
            exp_f := 0;
        ELSIF x =- 23980 THEN
            exp_f := 0;
        ELSIF x =- 23979 THEN
            exp_f := 0;
        ELSIF x =- 23978 THEN
            exp_f := 0;
        ELSIF x =- 23977 THEN
            exp_f := 0;
        ELSIF x =- 23976 THEN
            exp_f := 0;
        ELSIF x =- 23975 THEN
            exp_f := 0;
        ELSIF x =- 23974 THEN
            exp_f := 0;
        ELSIF x =- 23973 THEN
            exp_f := 0;
        ELSIF x =- 23972 THEN
            exp_f := 0;
        ELSIF x =- 23971 THEN
            exp_f := 0;
        ELSIF x =- 23970 THEN
            exp_f := 0;
        ELSIF x =- 23969 THEN
            exp_f := 0;
        ELSIF x =- 23968 THEN
            exp_f := 0;
        ELSIF x =- 23967 THEN
            exp_f := 0;
        ELSIF x =- 23966 THEN
            exp_f := 0;
        ELSIF x =- 23965 THEN
            exp_f := 0;
        ELSIF x =- 23964 THEN
            exp_f := 0;
        ELSIF x =- 23963 THEN
            exp_f := 0;
        ELSIF x =- 23962 THEN
            exp_f := 0;
        ELSIF x =- 23961 THEN
            exp_f := 0;
        ELSIF x =- 23960 THEN
            exp_f := 0;
        ELSIF x =- 23959 THEN
            exp_f := 0;
        ELSIF x =- 23958 THEN
            exp_f := 0;
        ELSIF x =- 23957 THEN
            exp_f := 0;
        ELSIF x =- 23956 THEN
            exp_f := 0;
        ELSIF x =- 23955 THEN
            exp_f := 0;
        ELSIF x =- 23954 THEN
            exp_f := 0;
        ELSIF x =- 23953 THEN
            exp_f := 0;
        ELSIF x =- 23952 THEN
            exp_f := 0;
        ELSIF x =- 23951 THEN
            exp_f := 0;
        ELSIF x =- 23950 THEN
            exp_f := 0;
        ELSIF x =- 23949 THEN
            exp_f := 0;
        ELSIF x =- 23948 THEN
            exp_f := 0;
        ELSIF x =- 23947 THEN
            exp_f := 0;
        ELSIF x =- 23946 THEN
            exp_f := 0;
        ELSIF x =- 23945 THEN
            exp_f := 0;
        ELSIF x =- 23944 THEN
            exp_f := 0;
        ELSIF x =- 23943 THEN
            exp_f := 0;
        ELSIF x =- 23942 THEN
            exp_f := 0;
        ELSIF x =- 23941 THEN
            exp_f := 0;
        ELSIF x =- 23940 THEN
            exp_f := 0;
        ELSIF x =- 23939 THEN
            exp_f := 0;
        ELSIF x =- 23938 THEN
            exp_f := 0;
        ELSIF x =- 23937 THEN
            exp_f := 0;
        ELSIF x =- 23936 THEN
            exp_f := 0;
        ELSIF x =- 23935 THEN
            exp_f := 0;
        ELSIF x =- 23934 THEN
            exp_f := 0;
        ELSIF x =- 23933 THEN
            exp_f := 0;
        ELSIF x =- 23932 THEN
            exp_f := 0;
        ELSIF x =- 23931 THEN
            exp_f := 0;
        ELSIF x =- 23930 THEN
            exp_f := 0;
        ELSIF x =- 23929 THEN
            exp_f := 0;
        ELSIF x =- 23928 THEN
            exp_f := 0;
        ELSIF x =- 23927 THEN
            exp_f := 0;
        ELSIF x =- 23926 THEN
            exp_f := 0;
        ELSIF x =- 23925 THEN
            exp_f := 0;
        ELSIF x =- 23924 THEN
            exp_f := 0;
        ELSIF x =- 23923 THEN
            exp_f := 0;
        ELSIF x =- 23922 THEN
            exp_f := 0;
        ELSIF x =- 23921 THEN
            exp_f := 0;
        ELSIF x =- 23920 THEN
            exp_f := 0;
        ELSIF x =- 23919 THEN
            exp_f := 0;
        ELSIF x =- 23918 THEN
            exp_f := 0;
        ELSIF x =- 23917 THEN
            exp_f := 0;
        ELSIF x =- 23916 THEN
            exp_f := 0;
        ELSIF x =- 23915 THEN
            exp_f := 0;
        ELSIF x =- 23914 THEN
            exp_f := 0;
        ELSIF x =- 23913 THEN
            exp_f := 0;
        ELSIF x =- 23912 THEN
            exp_f := 0;
        ELSIF x =- 23911 THEN
            exp_f := 0;
        ELSIF x =- 23910 THEN
            exp_f := 0;
        ELSIF x =- 23909 THEN
            exp_f := 0;
        ELSIF x =- 23908 THEN
            exp_f := 0;
        ELSIF x =- 23907 THEN
            exp_f := 0;
        ELSIF x =- 23906 THEN
            exp_f := 0;
        ELSIF x =- 23905 THEN
            exp_f := 0;
        ELSIF x =- 23904 THEN
            exp_f := 0;
        ELSIF x =- 23903 THEN
            exp_f := 0;
        ELSIF x =- 23902 THEN
            exp_f := 0;
        ELSIF x =- 23901 THEN
            exp_f := 0;
        ELSIF x =- 23900 THEN
            exp_f := 0;
        ELSIF x =- 23899 THEN
            exp_f := 0;
        ELSIF x =- 23898 THEN
            exp_f := 0;
        ELSIF x =- 23897 THEN
            exp_f := 0;
        ELSIF x =- 23896 THEN
            exp_f := 0;
        ELSIF x =- 23895 THEN
            exp_f := 0;
        ELSIF x =- 23894 THEN
            exp_f := 0;
        ELSIF x =- 23893 THEN
            exp_f := 0;
        ELSIF x =- 23892 THEN
            exp_f := 0;
        ELSIF x =- 23891 THEN
            exp_f := 0;
        ELSIF x =- 23890 THEN
            exp_f := 0;
        ELSIF x =- 23889 THEN
            exp_f := 0;
        ELSIF x =- 23888 THEN
            exp_f := 0;
        ELSIF x =- 23887 THEN
            exp_f := 0;
        ELSIF x =- 23886 THEN
            exp_f := 0;
        ELSIF x =- 23885 THEN
            exp_f := 0;
        ELSIF x =- 23884 THEN
            exp_f := 0;
        ELSIF x =- 23883 THEN
            exp_f := 0;
        ELSIF x =- 23882 THEN
            exp_f := 0;
        ELSIF x =- 23881 THEN
            exp_f := 0;
        ELSIF x =- 23880 THEN
            exp_f := 0;
        ELSIF x =- 23879 THEN
            exp_f := 0;
        ELSIF x =- 23878 THEN
            exp_f := 0;
        ELSIF x =- 23877 THEN
            exp_f := 0;
        ELSIF x =- 23876 THEN
            exp_f := 0;
        ELSIF x =- 23875 THEN
            exp_f := 0;
        ELSIF x =- 23874 THEN
            exp_f := 0;
        ELSIF x =- 23873 THEN
            exp_f := 0;
        ELSIF x =- 23872 THEN
            exp_f := 0;
        ELSIF x =- 23871 THEN
            exp_f := 0;
        ELSIF x =- 23870 THEN
            exp_f := 0;
        ELSIF x =- 23869 THEN
            exp_f := 0;
        ELSIF x =- 23868 THEN
            exp_f := 0;
        ELSIF x =- 23867 THEN
            exp_f := 0;
        ELSIF x =- 23866 THEN
            exp_f := 0;
        ELSIF x =- 23865 THEN
            exp_f := 0;
        ELSIF x =- 23864 THEN
            exp_f := 0;
        ELSIF x =- 23863 THEN
            exp_f := 0;
        ELSIF x =- 23862 THEN
            exp_f := 0;
        ELSIF x =- 23861 THEN
            exp_f := 0;
        ELSIF x =- 23860 THEN
            exp_f := 0;
        ELSIF x =- 23859 THEN
            exp_f := 0;
        ELSIF x =- 23858 THEN
            exp_f := 0;
        ELSIF x =- 23857 THEN
            exp_f := 0;
        ELSIF x =- 23856 THEN
            exp_f := 0;
        ELSIF x =- 23855 THEN
            exp_f := 0;
        ELSIF x =- 23854 THEN
            exp_f := 0;
        ELSIF x =- 23853 THEN
            exp_f := 0;
        ELSIF x =- 23852 THEN
            exp_f := 0;
        ELSIF x =- 23851 THEN
            exp_f := 0;
        ELSIF x =- 23850 THEN
            exp_f := 0;
        ELSIF x =- 23849 THEN
            exp_f := 0;
        ELSIF x =- 23848 THEN
            exp_f := 0;
        ELSIF x =- 23847 THEN
            exp_f := 0;
        ELSIF x =- 23846 THEN
            exp_f := 0;
        ELSIF x =- 23845 THEN
            exp_f := 0;
        ELSIF x =- 23844 THEN
            exp_f := 0;
        ELSIF x =- 23843 THEN
            exp_f := 0;
        ELSIF x =- 23842 THEN
            exp_f := 0;
        ELSIF x =- 23841 THEN
            exp_f := 0;
        ELSIF x =- 23840 THEN
            exp_f := 0;
        ELSIF x =- 23839 THEN
            exp_f := 0;
        ELSIF x =- 23838 THEN
            exp_f := 0;
        ELSIF x =- 23837 THEN
            exp_f := 0;
        ELSIF x =- 23836 THEN
            exp_f := 0;
        ELSIF x =- 23835 THEN
            exp_f := 0;
        ELSIF x =- 23834 THEN
            exp_f := 0;
        ELSIF x =- 23833 THEN
            exp_f := 0;
        ELSIF x =- 23832 THEN
            exp_f := 0;
        ELSIF x =- 23831 THEN
            exp_f := 0;
        ELSIF x =- 23830 THEN
            exp_f := 0;
        ELSIF x =- 23829 THEN
            exp_f := 0;
        ELSIF x =- 23828 THEN
            exp_f := 0;
        ELSIF x =- 23827 THEN
            exp_f := 0;
        ELSIF x =- 23826 THEN
            exp_f := 0;
        ELSIF x =- 23825 THEN
            exp_f := 0;
        ELSIF x =- 23824 THEN
            exp_f := 0;
        ELSIF x =- 23823 THEN
            exp_f := 0;
        ELSIF x =- 23822 THEN
            exp_f := 0;
        ELSIF x =- 23821 THEN
            exp_f := 0;
        ELSIF x =- 23820 THEN
            exp_f := 0;
        ELSIF x =- 23819 THEN
            exp_f := 0;
        ELSIF x =- 23818 THEN
            exp_f := 0;
        ELSIF x =- 23817 THEN
            exp_f := 0;
        ELSIF x =- 23816 THEN
            exp_f := 0;
        ELSIF x =- 23815 THEN
            exp_f := 0;
        ELSIF x =- 23814 THEN
            exp_f := 0;
        ELSIF x =- 23813 THEN
            exp_f := 0;
        ELSIF x =- 23812 THEN
            exp_f := 0;
        ELSIF x =- 23811 THEN
            exp_f := 0;
        ELSIF x =- 23810 THEN
            exp_f := 0;
        ELSIF x =- 23809 THEN
            exp_f := 0;
        ELSIF x =- 23808 THEN
            exp_f := 0;
        ELSIF x =- 23807 THEN
            exp_f := 0;
        ELSIF x =- 23806 THEN
            exp_f := 0;
        ELSIF x =- 23805 THEN
            exp_f := 0;
        ELSIF x =- 23804 THEN
            exp_f := 0;
        ELSIF x =- 23803 THEN
            exp_f := 0;
        ELSIF x =- 23802 THEN
            exp_f := 0;
        ELSIF x =- 23801 THEN
            exp_f := 0;
        ELSIF x =- 23800 THEN
            exp_f := 0;
        ELSIF x =- 23799 THEN
            exp_f := 0;
        ELSIF x =- 23798 THEN
            exp_f := 0;
        ELSIF x =- 23797 THEN
            exp_f := 0;
        ELSIF x =- 23796 THEN
            exp_f := 0;
        ELSIF x =- 23795 THEN
            exp_f := 0;
        ELSIF x =- 23794 THEN
            exp_f := 0;
        ELSIF x =- 23793 THEN
            exp_f := 0;
        ELSIF x =- 23792 THEN
            exp_f := 0;
        ELSIF x =- 23791 THEN
            exp_f := 0;
        ELSIF x =- 23790 THEN
            exp_f := 0;
        ELSIF x =- 23789 THEN
            exp_f := 0;
        ELSIF x =- 23788 THEN
            exp_f := 0;
        ELSIF x =- 23787 THEN
            exp_f := 0;
        ELSIF x =- 23786 THEN
            exp_f := 0;
        ELSIF x =- 23785 THEN
            exp_f := 0;
        ELSIF x =- 23784 THEN
            exp_f := 0;
        ELSIF x =- 23783 THEN
            exp_f := 0;
        ELSIF x =- 23782 THEN
            exp_f := 0;
        ELSIF x =- 23781 THEN
            exp_f := 0;
        ELSIF x =- 23780 THEN
            exp_f := 0;
        ELSIF x =- 23779 THEN
            exp_f := 0;
        ELSIF x =- 23778 THEN
            exp_f := 0;
        ELSIF x =- 23777 THEN
            exp_f := 0;
        ELSIF x =- 23776 THEN
            exp_f := 0;
        ELSIF x =- 23775 THEN
            exp_f := 0;
        ELSIF x =- 23774 THEN
            exp_f := 0;
        ELSIF x =- 23773 THEN
            exp_f := 0;
        ELSIF x =- 23772 THEN
            exp_f := 0;
        ELSIF x =- 23771 THEN
            exp_f := 0;
        ELSIF x =- 23770 THEN
            exp_f := 0;
        ELSIF x =- 23769 THEN
            exp_f := 0;
        ELSIF x =- 23768 THEN
            exp_f := 0;
        ELSIF x =- 23767 THEN
            exp_f := 0;
        ELSIF x =- 23766 THEN
            exp_f := 0;
        ELSIF x =- 23765 THEN
            exp_f := 0;
        ELSIF x =- 23764 THEN
            exp_f := 0;
        ELSIF x =- 23763 THEN
            exp_f := 0;
        ELSIF x =- 23762 THEN
            exp_f := 0;
        ELSIF x =- 23761 THEN
            exp_f := 0;
        ELSIF x =- 23760 THEN
            exp_f := 0;
        ELSIF x =- 23759 THEN
            exp_f := 0;
        ELSIF x =- 23758 THEN
            exp_f := 0;
        ELSIF x =- 23757 THEN
            exp_f := 0;
        ELSIF x =- 23756 THEN
            exp_f := 0;
        ELSIF x =- 23755 THEN
            exp_f := 0;
        ELSIF x =- 23754 THEN
            exp_f := 0;
        ELSIF x =- 23753 THEN
            exp_f := 0;
        ELSIF x =- 23752 THEN
            exp_f := 0;
        ELSIF x =- 23751 THEN
            exp_f := 0;
        ELSIF x =- 23750 THEN
            exp_f := 0;
        ELSIF x =- 23749 THEN
            exp_f := 0;
        ELSIF x =- 23748 THEN
            exp_f := 0;
        ELSIF x =- 23747 THEN
            exp_f := 0;
        ELSIF x =- 23746 THEN
            exp_f := 0;
        ELSIF x =- 23745 THEN
            exp_f := 0;
        ELSIF x =- 23744 THEN
            exp_f := 0;
        ELSIF x =- 23743 THEN
            exp_f := 0;
        ELSIF x =- 23742 THEN
            exp_f := 0;
        ELSIF x =- 23741 THEN
            exp_f := 0;
        ELSIF x =- 23740 THEN
            exp_f := 0;
        ELSIF x =- 23739 THEN
            exp_f := 0;
        ELSIF x =- 23738 THEN
            exp_f := 0;
        ELSIF x =- 23737 THEN
            exp_f := 0;
        ELSIF x =- 23736 THEN
            exp_f := 0;
        ELSIF x =- 23735 THEN
            exp_f := 0;
        ELSIF x =- 23734 THEN
            exp_f := 0;
        ELSIF x =- 23733 THEN
            exp_f := 0;
        ELSIF x =- 23732 THEN
            exp_f := 0;
        ELSIF x =- 23731 THEN
            exp_f := 0;
        ELSIF x =- 23730 THEN
            exp_f := 0;
        ELSIF x =- 23729 THEN
            exp_f := 0;
        ELSIF x =- 23728 THEN
            exp_f := 0;
        ELSIF x =- 23727 THEN
            exp_f := 0;
        ELSIF x =- 23726 THEN
            exp_f := 0;
        ELSIF x =- 23725 THEN
            exp_f := 0;
        ELSIF x =- 23724 THEN
            exp_f := 0;
        ELSIF x =- 23723 THEN
            exp_f := 0;
        ELSIF x =- 23722 THEN
            exp_f := 0;
        ELSIF x =- 23721 THEN
            exp_f := 0;
        ELSIF x =- 23720 THEN
            exp_f := 0;
        ELSIF x =- 23719 THEN
            exp_f := 0;
        ELSIF x =- 23718 THEN
            exp_f := 0;
        ELSIF x =- 23717 THEN
            exp_f := 0;
        ELSIF x =- 23716 THEN
            exp_f := 0;
        ELSIF x =- 23715 THEN
            exp_f := 0;
        ELSIF x =- 23714 THEN
            exp_f := 0;
        ELSIF x =- 23713 THEN
            exp_f := 0;
        ELSIF x =- 23712 THEN
            exp_f := 0;
        ELSIF x =- 23711 THEN
            exp_f := 0;
        ELSIF x =- 23710 THEN
            exp_f := 0;
        ELSIF x =- 23709 THEN
            exp_f := 0;
        ELSIF x =- 23708 THEN
            exp_f := 0;
        ELSIF x =- 23707 THEN
            exp_f := 0;
        ELSIF x =- 23706 THEN
            exp_f := 0;
        ELSIF x =- 23705 THEN
            exp_f := 0;
        ELSIF x =- 23704 THEN
            exp_f := 0;
        ELSIF x =- 23703 THEN
            exp_f := 0;
        ELSIF x =- 23702 THEN
            exp_f := 0;
        ELSIF x =- 23701 THEN
            exp_f := 0;
        ELSIF x =- 23700 THEN
            exp_f := 0;
        ELSIF x =- 23699 THEN
            exp_f := 0;
        ELSIF x =- 23698 THEN
            exp_f := 0;
        ELSIF x =- 23697 THEN
            exp_f := 0;
        ELSIF x =- 23696 THEN
            exp_f := 0;
        ELSIF x =- 23695 THEN
            exp_f := 0;
        ELSIF x =- 23694 THEN
            exp_f := 0;
        ELSIF x =- 23693 THEN
            exp_f := 0;
        ELSIF x =- 23692 THEN
            exp_f := 0;
        ELSIF x =- 23691 THEN
            exp_f := 0;
        ELSIF x =- 23690 THEN
            exp_f := 0;
        ELSIF x =- 23689 THEN
            exp_f := 0;
        ELSIF x =- 23688 THEN
            exp_f := 0;
        ELSIF x =- 23687 THEN
            exp_f := 0;
        ELSIF x =- 23686 THEN
            exp_f := 0;
        ELSIF x =- 23685 THEN
            exp_f := 0;
        ELSIF x =- 23684 THEN
            exp_f := 0;
        ELSIF x =- 23683 THEN
            exp_f := 0;
        ELSIF x =- 23682 THEN
            exp_f := 0;
        ELSIF x =- 23681 THEN
            exp_f := 0;
        ELSIF x =- 23680 THEN
            exp_f := 0;
        ELSIF x =- 23679 THEN
            exp_f := 0;
        ELSIF x =- 23678 THEN
            exp_f := 0;
        ELSIF x =- 23677 THEN
            exp_f := 0;
        ELSIF x =- 23676 THEN
            exp_f := 0;
        ELSIF x =- 23675 THEN
            exp_f := 0;
        ELSIF x =- 23674 THEN
            exp_f := 0;
        ELSIF x =- 23673 THEN
            exp_f := 0;
        ELSIF x =- 23672 THEN
            exp_f := 0;
        ELSIF x =- 23671 THEN
            exp_f := 0;
        ELSIF x =- 23670 THEN
            exp_f := 0;
        ELSIF x =- 23669 THEN
            exp_f := 0;
        ELSIF x =- 23668 THEN
            exp_f := 0;
        ELSIF x =- 23667 THEN
            exp_f := 0;
        ELSIF x =- 23666 THEN
            exp_f := 0;
        ELSIF x =- 23665 THEN
            exp_f := 0;
        ELSIF x =- 23664 THEN
            exp_f := 0;
        ELSIF x =- 23663 THEN
            exp_f := 0;
        ELSIF x =- 23662 THEN
            exp_f := 0;
        ELSIF x =- 23661 THEN
            exp_f := 0;
        ELSIF x =- 23660 THEN
            exp_f := 0;
        ELSIF x =- 23659 THEN
            exp_f := 0;
        ELSIF x =- 23658 THEN
            exp_f := 0;
        ELSIF x =- 23657 THEN
            exp_f := 0;
        ELSIF x =- 23656 THEN
            exp_f := 0;
        ELSIF x =- 23655 THEN
            exp_f := 0;
        ELSIF x =- 23654 THEN
            exp_f := 0;
        ELSIF x =- 23653 THEN
            exp_f := 0;
        ELSIF x =- 23652 THEN
            exp_f := 0;
        ELSIF x =- 23651 THEN
            exp_f := 0;
        ELSIF x =- 23650 THEN
            exp_f := 0;
        ELSIF x =- 23649 THEN
            exp_f := 0;
        ELSIF x =- 23648 THEN
            exp_f := 0;
        ELSIF x =- 23647 THEN
            exp_f := 0;
        ELSIF x =- 23646 THEN
            exp_f := 0;
        ELSIF x =- 23645 THEN
            exp_f := 0;
        ELSIF x =- 23644 THEN
            exp_f := 0;
        ELSIF x =- 23643 THEN
            exp_f := 0;
        ELSIF x =- 23642 THEN
            exp_f := 0;
        ELSIF x =- 23641 THEN
            exp_f := 0;
        ELSIF x =- 23640 THEN
            exp_f := 0;
        ELSIF x =- 23639 THEN
            exp_f := 0;
        ELSIF x =- 23638 THEN
            exp_f := 0;
        ELSIF x =- 23637 THEN
            exp_f := 0;
        ELSIF x =- 23636 THEN
            exp_f := 0;
        ELSIF x =- 23635 THEN
            exp_f := 0;
        ELSIF x =- 23634 THEN
            exp_f := 0;
        ELSIF x =- 23633 THEN
            exp_f := 0;
        ELSIF x =- 23632 THEN
            exp_f := 0;
        ELSIF x =- 23631 THEN
            exp_f := 0;
        ELSIF x =- 23630 THEN
            exp_f := 0;
        ELSIF x =- 23629 THEN
            exp_f := 0;
        ELSIF x =- 23628 THEN
            exp_f := 0;
        ELSIF x =- 23627 THEN
            exp_f := 0;
        ELSIF x =- 23626 THEN
            exp_f := 0;
        ELSIF x =- 23625 THEN
            exp_f := 0;
        ELSIF x =- 23624 THEN
            exp_f := 0;
        ELSIF x =- 23623 THEN
            exp_f := 0;
        ELSIF x =- 23622 THEN
            exp_f := 0;
        ELSIF x =- 23621 THEN
            exp_f := 0;
        ELSIF x =- 23620 THEN
            exp_f := 0;
        ELSIF x =- 23619 THEN
            exp_f := 0;
        ELSIF x =- 23618 THEN
            exp_f := 0;
        ELSIF x =- 23617 THEN
            exp_f := 0;
        ELSIF x =- 23616 THEN
            exp_f := 0;
        ELSIF x =- 23615 THEN
            exp_f := 0;
        ELSIF x =- 23614 THEN
            exp_f := 0;
        ELSIF x =- 23613 THEN
            exp_f := 0;
        ELSIF x =- 23612 THEN
            exp_f := 0;
        ELSIF x =- 23611 THEN
            exp_f := 0;
        ELSIF x =- 23610 THEN
            exp_f := 0;
        ELSIF x =- 23609 THEN
            exp_f := 0;
        ELSIF x =- 23608 THEN
            exp_f := 0;
        ELSIF x =- 23607 THEN
            exp_f := 0;
        ELSIF x =- 23606 THEN
            exp_f := 0;
        ELSIF x =- 23605 THEN
            exp_f := 0;
        ELSIF x =- 23604 THEN
            exp_f := 0;
        ELSIF x =- 23603 THEN
            exp_f := 0;
        ELSIF x =- 23602 THEN
            exp_f := 0;
        ELSIF x =- 23601 THEN
            exp_f := 0;
        ELSIF x =- 23600 THEN
            exp_f := 0;
        ELSIF x =- 23599 THEN
            exp_f := 0;
        ELSIF x =- 23598 THEN
            exp_f := 0;
        ELSIF x =- 23597 THEN
            exp_f := 0;
        ELSIF x =- 23596 THEN
            exp_f := 0;
        ELSIF x =- 23595 THEN
            exp_f := 0;
        ELSIF x =- 23594 THEN
            exp_f := 0;
        ELSIF x =- 23593 THEN
            exp_f := 0;
        ELSIF x =- 23592 THEN
            exp_f := 0;
        ELSIF x =- 23591 THEN
            exp_f := 0;
        ELSIF x =- 23590 THEN
            exp_f := 0;
        ELSIF x =- 23589 THEN
            exp_f := 0;
        ELSIF x =- 23588 THEN
            exp_f := 0;
        ELSIF x =- 23587 THEN
            exp_f := 0;
        ELSIF x =- 23586 THEN
            exp_f := 0;
        ELSIF x =- 23585 THEN
            exp_f := 0;
        ELSIF x =- 23584 THEN
            exp_f := 0;
        ELSIF x =- 23583 THEN
            exp_f := 0;
        ELSIF x =- 23582 THEN
            exp_f := 0;
        ELSIF x =- 23581 THEN
            exp_f := 0;
        ELSIF x =- 23580 THEN
            exp_f := 0;
        ELSIF x =- 23579 THEN
            exp_f := 0;
        ELSIF x =- 23578 THEN
            exp_f := 0;
        ELSIF x =- 23577 THEN
            exp_f := 0;
        ELSIF x =- 23576 THEN
            exp_f := 0;
        ELSIF x =- 23575 THEN
            exp_f := 0;
        ELSIF x =- 23574 THEN
            exp_f := 0;
        ELSIF x =- 23573 THEN
            exp_f := 0;
        ELSIF x =- 23572 THEN
            exp_f := 0;
        ELSIF x =- 23571 THEN
            exp_f := 0;
        ELSIF x =- 23570 THEN
            exp_f := 0;
        ELSIF x =- 23569 THEN
            exp_f := 0;
        ELSIF x =- 23568 THEN
            exp_f := 0;
        ELSIF x =- 23567 THEN
            exp_f := 0;
        ELSIF x =- 23566 THEN
            exp_f := 0;
        ELSIF x =- 23565 THEN
            exp_f := 0;
        ELSIF x =- 23564 THEN
            exp_f := 0;
        ELSIF x =- 23563 THEN
            exp_f := 0;
        ELSIF x =- 23562 THEN
            exp_f := 0;
        ELSIF x =- 23561 THEN
            exp_f := 0;
        ELSIF x =- 23560 THEN
            exp_f := 0;
        ELSIF x =- 23559 THEN
            exp_f := 0;
        ELSIF x =- 23558 THEN
            exp_f := 0;
        ELSIF x =- 23557 THEN
            exp_f := 0;
        ELSIF x =- 23556 THEN
            exp_f := 0;
        ELSIF x =- 23555 THEN
            exp_f := 0;
        ELSIF x =- 23554 THEN
            exp_f := 0;
        ELSIF x =- 23553 THEN
            exp_f := 0;
        ELSIF x =- 23552 THEN
            exp_f := 0;
        ELSIF x =- 23551 THEN
            exp_f := 0;
        ELSIF x =- 23550 THEN
            exp_f := 0;
        ELSIF x =- 23549 THEN
            exp_f := 0;
        ELSIF x =- 23548 THEN
            exp_f := 0;
        ELSIF x =- 23547 THEN
            exp_f := 0;
        ELSIF x =- 23546 THEN
            exp_f := 0;
        ELSIF x =- 23545 THEN
            exp_f := 0;
        ELSIF x =- 23544 THEN
            exp_f := 0;
        ELSIF x =- 23543 THEN
            exp_f := 0;
        ELSIF x =- 23542 THEN
            exp_f := 0;
        ELSIF x =- 23541 THEN
            exp_f := 0;
        ELSIF x =- 23540 THEN
            exp_f := 0;
        ELSIF x =- 23539 THEN
            exp_f := 0;
        ELSIF x =- 23538 THEN
            exp_f := 0;
        ELSIF x =- 23537 THEN
            exp_f := 0;
        ELSIF x =- 23536 THEN
            exp_f := 0;
        ELSIF x =- 23535 THEN
            exp_f := 0;
        ELSIF x =- 23534 THEN
            exp_f := 0;
        ELSIF x =- 23533 THEN
            exp_f := 0;
        ELSIF x =- 23532 THEN
            exp_f := 0;
        ELSIF x =- 23531 THEN
            exp_f := 0;
        ELSIF x =- 23530 THEN
            exp_f := 0;
        ELSIF x =- 23529 THEN
            exp_f := 0;
        ELSIF x =- 23528 THEN
            exp_f := 0;
        ELSIF x =- 23527 THEN
            exp_f := 0;
        ELSIF x =- 23526 THEN
            exp_f := 0;
        ELSIF x =- 23525 THEN
            exp_f := 0;
        ELSIF x =- 23524 THEN
            exp_f := 0;
        ELSIF x =- 23523 THEN
            exp_f := 0;
        ELSIF x =- 23522 THEN
            exp_f := 0;
        ELSIF x =- 23521 THEN
            exp_f := 0;
        ELSIF x =- 23520 THEN
            exp_f := 0;
        ELSIF x =- 23519 THEN
            exp_f := 0;
        ELSIF x =- 23518 THEN
            exp_f := 0;
        ELSIF x =- 23517 THEN
            exp_f := 0;
        ELSIF x =- 23516 THEN
            exp_f := 0;
        ELSIF x =- 23515 THEN
            exp_f := 0;
        ELSIF x =- 23514 THEN
            exp_f := 0;
        ELSIF x =- 23513 THEN
            exp_f := 0;
        ELSIF x =- 23512 THEN
            exp_f := 0;
        ELSIF x =- 23511 THEN
            exp_f := 0;
        ELSIF x =- 23510 THEN
            exp_f := 0;
        ELSIF x =- 23509 THEN
            exp_f := 0;
        ELSIF x =- 23508 THEN
            exp_f := 0;
        ELSIF x =- 23507 THEN
            exp_f := 0;
        ELSIF x =- 23506 THEN
            exp_f := 0;
        ELSIF x =- 23505 THEN
            exp_f := 0;
        ELSIF x =- 23504 THEN
            exp_f := 0;
        ELSIF x =- 23503 THEN
            exp_f := 0;
        ELSIF x =- 23502 THEN
            exp_f := 0;
        ELSIF x =- 23501 THEN
            exp_f := 0;
        ELSIF x =- 23500 THEN
            exp_f := 0;
        ELSIF x =- 23499 THEN
            exp_f := 0;
        ELSIF x =- 23498 THEN
            exp_f := 0;
        ELSIF x =- 23497 THEN
            exp_f := 0;
        ELSIF x =- 23496 THEN
            exp_f := 0;
        ELSIF x =- 23495 THEN
            exp_f := 0;
        ELSIF x =- 23494 THEN
            exp_f := 0;
        ELSIF x =- 23493 THEN
            exp_f := 0;
        ELSIF x =- 23492 THEN
            exp_f := 0;
        ELSIF x =- 23491 THEN
            exp_f := 0;
        ELSIF x =- 23490 THEN
            exp_f := 0;
        ELSIF x =- 23489 THEN
            exp_f := 0;
        ELSIF x =- 23488 THEN
            exp_f := 0;
        ELSIF x =- 23487 THEN
            exp_f := 0;
        ELSIF x =- 23486 THEN
            exp_f := 0;
        ELSIF x =- 23485 THEN
            exp_f := 0;
        ELSIF x =- 23484 THEN
            exp_f := 0;
        ELSIF x =- 23483 THEN
            exp_f := 0;
        ELSIF x =- 23482 THEN
            exp_f := 0;
        ELSIF x =- 23481 THEN
            exp_f := 0;
        ELSIF x =- 23480 THEN
            exp_f := 0;
        ELSIF x =- 23479 THEN
            exp_f := 0;
        ELSIF x =- 23478 THEN
            exp_f := 0;
        ELSIF x =- 23477 THEN
            exp_f := 0;
        ELSIF x =- 23476 THEN
            exp_f := 0;
        ELSIF x =- 23475 THEN
            exp_f := 0;
        ELSIF x =- 23474 THEN
            exp_f := 0;
        ELSIF x =- 23473 THEN
            exp_f := 0;
        ELSIF x =- 23472 THEN
            exp_f := 0;
        ELSIF x =- 23471 THEN
            exp_f := 0;
        ELSIF x =- 23470 THEN
            exp_f := 0;
        ELSIF x =- 23469 THEN
            exp_f := 0;
        ELSIF x =- 23468 THEN
            exp_f := 0;
        ELSIF x =- 23467 THEN
            exp_f := 0;
        ELSIF x =- 23466 THEN
            exp_f := 0;
        ELSIF x =- 23465 THEN
            exp_f := 0;
        ELSIF x =- 23464 THEN
            exp_f := 0;
        ELSIF x =- 23463 THEN
            exp_f := 0;
        ELSIF x =- 23462 THEN
            exp_f := 0;
        ELSIF x =- 23461 THEN
            exp_f := 0;
        ELSIF x =- 23460 THEN
            exp_f := 0;
        ELSIF x =- 23459 THEN
            exp_f := 0;
        ELSIF x =- 23458 THEN
            exp_f := 0;
        ELSIF x =- 23457 THEN
            exp_f := 0;
        ELSIF x =- 23456 THEN
            exp_f := 0;
        ELSIF x =- 23455 THEN
            exp_f := 0;
        ELSIF x =- 23454 THEN
            exp_f := 0;
        ELSIF x =- 23453 THEN
            exp_f := 0;
        ELSIF x =- 23452 THEN
            exp_f := 0;
        ELSIF x =- 23451 THEN
            exp_f := 0;
        ELSIF x =- 23450 THEN
            exp_f := 0;
        ELSIF x =- 23449 THEN
            exp_f := 0;
        ELSIF x =- 23448 THEN
            exp_f := 0;
        ELSIF x =- 23447 THEN
            exp_f := 0;
        ELSIF x =- 23446 THEN
            exp_f := 0;
        ELSIF x =- 23445 THEN
            exp_f := 0;
        ELSIF x =- 23444 THEN
            exp_f := 0;
        ELSIF x =- 23443 THEN
            exp_f := 0;
        ELSIF x =- 23442 THEN
            exp_f := 0;
        ELSIF x =- 23441 THEN
            exp_f := 0;
        ELSIF x =- 23440 THEN
            exp_f := 0;
        ELSIF x =- 23439 THEN
            exp_f := 0;
        ELSIF x =- 23438 THEN
            exp_f := 0;
        ELSIF x =- 23437 THEN
            exp_f := 0;
        ELSIF x =- 23436 THEN
            exp_f := 0;
        ELSIF x =- 23435 THEN
            exp_f := 0;
        ELSIF x =- 23434 THEN
            exp_f := 0;
        ELSIF x =- 23433 THEN
            exp_f := 0;
        ELSIF x =- 23432 THEN
            exp_f := 0;
        ELSIF x =- 23431 THEN
            exp_f := 0;
        ELSIF x =- 23430 THEN
            exp_f := 0;
        ELSIF x =- 23429 THEN
            exp_f := 0;
        ELSIF x =- 23428 THEN
            exp_f := 0;
        ELSIF x =- 23427 THEN
            exp_f := 0;
        ELSIF x =- 23426 THEN
            exp_f := 0;
        ELSIF x =- 23425 THEN
            exp_f := 0;
        ELSIF x =- 23424 THEN
            exp_f := 0;
        ELSIF x =- 23423 THEN
            exp_f := 0;
        ELSIF x =- 23422 THEN
            exp_f := 0;
        ELSIF x =- 23421 THEN
            exp_f := 0;
        ELSIF x =- 23420 THEN
            exp_f := 0;
        ELSIF x =- 23419 THEN
            exp_f := 0;
        ELSIF x =- 23418 THEN
            exp_f := 0;
        ELSIF x =- 23417 THEN
            exp_f := 0;
        ELSIF x =- 23416 THEN
            exp_f := 0;
        ELSIF x =- 23415 THEN
            exp_f := 0;
        ELSIF x =- 23414 THEN
            exp_f := 0;
        ELSIF x =- 23413 THEN
            exp_f := 0;
        ELSIF x =- 23412 THEN
            exp_f := 0;
        ELSIF x =- 23411 THEN
            exp_f := 0;
        ELSIF x =- 23410 THEN
            exp_f := 0;
        ELSIF x =- 23409 THEN
            exp_f := 0;
        ELSIF x =- 23408 THEN
            exp_f := 0;
        ELSIF x =- 23407 THEN
            exp_f := 0;
        ELSIF x =- 23406 THEN
            exp_f := 0;
        ELSIF x =- 23405 THEN
            exp_f := 0;
        ELSIF x =- 23404 THEN
            exp_f := 0;
        ELSIF x =- 23403 THEN
            exp_f := 0;
        ELSIF x =- 23402 THEN
            exp_f := 0;
        ELSIF x =- 23401 THEN
            exp_f := 0;
        ELSIF x =- 23400 THEN
            exp_f := 0;
        ELSIF x =- 23399 THEN
            exp_f := 0;
        ELSIF x =- 23398 THEN
            exp_f := 0;
        ELSIF x =- 23397 THEN
            exp_f := 0;
        ELSIF x =- 23396 THEN
            exp_f := 0;
        ELSIF x =- 23395 THEN
            exp_f := 0;
        ELSIF x =- 23394 THEN
            exp_f := 0;
        ELSIF x =- 23393 THEN
            exp_f := 0;
        ELSIF x =- 23392 THEN
            exp_f := 0;
        ELSIF x =- 23391 THEN
            exp_f := 0;
        ELSIF x =- 23390 THEN
            exp_f := 0;
        ELSIF x =- 23389 THEN
            exp_f := 0;
        ELSIF x =- 23388 THEN
            exp_f := 0;
        ELSIF x =- 23387 THEN
            exp_f := 0;
        ELSIF x =- 23386 THEN
            exp_f := 0;
        ELSIF x =- 23385 THEN
            exp_f := 0;
        ELSIF x =- 23384 THEN
            exp_f := 0;
        ELSIF x =- 23383 THEN
            exp_f := 0;
        ELSIF x =- 23382 THEN
            exp_f := 0;
        ELSIF x =- 23381 THEN
            exp_f := 0;
        ELSIF x =- 23380 THEN
            exp_f := 0;
        ELSIF x =- 23379 THEN
            exp_f := 0;
        ELSIF x =- 23378 THEN
            exp_f := 0;
        ELSIF x =- 23377 THEN
            exp_f := 0;
        ELSIF x =- 23376 THEN
            exp_f := 0;
        ELSIF x =- 23375 THEN
            exp_f := 0;
        ELSIF x =- 23374 THEN
            exp_f := 0;
        ELSIF x =- 23373 THEN
            exp_f := 0;
        ELSIF x =- 23372 THEN
            exp_f := 0;
        ELSIF x =- 23371 THEN
            exp_f := 0;
        ELSIF x =- 23370 THEN
            exp_f := 0;
        ELSIF x =- 23369 THEN
            exp_f := 0;
        ELSIF x =- 23368 THEN
            exp_f := 0;
        ELSIF x =- 23367 THEN
            exp_f := 0;
        ELSIF x =- 23366 THEN
            exp_f := 0;
        ELSIF x =- 23365 THEN
            exp_f := 0;
        ELSIF x =- 23364 THEN
            exp_f := 0;
        ELSIF x =- 23363 THEN
            exp_f := 0;
        ELSIF x =- 23362 THEN
            exp_f := 0;
        ELSIF x =- 23361 THEN
            exp_f := 0;
        ELSIF x =- 23360 THEN
            exp_f := 0;
        ELSIF x =- 23359 THEN
            exp_f := 0;
        ELSIF x =- 23358 THEN
            exp_f := 0;
        ELSIF x =- 23357 THEN
            exp_f := 0;
        ELSIF x =- 23356 THEN
            exp_f := 0;
        ELSIF x =- 23355 THEN
            exp_f := 0;
        ELSIF x =- 23354 THEN
            exp_f := 0;
        ELSIF x =- 23353 THEN
            exp_f := 0;
        ELSIF x =- 23352 THEN
            exp_f := 0;
        ELSIF x =- 23351 THEN
            exp_f := 0;
        ELSIF x =- 23350 THEN
            exp_f := 0;
        ELSIF x =- 23349 THEN
            exp_f := 0;
        ELSIF x =- 23348 THEN
            exp_f := 0;
        ELSIF x =- 23347 THEN
            exp_f := 0;
        ELSIF x =- 23346 THEN
            exp_f := 0;
        ELSIF x =- 23345 THEN
            exp_f := 0;
        ELSIF x =- 23344 THEN
            exp_f := 0;
        ELSIF x =- 23343 THEN
            exp_f := 0;
        ELSIF x =- 23342 THEN
            exp_f := 0;
        ELSIF x =- 23341 THEN
            exp_f := 0;
        ELSIF x =- 23340 THEN
            exp_f := 0;
        ELSIF x =- 23339 THEN
            exp_f := 0;
        ELSIF x =- 23338 THEN
            exp_f := 0;
        ELSIF x =- 23337 THEN
            exp_f := 0;
        ELSIF x =- 23336 THEN
            exp_f := 0;
        ELSIF x =- 23335 THEN
            exp_f := 0;
        ELSIF x =- 23334 THEN
            exp_f := 0;
        ELSIF x =- 23333 THEN
            exp_f := 0;
        ELSIF x =- 23332 THEN
            exp_f := 0;
        ELSIF x =- 23331 THEN
            exp_f := 0;
        ELSIF x =- 23330 THEN
            exp_f := 0;
        ELSIF x =- 23329 THEN
            exp_f := 0;
        ELSIF x =- 23328 THEN
            exp_f := 0;
        ELSIF x =- 23327 THEN
            exp_f := 0;
        ELSIF x =- 23326 THEN
            exp_f := 0;
        ELSIF x =- 23325 THEN
            exp_f := 0;
        ELSIF x =- 23324 THEN
            exp_f := 0;
        ELSIF x =- 23323 THEN
            exp_f := 0;
        ELSIF x =- 23322 THEN
            exp_f := 0;
        ELSIF x =- 23321 THEN
            exp_f := 0;
        ELSIF x =- 23320 THEN
            exp_f := 0;
        ELSIF x =- 23319 THEN
            exp_f := 0;
        ELSIF x =- 23318 THEN
            exp_f := 0;
        ELSIF x =- 23317 THEN
            exp_f := 0;
        ELSIF x =- 23316 THEN
            exp_f := 0;
        ELSIF x =- 23315 THEN
            exp_f := 0;
        ELSIF x =- 23314 THEN
            exp_f := 0;
        ELSIF x =- 23313 THEN
            exp_f := 0;
        ELSIF x =- 23312 THEN
            exp_f := 0;
        ELSIF x =- 23311 THEN
            exp_f := 0;
        ELSIF x =- 23310 THEN
            exp_f := 0;
        ELSIF x =- 23309 THEN
            exp_f := 0;
        ELSIF x =- 23308 THEN
            exp_f := 0;
        ELSIF x =- 23307 THEN
            exp_f := 0;
        ELSIF x =- 23306 THEN
            exp_f := 0;
        ELSIF x =- 23305 THEN
            exp_f := 0;
        ELSIF x =- 23304 THEN
            exp_f := 0;
        ELSIF x =- 23303 THEN
            exp_f := 0;
        ELSIF x =- 23302 THEN
            exp_f := 0;
        ELSIF x =- 23301 THEN
            exp_f := 0;
        ELSIF x =- 23300 THEN
            exp_f := 0;
        ELSIF x =- 23299 THEN
            exp_f := 0;
        ELSIF x =- 23298 THEN
            exp_f := 0;
        ELSIF x =- 23297 THEN
            exp_f := 0;
        ELSIF x =- 23296 THEN
            exp_f := 0;
        ELSIF x =- 23295 THEN
            exp_f := 0;
        ELSIF x =- 23294 THEN
            exp_f := 0;
        ELSIF x =- 23293 THEN
            exp_f := 0;
        ELSIF x =- 23292 THEN
            exp_f := 0;
        ELSIF x =- 23291 THEN
            exp_f := 0;
        ELSIF x =- 23290 THEN
            exp_f := 0;
        ELSIF x =- 23289 THEN
            exp_f := 0;
        ELSIF x =- 23288 THEN
            exp_f := 0;
        ELSIF x =- 23287 THEN
            exp_f := 0;
        ELSIF x =- 23286 THEN
            exp_f := 0;
        ELSIF x =- 23285 THEN
            exp_f := 0;
        ELSIF x =- 23284 THEN
            exp_f := 0;
        ELSIF x =- 23283 THEN
            exp_f := 0;
        ELSIF x =- 23282 THEN
            exp_f := 0;
        ELSIF x =- 23281 THEN
            exp_f := 0;
        ELSIF x =- 23280 THEN
            exp_f := 0;
        ELSIF x =- 23279 THEN
            exp_f := 0;
        ELSIF x =- 23278 THEN
            exp_f := 0;
        ELSIF x =- 23277 THEN
            exp_f := 0;
        ELSIF x =- 23276 THEN
            exp_f := 0;
        ELSIF x =- 23275 THEN
            exp_f := 0;
        ELSIF x =- 23274 THEN
            exp_f := 0;
        ELSIF x =- 23273 THEN
            exp_f := 0;
        ELSIF x =- 23272 THEN
            exp_f := 0;
        ELSIF x =- 23271 THEN
            exp_f := 0;
        ELSIF x =- 23270 THEN
            exp_f := 0;
        ELSIF x =- 23269 THEN
            exp_f := 0;
        ELSIF x =- 23268 THEN
            exp_f := 0;
        ELSIF x =- 23267 THEN
            exp_f := 0;
        ELSIF x =- 23266 THEN
            exp_f := 0;
        ELSIF x =- 23265 THEN
            exp_f := 0;
        ELSIF x =- 23264 THEN
            exp_f := 0;
        ELSIF x =- 23263 THEN
            exp_f := 0;
        ELSIF x =- 23262 THEN
            exp_f := 0;
        ELSIF x =- 23261 THEN
            exp_f := 0;
        ELSIF x =- 23260 THEN
            exp_f := 0;
        ELSIF x =- 23259 THEN
            exp_f := 0;
        ELSIF x =- 23258 THEN
            exp_f := 0;
        ELSIF x =- 23257 THEN
            exp_f := 0;
        ELSIF x =- 23256 THEN
            exp_f := 0;
        ELSIF x =- 23255 THEN
            exp_f := 0;
        ELSIF x =- 23254 THEN
            exp_f := 0;
        ELSIF x =- 23253 THEN
            exp_f := 0;
        ELSIF x =- 23252 THEN
            exp_f := 0;
        ELSIF x =- 23251 THEN
            exp_f := 0;
        ELSIF x =- 23250 THEN
            exp_f := 0;
        ELSIF x =- 23249 THEN
            exp_f := 0;
        ELSIF x =- 23248 THEN
            exp_f := 0;
        ELSIF x =- 23247 THEN
            exp_f := 0;
        ELSIF x =- 23246 THEN
            exp_f := 0;
        ELSIF x =- 23245 THEN
            exp_f := 0;
        ELSIF x =- 23244 THEN
            exp_f := 0;
        ELSIF x =- 23243 THEN
            exp_f := 0;
        ELSIF x =- 23242 THEN
            exp_f := 0;
        ELSIF x =- 23241 THEN
            exp_f := 0;
        ELSIF x =- 23240 THEN
            exp_f := 0;
        ELSIF x =- 23239 THEN
            exp_f := 0;
        ELSIF x =- 23238 THEN
            exp_f := 0;
        ELSIF x =- 23237 THEN
            exp_f := 0;
        ELSIF x =- 23236 THEN
            exp_f := 0;
        ELSIF x =- 23235 THEN
            exp_f := 0;
        ELSIF x =- 23234 THEN
            exp_f := 0;
        ELSIF x =- 23233 THEN
            exp_f := 0;
        ELSIF x =- 23232 THEN
            exp_f := 0;
        ELSIF x =- 23231 THEN
            exp_f := 0;
        ELSIF x =- 23230 THEN
            exp_f := 0;
        ELSIF x =- 23229 THEN
            exp_f := 0;
        ELSIF x =- 23228 THEN
            exp_f := 0;
        ELSIF x =- 23227 THEN
            exp_f := 0;
        ELSIF x =- 23226 THEN
            exp_f := 0;
        ELSIF x =- 23225 THEN
            exp_f := 0;
        ELSIF x =- 23224 THEN
            exp_f := 0;
        ELSIF x =- 23223 THEN
            exp_f := 0;
        ELSIF x =- 23222 THEN
            exp_f := 0;
        ELSIF x =- 23221 THEN
            exp_f := 0;
        ELSIF x =- 23220 THEN
            exp_f := 0;
        ELSIF x =- 23219 THEN
            exp_f := 0;
        ELSIF x =- 23218 THEN
            exp_f := 0;
        ELSIF x =- 23217 THEN
            exp_f := 0;
        ELSIF x =- 23216 THEN
            exp_f := 0;
        ELSIF x =- 23215 THEN
            exp_f := 0;
        ELSIF x =- 23214 THEN
            exp_f := 0;
        ELSIF x =- 23213 THEN
            exp_f := 0;
        ELSIF x =- 23212 THEN
            exp_f := 0;
        ELSIF x =- 23211 THEN
            exp_f := 0;
        ELSIF x =- 23210 THEN
            exp_f := 0;
        ELSIF x =- 23209 THEN
            exp_f := 0;
        ELSIF x =- 23208 THEN
            exp_f := 0;
        ELSIF x =- 23207 THEN
            exp_f := 0;
        ELSIF x =- 23206 THEN
            exp_f := 0;
        ELSIF x =- 23205 THEN
            exp_f := 0;
        ELSIF x =- 23204 THEN
            exp_f := 0;
        ELSIF x =- 23203 THEN
            exp_f := 0;
        ELSIF x =- 23202 THEN
            exp_f := 0;
        ELSIF x =- 23201 THEN
            exp_f := 0;
        ELSIF x =- 23200 THEN
            exp_f := 0;
        ELSIF x =- 23199 THEN
            exp_f := 0;
        ELSIF x =- 23198 THEN
            exp_f := 0;
        ELSIF x =- 23197 THEN
            exp_f := 0;
        ELSIF x =- 23196 THEN
            exp_f := 0;
        ELSIF x =- 23195 THEN
            exp_f := 0;
        ELSIF x =- 23194 THEN
            exp_f := 0;
        ELSIF x =- 23193 THEN
            exp_f := 0;
        ELSIF x =- 23192 THEN
            exp_f := 0;
        ELSIF x =- 23191 THEN
            exp_f := 0;
        ELSIF x =- 23190 THEN
            exp_f := 0;
        ELSIF x =- 23189 THEN
            exp_f := 0;
        ELSIF x =- 23188 THEN
            exp_f := 0;
        ELSIF x =- 23187 THEN
            exp_f := 0;
        ELSIF x =- 23186 THEN
            exp_f := 0;
        ELSIF x =- 23185 THEN
            exp_f := 0;
        ELSIF x =- 23184 THEN
            exp_f := 0;
        ELSIF x =- 23183 THEN
            exp_f := 0;
        ELSIF x =- 23182 THEN
            exp_f := 0;
        ELSIF x =- 23181 THEN
            exp_f := 0;
        ELSIF x =- 23180 THEN
            exp_f := 0;
        ELSIF x =- 23179 THEN
            exp_f := 0;
        ELSIF x =- 23178 THEN
            exp_f := 0;
        ELSIF x =- 23177 THEN
            exp_f := 0;
        ELSIF x =- 23176 THEN
            exp_f := 0;
        ELSIF x =- 23175 THEN
            exp_f := 0;
        ELSIF x =- 23174 THEN
            exp_f := 0;
        ELSIF x =- 23173 THEN
            exp_f := 0;
        ELSIF x =- 23172 THEN
            exp_f := 0;
        ELSIF x =- 23171 THEN
            exp_f := 0;
        ELSIF x =- 23170 THEN
            exp_f := 0;
        ELSIF x =- 23169 THEN
            exp_f := 0;
        ELSIF x =- 23168 THEN
            exp_f := 0;
        ELSIF x =- 23167 THEN
            exp_f := 0;
        ELSIF x =- 23166 THEN
            exp_f := 0;
        ELSIF x =- 23165 THEN
            exp_f := 0;
        ELSIF x =- 23164 THEN
            exp_f := 0;
        ELSIF x =- 23163 THEN
            exp_f := 0;
        ELSIF x =- 23162 THEN
            exp_f := 0;
        ELSIF x =- 23161 THEN
            exp_f := 0;
        ELSIF x =- 23160 THEN
            exp_f := 0;
        ELSIF x =- 23159 THEN
            exp_f := 0;
        ELSIF x =- 23158 THEN
            exp_f := 0;
        ELSIF x =- 23157 THEN
            exp_f := 0;
        ELSIF x =- 23156 THEN
            exp_f := 0;
        ELSIF x =- 23155 THEN
            exp_f := 0;
        ELSIF x =- 23154 THEN
            exp_f := 0;
        ELSIF x =- 23153 THEN
            exp_f := 0;
        ELSIF x =- 23152 THEN
            exp_f := 0;
        ELSIF x =- 23151 THEN
            exp_f := 0;
        ELSIF x =- 23150 THEN
            exp_f := 0;
        ELSIF x =- 23149 THEN
            exp_f := 0;
        ELSIF x =- 23148 THEN
            exp_f := 0;
        ELSIF x =- 23147 THEN
            exp_f := 0;
        ELSIF x =- 23146 THEN
            exp_f := 0;
        ELSIF x =- 23145 THEN
            exp_f := 0;
        ELSIF x =- 23144 THEN
            exp_f := 0;
        ELSIF x =- 23143 THEN
            exp_f := 0;
        ELSIF x =- 23142 THEN
            exp_f := 0;
        ELSIF x =- 23141 THEN
            exp_f := 0;
        ELSIF x =- 23140 THEN
            exp_f := 0;
        ELSIF x =- 23139 THEN
            exp_f := 0;
        ELSIF x =- 23138 THEN
            exp_f := 0;
        ELSIF x =- 23137 THEN
            exp_f := 0;
        ELSIF x =- 23136 THEN
            exp_f := 0;
        ELSIF x =- 23135 THEN
            exp_f := 0;
        ELSIF x =- 23134 THEN
            exp_f := 0;
        ELSIF x =- 23133 THEN
            exp_f := 0;
        ELSIF x =- 23132 THEN
            exp_f := 0;
        ELSIF x =- 23131 THEN
            exp_f := 0;
        ELSIF x =- 23130 THEN
            exp_f := 0;
        ELSIF x =- 23129 THEN
            exp_f := 0;
        ELSIF x =- 23128 THEN
            exp_f := 0;
        ELSIF x =- 23127 THEN
            exp_f := 0;
        ELSIF x =- 23126 THEN
            exp_f := 0;
        ELSIF x =- 23125 THEN
            exp_f := 0;
        ELSIF x =- 23124 THEN
            exp_f := 0;
        ELSIF x =- 23123 THEN
            exp_f := 0;
        ELSIF x =- 23122 THEN
            exp_f := 0;
        ELSIF x =- 23121 THEN
            exp_f := 0;
        ELSIF x =- 23120 THEN
            exp_f := 0;
        ELSIF x =- 23119 THEN
            exp_f := 0;
        ELSIF x =- 23118 THEN
            exp_f := 0;
        ELSIF x =- 23117 THEN
            exp_f := 0;
        ELSIF x =- 23116 THEN
            exp_f := 0;
        ELSIF x =- 23115 THEN
            exp_f := 0;
        ELSIF x =- 23114 THEN
            exp_f := 0;
        ELSIF x =- 23113 THEN
            exp_f := 0;
        ELSIF x =- 23112 THEN
            exp_f := 0;
        ELSIF x =- 23111 THEN
            exp_f := 0;
        ELSIF x =- 23110 THEN
            exp_f := 0;
        ELSIF x =- 23109 THEN
            exp_f := 0;
        ELSIF x =- 23108 THEN
            exp_f := 0;
        ELSIF x =- 23107 THEN
            exp_f := 0;
        ELSIF x =- 23106 THEN
            exp_f := 0;
        ELSIF x =- 23105 THEN
            exp_f := 0;
        ELSIF x =- 23104 THEN
            exp_f := 0;
        ELSIF x =- 23103 THEN
            exp_f := 0;
        ELSIF x =- 23102 THEN
            exp_f := 0;
        ELSIF x =- 23101 THEN
            exp_f := 0;
        ELSIF x =- 23100 THEN
            exp_f := 0;
        ELSIF x =- 23099 THEN
            exp_f := 0;
        ELSIF x =- 23098 THEN
            exp_f := 0;
        ELSIF x =- 23097 THEN
            exp_f := 0;
        ELSIF x =- 23096 THEN
            exp_f := 0;
        ELSIF x =- 23095 THEN
            exp_f := 0;
        ELSIF x =- 23094 THEN
            exp_f := 0;
        ELSIF x =- 23093 THEN
            exp_f := 0;
        ELSIF x =- 23092 THEN
            exp_f := 0;
        ELSIF x =- 23091 THEN
            exp_f := 0;
        ELSIF x =- 23090 THEN
            exp_f := 0;
        ELSIF x =- 23089 THEN
            exp_f := 0;
        ELSIF x =- 23088 THEN
            exp_f := 0;
        ELSIF x =- 23087 THEN
            exp_f := 0;
        ELSIF x =- 23086 THEN
            exp_f := 0;
        ELSIF x =- 23085 THEN
            exp_f := 0;
        ELSIF x =- 23084 THEN
            exp_f := 0;
        ELSIF x =- 23083 THEN
            exp_f := 0;
        ELSIF x =- 23082 THEN
            exp_f := 0;
        ELSIF x =- 23081 THEN
            exp_f := 0;
        ELSIF x =- 23080 THEN
            exp_f := 0;
        ELSIF x =- 23079 THEN
            exp_f := 0;
        ELSIF x =- 23078 THEN
            exp_f := 0;
        ELSIF x =- 23077 THEN
            exp_f := 0;
        ELSIF x =- 23076 THEN
            exp_f := 0;
        ELSIF x =- 23075 THEN
            exp_f := 0;
        ELSIF x =- 23074 THEN
            exp_f := 0;
        ELSIF x =- 23073 THEN
            exp_f := 0;
        ELSIF x =- 23072 THEN
            exp_f := 0;
        ELSIF x =- 23071 THEN
            exp_f := 0;
        ELSIF x =- 23070 THEN
            exp_f := 0;
        ELSIF x =- 23069 THEN
            exp_f := 0;
        ELSIF x =- 23068 THEN
            exp_f := 0;
        ELSIF x =- 23067 THEN
            exp_f := 0;
        ELSIF x =- 23066 THEN
            exp_f := 0;
        ELSIF x =- 23065 THEN
            exp_f := 0;
        ELSIF x =- 23064 THEN
            exp_f := 0;
        ELSIF x =- 23063 THEN
            exp_f := 0;
        ELSIF x =- 23062 THEN
            exp_f := 0;
        ELSIF x =- 23061 THEN
            exp_f := 0;
        ELSIF x =- 23060 THEN
            exp_f := 0;
        ELSIF x =- 23059 THEN
            exp_f := 0;
        ELSIF x =- 23058 THEN
            exp_f := 0;
        ELSIF x =- 23057 THEN
            exp_f := 0;
        ELSIF x =- 23056 THEN
            exp_f := 0;
        ELSIF x =- 23055 THEN
            exp_f := 0;
        ELSIF x =- 23054 THEN
            exp_f := 0;
        ELSIF x =- 23053 THEN
            exp_f := 0;
        ELSIF x =- 23052 THEN
            exp_f := 0;
        ELSIF x =- 23051 THEN
            exp_f := 0;
        ELSIF x =- 23050 THEN
            exp_f := 0;
        ELSIF x =- 23049 THEN
            exp_f := 0;
        ELSIF x =- 23048 THEN
            exp_f := 0;
        ELSIF x =- 23047 THEN
            exp_f := 0;
        ELSIF x =- 23046 THEN
            exp_f := 0;
        ELSIF x =- 23045 THEN
            exp_f := 0;
        ELSIF x =- 23044 THEN
            exp_f := 0;
        ELSIF x =- 23043 THEN
            exp_f := 0;
        ELSIF x =- 23042 THEN
            exp_f := 0;
        ELSIF x =- 23041 THEN
            exp_f := 0;
        ELSIF x =- 23040 THEN
            exp_f := 0;
        ELSIF x =- 23039 THEN
            exp_f := 0;
        ELSIF x =- 23038 THEN
            exp_f := 0;
        ELSIF x =- 23037 THEN
            exp_f := 0;
        ELSIF x =- 23036 THEN
            exp_f := 0;
        ELSIF x =- 23035 THEN
            exp_f := 0;
        ELSIF x =- 23034 THEN
            exp_f := 0;
        ELSIF x =- 23033 THEN
            exp_f := 0;
        ELSIF x =- 23032 THEN
            exp_f := 0;
        ELSIF x =- 23031 THEN
            exp_f := 0;
        ELSIF x =- 23030 THEN
            exp_f := 0;
        ELSIF x =- 23029 THEN
            exp_f := 0;
        ELSIF x =- 23028 THEN
            exp_f := 0;
        ELSIF x =- 23027 THEN
            exp_f := 0;
        ELSIF x =- 23026 THEN
            exp_f := 0;
        ELSIF x =- 23025 THEN
            exp_f := 0;
        ELSIF x =- 23024 THEN
            exp_f := 0;
        ELSIF x =- 23023 THEN
            exp_f := 0;
        ELSIF x =- 23022 THEN
            exp_f := 0;
        ELSIF x =- 23021 THEN
            exp_f := 0;
        ELSIF x =- 23020 THEN
            exp_f := 0;
        ELSIF x =- 23019 THEN
            exp_f := 0;
        ELSIF x =- 23018 THEN
            exp_f := 0;
        ELSIF x =- 23017 THEN
            exp_f := 0;
        ELSIF x =- 23016 THEN
            exp_f := 0;
        ELSIF x =- 23015 THEN
            exp_f := 0;
        ELSIF x =- 23014 THEN
            exp_f := 0;
        ELSIF x =- 23013 THEN
            exp_f := 0;
        ELSIF x =- 23012 THEN
            exp_f := 0;
        ELSIF x =- 23011 THEN
            exp_f := 0;
        ELSIF x =- 23010 THEN
            exp_f := 0;
        ELSIF x =- 23009 THEN
            exp_f := 0;
        ELSIF x =- 23008 THEN
            exp_f := 0;
        ELSIF x =- 23007 THEN
            exp_f := 0;
        ELSIF x =- 23006 THEN
            exp_f := 0;
        ELSIF x =- 23005 THEN
            exp_f := 0;
        ELSIF x =- 23004 THEN
            exp_f := 0;
        ELSIF x =- 23003 THEN
            exp_f := 0;
        ELSIF x =- 23002 THEN
            exp_f := 0;
        ELSIF x =- 23001 THEN
            exp_f := 0;
        ELSIF x =- 23000 THEN
            exp_f := 0;
        ELSIF x =- 22999 THEN
            exp_f := 0;
        ELSIF x =- 22998 THEN
            exp_f := 0;
        ELSIF x =- 22997 THEN
            exp_f := 0;
        ELSIF x =- 22996 THEN
            exp_f := 0;
        ELSIF x =- 22995 THEN
            exp_f := 0;
        ELSIF x =- 22994 THEN
            exp_f := 0;
        ELSIF x =- 22993 THEN
            exp_f := 0;
        ELSIF x =- 22992 THEN
            exp_f := 0;
        ELSIF x =- 22991 THEN
            exp_f := 0;
        ELSIF x =- 22990 THEN
            exp_f := 0;
        ELSIF x =- 22989 THEN
            exp_f := 0;
        ELSIF x =- 22988 THEN
            exp_f := 0;
        ELSIF x =- 22987 THEN
            exp_f := 0;
        ELSIF x =- 22986 THEN
            exp_f := 0;
        ELSIF x =- 22985 THEN
            exp_f := 0;
        ELSIF x =- 22984 THEN
            exp_f := 0;
        ELSIF x =- 22983 THEN
            exp_f := 0;
        ELSIF x =- 22982 THEN
            exp_f := 0;
        ELSIF x =- 22981 THEN
            exp_f := 0;
        ELSIF x =- 22980 THEN
            exp_f := 0;
        ELSIF x =- 22979 THEN
            exp_f := 0;
        ELSIF x =- 22978 THEN
            exp_f := 0;
        ELSIF x =- 22977 THEN
            exp_f := 0;
        ELSIF x =- 22976 THEN
            exp_f := 0;
        ELSIF x =- 22975 THEN
            exp_f := 0;
        ELSIF x =- 22974 THEN
            exp_f := 0;
        ELSIF x =- 22973 THEN
            exp_f := 0;
        ELSIF x =- 22972 THEN
            exp_f := 0;
        ELSIF x =- 22971 THEN
            exp_f := 0;
        ELSIF x =- 22970 THEN
            exp_f := 0;
        ELSIF x =- 22969 THEN
            exp_f := 0;
        ELSIF x =- 22968 THEN
            exp_f := 0;
        ELSIF x =- 22967 THEN
            exp_f := 0;
        ELSIF x =- 22966 THEN
            exp_f := 0;
        ELSIF x =- 22965 THEN
            exp_f := 0;
        ELSIF x =- 22964 THEN
            exp_f := 0;
        ELSIF x =- 22963 THEN
            exp_f := 0;
        ELSIF x =- 22962 THEN
            exp_f := 0;
        ELSIF x =- 22961 THEN
            exp_f := 0;
        ELSIF x =- 22960 THEN
            exp_f := 0;
        ELSIF x =- 22959 THEN
            exp_f := 0;
        ELSIF x =- 22958 THEN
            exp_f := 0;
        ELSIF x =- 22957 THEN
            exp_f := 0;
        ELSIF x =- 22956 THEN
            exp_f := 0;
        ELSIF x =- 22955 THEN
            exp_f := 0;
        ELSIF x =- 22954 THEN
            exp_f := 0;
        ELSIF x =- 22953 THEN
            exp_f := 0;
        ELSIF x =- 22952 THEN
            exp_f := 0;
        ELSIF x =- 22951 THEN
            exp_f := 0;
        ELSIF x =- 22950 THEN
            exp_f := 0;
        ELSIF x =- 22949 THEN
            exp_f := 0;
        ELSIF x =- 22948 THEN
            exp_f := 0;
        ELSIF x =- 22947 THEN
            exp_f := 0;
        ELSIF x =- 22946 THEN
            exp_f := 0;
        ELSIF x =- 22945 THEN
            exp_f := 0;
        ELSIF x =- 22944 THEN
            exp_f := 0;
        ELSIF x =- 22943 THEN
            exp_f := 0;
        ELSIF x =- 22942 THEN
            exp_f := 0;
        ELSIF x =- 22941 THEN
            exp_f := 0;
        ELSIF x =- 22940 THEN
            exp_f := 0;
        ELSIF x =- 22939 THEN
            exp_f := 0;
        ELSIF x =- 22938 THEN
            exp_f := 0;
        ELSIF x =- 22937 THEN
            exp_f := 0;
        ELSIF x =- 22936 THEN
            exp_f := 0;
        ELSIF x =- 22935 THEN
            exp_f := 0;
        ELSIF x =- 22934 THEN
            exp_f := 0;
        ELSIF x =- 22933 THEN
            exp_f := 0;
        ELSIF x =- 22932 THEN
            exp_f := 0;
        ELSIF x =- 22931 THEN
            exp_f := 0;
        ELSIF x =- 22930 THEN
            exp_f := 0;
        ELSIF x =- 22929 THEN
            exp_f := 0;
        ELSIF x =- 22928 THEN
            exp_f := 0;
        ELSIF x =- 22927 THEN
            exp_f := 0;
        ELSIF x =- 22926 THEN
            exp_f := 0;
        ELSIF x =- 22925 THEN
            exp_f := 0;
        ELSIF x =- 22924 THEN
            exp_f := 0;
        ELSIF x =- 22923 THEN
            exp_f := 0;
        ELSIF x =- 22922 THEN
            exp_f := 0;
        ELSIF x =- 22921 THEN
            exp_f := 0;
        ELSIF x =- 22920 THEN
            exp_f := 0;
        ELSIF x =- 22919 THEN
            exp_f := 0;
        ELSIF x =- 22918 THEN
            exp_f := 0;
        ELSIF x =- 22917 THEN
            exp_f := 0;
        ELSIF x =- 22916 THEN
            exp_f := 0;
        ELSIF x =- 22915 THEN
            exp_f := 0;
        ELSIF x =- 22914 THEN
            exp_f := 0;
        ELSIF x =- 22913 THEN
            exp_f := 0;
        ELSIF x =- 22912 THEN
            exp_f := 0;
        ELSIF x =- 22911 THEN
            exp_f := 0;
        ELSIF x =- 22910 THEN
            exp_f := 0;
        ELSIF x =- 22909 THEN
            exp_f := 0;
        ELSIF x =- 22908 THEN
            exp_f := 0;
        ELSIF x =- 22907 THEN
            exp_f := 0;
        ELSIF x =- 22906 THEN
            exp_f := 0;
        ELSIF x =- 22905 THEN
            exp_f := 0;
        ELSIF x =- 22904 THEN
            exp_f := 0;
        ELSIF x =- 22903 THEN
            exp_f := 0;
        ELSIF x =- 22902 THEN
            exp_f := 0;
        ELSIF x =- 22901 THEN
            exp_f := 0;
        ELSIF x =- 22900 THEN
            exp_f := 0;
        ELSIF x =- 22899 THEN
            exp_f := 0;
        ELSIF x =- 22898 THEN
            exp_f := 0;
        ELSIF x =- 22897 THEN
            exp_f := 0;
        ELSIF x =- 22896 THEN
            exp_f := 0;
        ELSIF x =- 22895 THEN
            exp_f := 0;
        ELSIF x =- 22894 THEN
            exp_f := 0;
        ELSIF x =- 22893 THEN
            exp_f := 0;
        ELSIF x =- 22892 THEN
            exp_f := 0;
        ELSIF x =- 22891 THEN
            exp_f := 0;
        ELSIF x =- 22890 THEN
            exp_f := 0;
        ELSIF x =- 22889 THEN
            exp_f := 0;
        ELSIF x =- 22888 THEN
            exp_f := 0;
        ELSIF x =- 22887 THEN
            exp_f := 0;
        ELSIF x =- 22886 THEN
            exp_f := 0;
        ELSIF x =- 22885 THEN
            exp_f := 0;
        ELSIF x =- 22884 THEN
            exp_f := 0;
        ELSIF x =- 22883 THEN
            exp_f := 0;
        ELSIF x =- 22882 THEN
            exp_f := 0;
        ELSIF x =- 22881 THEN
            exp_f := 0;
        ELSIF x =- 22880 THEN
            exp_f := 0;
        ELSIF x =- 22879 THEN
            exp_f := 0;
        ELSIF x =- 22878 THEN
            exp_f := 0;
        ELSIF x =- 22877 THEN
            exp_f := 0;
        ELSIF x =- 22876 THEN
            exp_f := 0;
        ELSIF x =- 22875 THEN
            exp_f := 0;
        ELSIF x =- 22874 THEN
            exp_f := 0;
        ELSIF x =- 22873 THEN
            exp_f := 0;
        ELSIF x =- 22872 THEN
            exp_f := 0;
        ELSIF x =- 22871 THEN
            exp_f := 0;
        ELSIF x =- 22870 THEN
            exp_f := 0;
        ELSIF x =- 22869 THEN
            exp_f := 0;
        ELSIF x =- 22868 THEN
            exp_f := 0;
        ELSIF x =- 22867 THEN
            exp_f := 0;
        ELSIF x =- 22866 THEN
            exp_f := 0;
        ELSIF x =- 22865 THEN
            exp_f := 0;
        ELSIF x =- 22864 THEN
            exp_f := 0;
        ELSIF x =- 22863 THEN
            exp_f := 0;
        ELSIF x =- 22862 THEN
            exp_f := 0;
        ELSIF x =- 22861 THEN
            exp_f := 0;
        ELSIF x =- 22860 THEN
            exp_f := 0;
        ELSIF x =- 22859 THEN
            exp_f := 0;
        ELSIF x =- 22858 THEN
            exp_f := 0;
        ELSIF x =- 22857 THEN
            exp_f := 0;
        ELSIF x =- 22856 THEN
            exp_f := 0;
        ELSIF x =- 22855 THEN
            exp_f := 0;
        ELSIF x =- 22854 THEN
            exp_f := 0;
        ELSIF x =- 22853 THEN
            exp_f := 0;
        ELSIF x =- 22852 THEN
            exp_f := 0;
        ELSIF x =- 22851 THEN
            exp_f := 0;
        ELSIF x =- 22850 THEN
            exp_f := 0;
        ELSIF x =- 22849 THEN
            exp_f := 0;
        ELSIF x =- 22848 THEN
            exp_f := 0;
        ELSIF x =- 22847 THEN
            exp_f := 0;
        ELSIF x =- 22846 THEN
            exp_f := 0;
        ELSIF x =- 22845 THEN
            exp_f := 0;
        ELSIF x =- 22844 THEN
            exp_f := 0;
        ELSIF x =- 22843 THEN
            exp_f := 0;
        ELSIF x =- 22842 THEN
            exp_f := 0;
        ELSIF x =- 22841 THEN
            exp_f := 0;
        ELSIF x =- 22840 THEN
            exp_f := 0;
        ELSIF x =- 22839 THEN
            exp_f := 0;
        ELSIF x =- 22838 THEN
            exp_f := 0;
        ELSIF x =- 22837 THEN
            exp_f := 0;
        ELSIF x =- 22836 THEN
            exp_f := 0;
        ELSIF x =- 22835 THEN
            exp_f := 0;
        ELSIF x =- 22834 THEN
            exp_f := 0;
        ELSIF x =- 22833 THEN
            exp_f := 0;
        ELSIF x =- 22832 THEN
            exp_f := 0;
        ELSIF x =- 22831 THEN
            exp_f := 0;
        ELSIF x =- 22830 THEN
            exp_f := 0;
        ELSIF x =- 22829 THEN
            exp_f := 0;
        ELSIF x =- 22828 THEN
            exp_f := 0;
        ELSIF x =- 22827 THEN
            exp_f := 0;
        ELSIF x =- 22826 THEN
            exp_f := 0;
        ELSIF x =- 22825 THEN
            exp_f := 0;
        ELSIF x =- 22824 THEN
            exp_f := 0;
        ELSIF x =- 22823 THEN
            exp_f := 0;
        ELSIF x =- 22822 THEN
            exp_f := 0;
        ELSIF x =- 22821 THEN
            exp_f := 0;
        ELSIF x =- 22820 THEN
            exp_f := 0;
        ELSIF x =- 22819 THEN
            exp_f := 0;
        ELSIF x =- 22818 THEN
            exp_f := 0;
        ELSIF x =- 22817 THEN
            exp_f := 0;
        ELSIF x =- 22816 THEN
            exp_f := 0;
        ELSIF x =- 22815 THEN
            exp_f := 0;
        ELSIF x =- 22814 THEN
            exp_f := 0;
        ELSIF x =- 22813 THEN
            exp_f := 0;
        ELSIF x =- 22812 THEN
            exp_f := 0;
        ELSIF x =- 22811 THEN
            exp_f := 0;
        ELSIF x =- 22810 THEN
            exp_f := 0;
        ELSIF x =- 22809 THEN
            exp_f := 0;
        ELSIF x =- 22808 THEN
            exp_f := 0;
        ELSIF x =- 22807 THEN
            exp_f := 0;
        ELSIF x =- 22806 THEN
            exp_f := 0;
        ELSIF x =- 22805 THEN
            exp_f := 0;
        ELSIF x =- 22804 THEN
            exp_f := 0;
        ELSIF x =- 22803 THEN
            exp_f := 0;
        ELSIF x =- 22802 THEN
            exp_f := 0;
        ELSIF x =- 22801 THEN
            exp_f := 0;
        ELSIF x =- 22800 THEN
            exp_f := 0;
        ELSIF x =- 22799 THEN
            exp_f := 0;
        ELSIF x =- 22798 THEN
            exp_f := 0;
        ELSIF x =- 22797 THEN
            exp_f := 0;
        ELSIF x =- 22796 THEN
            exp_f := 0;
        ELSIF x =- 22795 THEN
            exp_f := 0;
        ELSIF x =- 22794 THEN
            exp_f := 0;
        ELSIF x =- 22793 THEN
            exp_f := 0;
        ELSIF x =- 22792 THEN
            exp_f := 0;
        ELSIF x =- 22791 THEN
            exp_f := 0;
        ELSIF x =- 22790 THEN
            exp_f := 0;
        ELSIF x =- 22789 THEN
            exp_f := 0;
        ELSIF x =- 22788 THEN
            exp_f := 0;
        ELSIF x =- 22787 THEN
            exp_f := 0;
        ELSIF x =- 22786 THEN
            exp_f := 0;
        ELSIF x =- 22785 THEN
            exp_f := 0;
        ELSIF x =- 22784 THEN
            exp_f := 0;
        ELSIF x =- 22783 THEN
            exp_f := 0;
        ELSIF x =- 22782 THEN
            exp_f := 0;
        ELSIF x =- 22781 THEN
            exp_f := 0;
        ELSIF x =- 22780 THEN
            exp_f := 0;
        ELSIF x =- 22779 THEN
            exp_f := 0;
        ELSIF x =- 22778 THEN
            exp_f := 0;
        ELSIF x =- 22777 THEN
            exp_f := 0;
        ELSIF x =- 22776 THEN
            exp_f := 0;
        ELSIF x =- 22775 THEN
            exp_f := 0;
        ELSIF x =- 22774 THEN
            exp_f := 0;
        ELSIF x =- 22773 THEN
            exp_f := 0;
        ELSIF x =- 22772 THEN
            exp_f := 0;
        ELSIF x =- 22771 THEN
            exp_f := 0;
        ELSIF x =- 22770 THEN
            exp_f := 0;
        ELSIF x =- 22769 THEN
            exp_f := 0;
        ELSIF x =- 22768 THEN
            exp_f := 0;
        ELSIF x =- 22767 THEN
            exp_f := 0;
        ELSIF x =- 22766 THEN
            exp_f := 0;
        ELSIF x =- 22765 THEN
            exp_f := 0;
        ELSIF x =- 22764 THEN
            exp_f := 0;
        ELSIF x =- 22763 THEN
            exp_f := 0;
        ELSIF x =- 22762 THEN
            exp_f := 0;
        ELSIF x =- 22761 THEN
            exp_f := 0;
        ELSIF x =- 22760 THEN
            exp_f := 0;
        ELSIF x =- 22759 THEN
            exp_f := 0;
        ELSIF x =- 22758 THEN
            exp_f := 0;
        ELSIF x =- 22757 THEN
            exp_f := 0;
        ELSIF x =- 22756 THEN
            exp_f := 0;
        ELSIF x =- 22755 THEN
            exp_f := 0;
        ELSIF x =- 22754 THEN
            exp_f := 0;
        ELSIF x =- 22753 THEN
            exp_f := 0;
        ELSIF x =- 22752 THEN
            exp_f := 0;
        ELSIF x =- 22751 THEN
            exp_f := 0;
        ELSIF x =- 22750 THEN
            exp_f := 0;
        ELSIF x =- 22749 THEN
            exp_f := 0;
        ELSIF x =- 22748 THEN
            exp_f := 0;
        ELSIF x =- 22747 THEN
            exp_f := 0;
        ELSIF x =- 22746 THEN
            exp_f := 0;
        ELSIF x =- 22745 THEN
            exp_f := 0;
        ELSIF x =- 22744 THEN
            exp_f := 0;
        ELSIF x =- 22743 THEN
            exp_f := 0;
        ELSIF x =- 22742 THEN
            exp_f := 0;
        ELSIF x =- 22741 THEN
            exp_f := 0;
        ELSIF x =- 22740 THEN
            exp_f := 0;
        ELSIF x =- 22739 THEN
            exp_f := 0;
        ELSIF x =- 22738 THEN
            exp_f := 0;
        ELSIF x =- 22737 THEN
            exp_f := 0;
        ELSIF x =- 22736 THEN
            exp_f := 0;
        ELSIF x =- 22735 THEN
            exp_f := 0;
        ELSIF x =- 22734 THEN
            exp_f := 0;
        ELSIF x =- 22733 THEN
            exp_f := 0;
        ELSIF x =- 22732 THEN
            exp_f := 0;
        ELSIF x =- 22731 THEN
            exp_f := 0;
        ELSIF x =- 22730 THEN
            exp_f := 0;
        ELSIF x =- 22729 THEN
            exp_f := 0;
        ELSIF x =- 22728 THEN
            exp_f := 0;
        ELSIF x =- 22727 THEN
            exp_f := 0;
        ELSIF x =- 22726 THEN
            exp_f := 0;
        ELSIF x =- 22725 THEN
            exp_f := 0;
        ELSIF x =- 22724 THEN
            exp_f := 0;
        ELSIF x =- 22723 THEN
            exp_f := 0;
        ELSIF x =- 22722 THEN
            exp_f := 0;
        ELSIF x =- 22721 THEN
            exp_f := 0;
        ELSIF x =- 22720 THEN
            exp_f := 0;
        ELSIF x =- 22719 THEN
            exp_f := 0;
        ELSIF x =- 22718 THEN
            exp_f := 0;
        ELSIF x =- 22717 THEN
            exp_f := 0;
        ELSIF x =- 22716 THEN
            exp_f := 0;
        ELSIF x =- 22715 THEN
            exp_f := 0;
        ELSIF x =- 22714 THEN
            exp_f := 0;
        ELSIF x =- 22713 THEN
            exp_f := 0;
        ELSIF x =- 22712 THEN
            exp_f := 0;
        ELSIF x =- 22711 THEN
            exp_f := 0;
        ELSIF x =- 22710 THEN
            exp_f := 0;
        ELSIF x =- 22709 THEN
            exp_f := 0;
        ELSIF x =- 22708 THEN
            exp_f := 0;
        ELSIF x =- 22707 THEN
            exp_f := 0;
        ELSIF x =- 22706 THEN
            exp_f := 0;
        ELSIF x =- 22705 THEN
            exp_f := 0;
        ELSIF x =- 22704 THEN
            exp_f := 0;
        ELSIF x =- 22703 THEN
            exp_f := 0;
        ELSIF x =- 22702 THEN
            exp_f := 0;
        ELSIF x =- 22701 THEN
            exp_f := 0;
        ELSIF x =- 22700 THEN
            exp_f := 0;
        ELSIF x =- 22699 THEN
            exp_f := 0;
        ELSIF x =- 22698 THEN
            exp_f := 0;
        ELSIF x =- 22697 THEN
            exp_f := 0;
        ELSIF x =- 22696 THEN
            exp_f := 0;
        ELSIF x =- 22695 THEN
            exp_f := 0;
        ELSIF x =- 22694 THEN
            exp_f := 0;
        ELSIF x =- 22693 THEN
            exp_f := 0;
        ELSIF x =- 22692 THEN
            exp_f := 0;
        ELSIF x =- 22691 THEN
            exp_f := 0;
        ELSIF x =- 22690 THEN
            exp_f := 0;
        ELSIF x =- 22689 THEN
            exp_f := 0;
        ELSIF x =- 22688 THEN
            exp_f := 0;
        ELSIF x =- 22687 THEN
            exp_f := 0;
        ELSIF x =- 22686 THEN
            exp_f := 0;
        ELSIF x =- 22685 THEN
            exp_f := 0;
        ELSIF x =- 22684 THEN
            exp_f := 0;
        ELSIF x =- 22683 THEN
            exp_f := 0;
        ELSIF x =- 22682 THEN
            exp_f := 0;
        ELSIF x =- 22681 THEN
            exp_f := 0;
        ELSIF x =- 22680 THEN
            exp_f := 0;
        ELSIF x =- 22679 THEN
            exp_f := 0;
        ELSIF x =- 22678 THEN
            exp_f := 0;
        ELSIF x =- 22677 THEN
            exp_f := 0;
        ELSIF x =- 22676 THEN
            exp_f := 0;
        ELSIF x =- 22675 THEN
            exp_f := 0;
        ELSIF x =- 22674 THEN
            exp_f := 0;
        ELSIF x =- 22673 THEN
            exp_f := 0;
        ELSIF x =- 22672 THEN
            exp_f := 0;
        ELSIF x =- 22671 THEN
            exp_f := 0;
        ELSIF x =- 22670 THEN
            exp_f := 0;
        ELSIF x =- 22669 THEN
            exp_f := 0;
        ELSIF x =- 22668 THEN
            exp_f := 0;
        ELSIF x =- 22667 THEN
            exp_f := 0;
        ELSIF x =- 22666 THEN
            exp_f := 0;
        ELSIF x =- 22665 THEN
            exp_f := 0;
        ELSIF x =- 22664 THEN
            exp_f := 0;
        ELSIF x =- 22663 THEN
            exp_f := 0;
        ELSIF x =- 22662 THEN
            exp_f := 0;
        ELSIF x =- 22661 THEN
            exp_f := 0;
        ELSIF x =- 22660 THEN
            exp_f := 0;
        ELSIF x =- 22659 THEN
            exp_f := 0;
        ELSIF x =- 22658 THEN
            exp_f := 0;
        ELSIF x =- 22657 THEN
            exp_f := 0;
        ELSIF x =- 22656 THEN
            exp_f := 0;
        ELSIF x =- 22655 THEN
            exp_f := 0;
        ELSIF x =- 22654 THEN
            exp_f := 0;
        ELSIF x =- 22653 THEN
            exp_f := 0;
        ELSIF x =- 22652 THEN
            exp_f := 0;
        ELSIF x =- 22651 THEN
            exp_f := 0;
        ELSIF x =- 22650 THEN
            exp_f := 0;
        ELSIF x =- 22649 THEN
            exp_f := 0;
        ELSIF x =- 22648 THEN
            exp_f := 0;
        ELSIF x =- 22647 THEN
            exp_f := 0;
        ELSIF x =- 22646 THEN
            exp_f := 0;
        ELSIF x =- 22645 THEN
            exp_f := 0;
        ELSIF x =- 22644 THEN
            exp_f := 0;
        ELSIF x =- 22643 THEN
            exp_f := 0;
        ELSIF x =- 22642 THEN
            exp_f := 0;
        ELSIF x =- 22641 THEN
            exp_f := 0;
        ELSIF x =- 22640 THEN
            exp_f := 0;
        ELSIF x =- 22639 THEN
            exp_f := 0;
        ELSIF x =- 22638 THEN
            exp_f := 0;
        ELSIF x =- 22637 THEN
            exp_f := 0;
        ELSIF x =- 22636 THEN
            exp_f := 0;
        ELSIF x =- 22635 THEN
            exp_f := 0;
        ELSIF x =- 22634 THEN
            exp_f := 0;
        ELSIF x =- 22633 THEN
            exp_f := 0;
        ELSIF x =- 22632 THEN
            exp_f := 0;
        ELSIF x =- 22631 THEN
            exp_f := 0;
        ELSIF x =- 22630 THEN
            exp_f := 0;
        ELSIF x =- 22629 THEN
            exp_f := 0;
        ELSIF x =- 22628 THEN
            exp_f := 0;
        ELSIF x =- 22627 THEN
            exp_f := 0;
        ELSIF x =- 22626 THEN
            exp_f := 0;
        ELSIF x =- 22625 THEN
            exp_f := 0;
        ELSIF x =- 22624 THEN
            exp_f := 0;
        ELSIF x =- 22623 THEN
            exp_f := 0;
        ELSIF x =- 22622 THEN
            exp_f := 0;
        ELSIF x =- 22621 THEN
            exp_f := 0;
        ELSIF x =- 22620 THEN
            exp_f := 0;
        ELSIF x =- 22619 THEN
            exp_f := 0;
        ELSIF x =- 22618 THEN
            exp_f := 0;
        ELSIF x =- 22617 THEN
            exp_f := 0;
        ELSIF x =- 22616 THEN
            exp_f := 0;
        ELSIF x =- 22615 THEN
            exp_f := 0;
        ELSIF x =- 22614 THEN
            exp_f := 0;
        ELSIF x =- 22613 THEN
            exp_f := 0;
        ELSIF x =- 22612 THEN
            exp_f := 0;
        ELSIF x =- 22611 THEN
            exp_f := 0;
        ELSIF x =- 22610 THEN
            exp_f := 0;
        ELSIF x =- 22609 THEN
            exp_f := 0;
        ELSIF x =- 22608 THEN
            exp_f := 0;
        ELSIF x =- 22607 THEN
            exp_f := 0;
        ELSIF x =- 22606 THEN
            exp_f := 0;
        ELSIF x =- 22605 THEN
            exp_f := 0;
        ELSIF x =- 22604 THEN
            exp_f := 0;
        ELSIF x =- 22603 THEN
            exp_f := 0;
        ELSIF x =- 22602 THEN
            exp_f := 0;
        ELSIF x =- 22601 THEN
            exp_f := 0;
        ELSIF x =- 22600 THEN
            exp_f := 0;
        ELSIF x =- 22599 THEN
            exp_f := 0;
        ELSIF x =- 22598 THEN
            exp_f := 0;
        ELSIF x =- 22597 THEN
            exp_f := 0;
        ELSIF x =- 22596 THEN
            exp_f := 0;
        ELSIF x =- 22595 THEN
            exp_f := 0;
        ELSIF x =- 22594 THEN
            exp_f := 0;
        ELSIF x =- 22593 THEN
            exp_f := 0;
        ELSIF x =- 22592 THEN
            exp_f := 0;
        ELSIF x =- 22591 THEN
            exp_f := 0;
        ELSIF x =- 22590 THEN
            exp_f := 0;
        ELSIF x =- 22589 THEN
            exp_f := 0;
        ELSIF x =- 22588 THEN
            exp_f := 0;
        ELSIF x =- 22587 THEN
            exp_f := 0;
        ELSIF x =- 22586 THEN
            exp_f := 0;
        ELSIF x =- 22585 THEN
            exp_f := 0;
        ELSIF x =- 22584 THEN
            exp_f := 0;
        ELSIF x =- 22583 THEN
            exp_f := 0;
        ELSIF x =- 22582 THEN
            exp_f := 0;
        ELSIF x =- 22581 THEN
            exp_f := 0;
        ELSIF x =- 22580 THEN
            exp_f := 0;
        ELSIF x =- 22579 THEN
            exp_f := 0;
        ELSIF x =- 22578 THEN
            exp_f := 0;
        ELSIF x =- 22577 THEN
            exp_f := 0;
        ELSIF x =- 22576 THEN
            exp_f := 0;
        ELSIF x =- 22575 THEN
            exp_f := 0;
        ELSIF x =- 22574 THEN
            exp_f := 0;
        ELSIF x =- 22573 THEN
            exp_f := 0;
        ELSIF x =- 22572 THEN
            exp_f := 0;
        ELSIF x =- 22571 THEN
            exp_f := 0;
        ELSIF x =- 22570 THEN
            exp_f := 0;
        ELSIF x =- 22569 THEN
            exp_f := 0;
        ELSIF x =- 22568 THEN
            exp_f := 0;
        ELSIF x =- 22567 THEN
            exp_f := 0;
        ELSIF x =- 22566 THEN
            exp_f := 0;
        ELSIF x =- 22565 THEN
            exp_f := 0;
        ELSIF x =- 22564 THEN
            exp_f := 0;
        ELSIF x =- 22563 THEN
            exp_f := 0;
        ELSIF x =- 22562 THEN
            exp_f := 0;
        ELSIF x =- 22561 THEN
            exp_f := 0;
        ELSIF x =- 22560 THEN
            exp_f := 0;
        ELSIF x =- 22559 THEN
            exp_f := 0;
        ELSIF x =- 22558 THEN
            exp_f := 0;
        ELSIF x =- 22557 THEN
            exp_f := 0;
        ELSIF x =- 22556 THEN
            exp_f := 0;
        ELSIF x =- 22555 THEN
            exp_f := 0;
        ELSIF x =- 22554 THEN
            exp_f := 0;
        ELSIF x =- 22553 THEN
            exp_f := 0;
        ELSIF x =- 22552 THEN
            exp_f := 0;
        ELSIF x =- 22551 THEN
            exp_f := 0;
        ELSIF x =- 22550 THEN
            exp_f := 0;
        ELSIF x =- 22549 THEN
            exp_f := 0;
        ELSIF x =- 22548 THEN
            exp_f := 0;
        ELSIF x =- 22547 THEN
            exp_f := 0;
        ELSIF x =- 22546 THEN
            exp_f := 0;
        ELSIF x =- 22545 THEN
            exp_f := 0;
        ELSIF x =- 22544 THEN
            exp_f := 0;
        ELSIF x =- 22543 THEN
            exp_f := 0;
        ELSIF x =- 22542 THEN
            exp_f := 0;
        ELSIF x =- 22541 THEN
            exp_f := 0;
        ELSIF x =- 22540 THEN
            exp_f := 0;
        ELSIF x =- 22539 THEN
            exp_f := 0;
        ELSIF x =- 22538 THEN
            exp_f := 0;
        ELSIF x =- 22537 THEN
            exp_f := 0;
        ELSIF x =- 22536 THEN
            exp_f := 0;
        ELSIF x =- 22535 THEN
            exp_f := 0;
        ELSIF x =- 22534 THEN
            exp_f := 0;
        ELSIF x =- 22533 THEN
            exp_f := 0;
        ELSIF x =- 22532 THEN
            exp_f := 0;
        ELSIF x =- 22531 THEN
            exp_f := 0;
        ELSIF x =- 22530 THEN
            exp_f := 0;
        ELSIF x =- 22529 THEN
            exp_f := 0;
        ELSIF x =- 22528 THEN
            exp_f := 0;
        ELSIF x =- 22527 THEN
            exp_f := 0;
        ELSIF x =- 22526 THEN
            exp_f := 0;
        ELSIF x =- 22525 THEN
            exp_f := 0;
        ELSIF x =- 22524 THEN
            exp_f := 0;
        ELSIF x =- 22523 THEN
            exp_f := 0;
        ELSIF x =- 22522 THEN
            exp_f := 0;
        ELSIF x =- 22521 THEN
            exp_f := 0;
        ELSIF x =- 22520 THEN
            exp_f := 0;
        ELSIF x =- 22519 THEN
            exp_f := 0;
        ELSIF x =- 22518 THEN
            exp_f := 0;
        ELSIF x =- 22517 THEN
            exp_f := 0;
        ELSIF x =- 22516 THEN
            exp_f := 0;
        ELSIF x =- 22515 THEN
            exp_f := 0;
        ELSIF x =- 22514 THEN
            exp_f := 0;
        ELSIF x =- 22513 THEN
            exp_f := 0;
        ELSIF x =- 22512 THEN
            exp_f := 0;
        ELSIF x =- 22511 THEN
            exp_f := 0;
        ELSIF x =- 22510 THEN
            exp_f := 0;
        ELSIF x =- 22509 THEN
            exp_f := 0;
        ELSIF x =- 22508 THEN
            exp_f := 0;
        ELSIF x =- 22507 THEN
            exp_f := 0;
        ELSIF x =- 22506 THEN
            exp_f := 0;
        ELSIF x =- 22505 THEN
            exp_f := 0;
        ELSIF x =- 22504 THEN
            exp_f := 0;
        ELSIF x =- 22503 THEN
            exp_f := 0;
        ELSIF x =- 22502 THEN
            exp_f := 0;
        ELSIF x =- 22501 THEN
            exp_f := 0;
        ELSIF x =- 22500 THEN
            exp_f := 0;
        ELSIF x =- 22499 THEN
            exp_f := 0;
        ELSIF x =- 22498 THEN
            exp_f := 0;
        ELSIF x =- 22497 THEN
            exp_f := 0;
        ELSIF x =- 22496 THEN
            exp_f := 0;
        ELSIF x =- 22495 THEN
            exp_f := 0;
        ELSIF x =- 22494 THEN
            exp_f := 0;
        ELSIF x =- 22493 THEN
            exp_f := 0;
        ELSIF x =- 22492 THEN
            exp_f := 0;
        ELSIF x =- 22491 THEN
            exp_f := 0;
        ELSIF x =- 22490 THEN
            exp_f := 0;
        ELSIF x =- 22489 THEN
            exp_f := 0;
        ELSIF x =- 22488 THEN
            exp_f := 0;
        ELSIF x =- 22487 THEN
            exp_f := 0;
        ELSIF x =- 22486 THEN
            exp_f := 0;
        ELSIF x =- 22485 THEN
            exp_f := 0;
        ELSIF x =- 22484 THEN
            exp_f := 0;
        ELSIF x =- 22483 THEN
            exp_f := 0;
        ELSIF x =- 22482 THEN
            exp_f := 0;
        ELSIF x =- 22481 THEN
            exp_f := 0;
        ELSIF x =- 22480 THEN
            exp_f := 0;
        ELSIF x =- 22479 THEN
            exp_f := 0;
        ELSIF x =- 22478 THEN
            exp_f := 0;
        ELSIF x =- 22477 THEN
            exp_f := 0;
        ELSIF x =- 22476 THEN
            exp_f := 0;
        ELSIF x =- 22475 THEN
            exp_f := 0;
        ELSIF x =- 22474 THEN
            exp_f := 0;
        ELSIF x =- 22473 THEN
            exp_f := 0;
        ELSIF x =- 22472 THEN
            exp_f := 0;
        ELSIF x =- 22471 THEN
            exp_f := 0;
        ELSIF x =- 22470 THEN
            exp_f := 0;
        ELSIF x =- 22469 THEN
            exp_f := 0;
        ELSIF x =- 22468 THEN
            exp_f := 0;
        ELSIF x =- 22467 THEN
            exp_f := 0;
        ELSIF x =- 22466 THEN
            exp_f := 0;
        ELSIF x =- 22465 THEN
            exp_f := 0;
        ELSIF x =- 22464 THEN
            exp_f := 0;
        ELSIF x =- 22463 THEN
            exp_f := 0;
        ELSIF x =- 22462 THEN
            exp_f := 0;
        ELSIF x =- 22461 THEN
            exp_f := 0;
        ELSIF x =- 22460 THEN
            exp_f := 0;
        ELSIF x =- 22459 THEN
            exp_f := 0;
        ELSIF x =- 22458 THEN
            exp_f := 0;
        ELSIF x =- 22457 THEN
            exp_f := 0;
        ELSIF x =- 22456 THEN
            exp_f := 0;
        ELSIF x =- 22455 THEN
            exp_f := 0;
        ELSIF x =- 22454 THEN
            exp_f := 0;
        ELSIF x =- 22453 THEN
            exp_f := 0;
        ELSIF x =- 22452 THEN
            exp_f := 0;
        ELSIF x =- 22451 THEN
            exp_f := 0;
        ELSIF x =- 22450 THEN
            exp_f := 0;
        ELSIF x =- 22449 THEN
            exp_f := 0;
        ELSIF x =- 22448 THEN
            exp_f := 0;
        ELSIF x =- 22447 THEN
            exp_f := 0;
        ELSIF x =- 22446 THEN
            exp_f := 0;
        ELSIF x =- 22445 THEN
            exp_f := 0;
        ELSIF x =- 22444 THEN
            exp_f := 0;
        ELSIF x =- 22443 THEN
            exp_f := 0;
        ELSIF x =- 22442 THEN
            exp_f := 0;
        ELSIF x =- 22441 THEN
            exp_f := 0;
        ELSIF x =- 22440 THEN
            exp_f := 0;
        ELSIF x =- 22439 THEN
            exp_f := 0;
        ELSIF x =- 22438 THEN
            exp_f := 0;
        ELSIF x =- 22437 THEN
            exp_f := 0;
        ELSIF x =- 22436 THEN
            exp_f := 0;
        ELSIF x =- 22435 THEN
            exp_f := 0;
        ELSIF x =- 22434 THEN
            exp_f := 0;
        ELSIF x =- 22433 THEN
            exp_f := 0;
        ELSIF x =- 22432 THEN
            exp_f := 0;
        ELSIF x =- 22431 THEN
            exp_f := 0;
        ELSIF x =- 22430 THEN
            exp_f := 0;
        ELSIF x =- 22429 THEN
            exp_f := 0;
        ELSIF x =- 22428 THEN
            exp_f := 0;
        ELSIF x =- 22427 THEN
            exp_f := 0;
        ELSIF x =- 22426 THEN
            exp_f := 0;
        ELSIF x =- 22425 THEN
            exp_f := 0;
        ELSIF x =- 22424 THEN
            exp_f := 0;
        ELSIF x =- 22423 THEN
            exp_f := 0;
        ELSIF x =- 22422 THEN
            exp_f := 0;
        ELSIF x =- 22421 THEN
            exp_f := 0;
        ELSIF x =- 22420 THEN
            exp_f := 0;
        ELSIF x =- 22419 THEN
            exp_f := 0;
        ELSIF x =- 22418 THEN
            exp_f := 0;
        ELSIF x =- 22417 THEN
            exp_f := 0;
        ELSIF x =- 22416 THEN
            exp_f := 0;
        ELSIF x =- 22415 THEN
            exp_f := 0;
        ELSIF x =- 22414 THEN
            exp_f := 0;
        ELSIF x =- 22413 THEN
            exp_f := 0;
        ELSIF x =- 22412 THEN
            exp_f := 0;
        ELSIF x =- 22411 THEN
            exp_f := 0;
        ELSIF x =- 22410 THEN
            exp_f := 0;
        ELSIF x =- 22409 THEN
            exp_f := 0;
        ELSIF x =- 22408 THEN
            exp_f := 0;
        ELSIF x =- 22407 THEN
            exp_f := 0;
        ELSIF x =- 22406 THEN
            exp_f := 0;
        ELSIF x =- 22405 THEN
            exp_f := 0;
        ELSIF x =- 22404 THEN
            exp_f := 0;
        ELSIF x =- 22403 THEN
            exp_f := 0;
        ELSIF x =- 22402 THEN
            exp_f := 0;
        ELSIF x =- 22401 THEN
            exp_f := 0;
        ELSIF x =- 22400 THEN
            exp_f := 0;
        ELSIF x =- 22399 THEN
            exp_f := 0;
        ELSIF x =- 22398 THEN
            exp_f := 0;
        ELSIF x =- 22397 THEN
            exp_f := 0;
        ELSIF x =- 22396 THEN
            exp_f := 0;
        ELSIF x =- 22395 THEN
            exp_f := 0;
        ELSIF x =- 22394 THEN
            exp_f := 0;
        ELSIF x =- 22393 THEN
            exp_f := 0;
        ELSIF x =- 22392 THEN
            exp_f := 0;
        ELSIF x =- 22391 THEN
            exp_f := 0;
        ELSIF x =- 22390 THEN
            exp_f := 0;
        ELSIF x =- 22389 THEN
            exp_f := 0;
        ELSIF x =- 22388 THEN
            exp_f := 0;
        ELSIF x =- 22387 THEN
            exp_f := 0;
        ELSIF x =- 22386 THEN
            exp_f := 0;
        ELSIF x =- 22385 THEN
            exp_f := 0;
        ELSIF x =- 22384 THEN
            exp_f := 0;
        ELSIF x =- 22383 THEN
            exp_f := 0;
        ELSIF x =- 22382 THEN
            exp_f := 0;
        ELSIF x =- 22381 THEN
            exp_f := 0;
        ELSIF x =- 22380 THEN
            exp_f := 0;
        ELSIF x =- 22379 THEN
            exp_f := 0;
        ELSIF x =- 22378 THEN
            exp_f := 0;
        ELSIF x =- 22377 THEN
            exp_f := 0;
        ELSIF x =- 22376 THEN
            exp_f := 0;
        ELSIF x =- 22375 THEN
            exp_f := 0;
        ELSIF x =- 22374 THEN
            exp_f := 0;
        ELSIF x =- 22373 THEN
            exp_f := 0;
        ELSIF x =- 22372 THEN
            exp_f := 0;
        ELSIF x =- 22371 THEN
            exp_f := 0;
        ELSIF x =- 22370 THEN
            exp_f := 0;
        ELSIF x =- 22369 THEN
            exp_f := 0;
        ELSIF x =- 22368 THEN
            exp_f := 0;
        ELSIF x =- 22367 THEN
            exp_f := 0;
        ELSIF x =- 22366 THEN
            exp_f := 0;
        ELSIF x =- 22365 THEN
            exp_f := 0;
        ELSIF x =- 22364 THEN
            exp_f := 0;
        ELSIF x =- 22363 THEN
            exp_f := 0;
        ELSIF x =- 22362 THEN
            exp_f := 0;
        ELSIF x =- 22361 THEN
            exp_f := 0;
        ELSIF x =- 22360 THEN
            exp_f := 0;
        ELSIF x =- 22359 THEN
            exp_f := 0;
        ELSIF x =- 22358 THEN
            exp_f := 0;
        ELSIF x =- 22357 THEN
            exp_f := 0;
        ELSIF x =- 22356 THEN
            exp_f := 0;
        ELSIF x =- 22355 THEN
            exp_f := 0;
        ELSIF x =- 22354 THEN
            exp_f := 0;
        ELSIF x =- 22353 THEN
            exp_f := 0;
        ELSIF x =- 22352 THEN
            exp_f := 0;
        ELSIF x =- 22351 THEN
            exp_f := 0;
        ELSIF x =- 22350 THEN
            exp_f := 0;
        ELSIF x =- 22349 THEN
            exp_f := 0;
        ELSIF x =- 22348 THEN
            exp_f := 0;
        ELSIF x =- 22347 THEN
            exp_f := 0;
        ELSIF x =- 22346 THEN
            exp_f := 0;
        ELSIF x =- 22345 THEN
            exp_f := 0;
        ELSIF x =- 22344 THEN
            exp_f := 0;
        ELSIF x =- 22343 THEN
            exp_f := 0;
        ELSIF x =- 22342 THEN
            exp_f := 0;
        ELSIF x =- 22341 THEN
            exp_f := 0;
        ELSIF x =- 22340 THEN
            exp_f := 0;
        ELSIF x =- 22339 THEN
            exp_f := 0;
        ELSIF x =- 22338 THEN
            exp_f := 0;
        ELSIF x =- 22337 THEN
            exp_f := 0;
        ELSIF x =- 22336 THEN
            exp_f := 0;
        ELSIF x =- 22335 THEN
            exp_f := 0;
        ELSIF x =- 22334 THEN
            exp_f := 0;
        ELSIF x =- 22333 THEN
            exp_f := 0;
        ELSIF x =- 22332 THEN
            exp_f := 0;
        ELSIF x =- 22331 THEN
            exp_f := 0;
        ELSIF x =- 22330 THEN
            exp_f := 0;
        ELSIF x =- 22329 THEN
            exp_f := 0;
        ELSIF x =- 22328 THEN
            exp_f := 0;
        ELSIF x =- 22327 THEN
            exp_f := 0;
        ELSIF x =- 22326 THEN
            exp_f := 0;
        ELSIF x =- 22325 THEN
            exp_f := 0;
        ELSIF x =- 22324 THEN
            exp_f := 0;
        ELSIF x =- 22323 THEN
            exp_f := 0;
        ELSIF x =- 22322 THEN
            exp_f := 0;
        ELSIF x =- 22321 THEN
            exp_f := 0;
        ELSIF x =- 22320 THEN
            exp_f := 0;
        ELSIF x =- 22319 THEN
            exp_f := 0;
        ELSIF x =- 22318 THEN
            exp_f := 0;
        ELSIF x =- 22317 THEN
            exp_f := 0;
        ELSIF x =- 22316 THEN
            exp_f := 0;
        ELSIF x =- 22315 THEN
            exp_f := 0;
        ELSIF x =- 22314 THEN
            exp_f := 0;
        ELSIF x =- 22313 THEN
            exp_f := 0;
        ELSIF x =- 22312 THEN
            exp_f := 0;
        ELSIF x =- 22311 THEN
            exp_f := 0;
        ELSIF x =- 22310 THEN
            exp_f := 0;
        ELSIF x =- 22309 THEN
            exp_f := 0;
        ELSIF x =- 22308 THEN
            exp_f := 0;
        ELSIF x =- 22307 THEN
            exp_f := 0;
        ELSIF x =- 22306 THEN
            exp_f := 0;
        ELSIF x =- 22305 THEN
            exp_f := 0;
        ELSIF x =- 22304 THEN
            exp_f := 0;
        ELSIF x =- 22303 THEN
            exp_f := 0;
        ELSIF x =- 22302 THEN
            exp_f := 0;
        ELSIF x =- 22301 THEN
            exp_f := 0;
        ELSIF x =- 22300 THEN
            exp_f := 0;
        ELSIF x =- 22299 THEN
            exp_f := 0;
        ELSIF x =- 22298 THEN
            exp_f := 0;
        ELSIF x =- 22297 THEN
            exp_f := 0;
        ELSIF x =- 22296 THEN
            exp_f := 0;
        ELSIF x =- 22295 THEN
            exp_f := 0;
        ELSIF x =- 22294 THEN
            exp_f := 0;
        ELSIF x =- 22293 THEN
            exp_f := 0;
        ELSIF x =- 22292 THEN
            exp_f := 0;
        ELSIF x =- 22291 THEN
            exp_f := 0;
        ELSIF x =- 22290 THEN
            exp_f := 0;
        ELSIF x =- 22289 THEN
            exp_f := 0;
        ELSIF x =- 22288 THEN
            exp_f := 0;
        ELSIF x =- 22287 THEN
            exp_f := 0;
        ELSIF x =- 22286 THEN
            exp_f := 0;
        ELSIF x =- 22285 THEN
            exp_f := 0;
        ELSIF x =- 22284 THEN
            exp_f := 0;
        ELSIF x =- 22283 THEN
            exp_f := 0;
        ELSIF x =- 22282 THEN
            exp_f := 0;
        ELSIF x =- 22281 THEN
            exp_f := 0;
        ELSIF x =- 22280 THEN
            exp_f := 0;
        ELSIF x =- 22279 THEN
            exp_f := 0;
        ELSIF x =- 22278 THEN
            exp_f := 0;
        ELSIF x =- 22277 THEN
            exp_f := 0;
        ELSIF x =- 22276 THEN
            exp_f := 0;
        ELSIF x =- 22275 THEN
            exp_f := 0;
        ELSIF x =- 22274 THEN
            exp_f := 0;
        ELSIF x =- 22273 THEN
            exp_f := 0;
        ELSIF x =- 22272 THEN
            exp_f := 0;
        ELSIF x =- 22271 THEN
            exp_f := 0;
        ELSIF x =- 22270 THEN
            exp_f := 0;
        ELSIF x =- 22269 THEN
            exp_f := 0;
        ELSIF x =- 22268 THEN
            exp_f := 0;
        ELSIF x =- 22267 THEN
            exp_f := 0;
        ELSIF x =- 22266 THEN
            exp_f := 0;
        ELSIF x =- 22265 THEN
            exp_f := 0;
        ELSIF x =- 22264 THEN
            exp_f := 0;
        ELSIF x =- 22263 THEN
            exp_f := 0;
        ELSIF x =- 22262 THEN
            exp_f := 0;
        ELSIF x =- 22261 THEN
            exp_f := 0;
        ELSIF x =- 22260 THEN
            exp_f := 0;
        ELSIF x =- 22259 THEN
            exp_f := 0;
        ELSIF x =- 22258 THEN
            exp_f := 0;
        ELSIF x =- 22257 THEN
            exp_f := 0;
        ELSIF x =- 22256 THEN
            exp_f := 0;
        ELSIF x =- 22255 THEN
            exp_f := 0;
        ELSIF x =- 22254 THEN
            exp_f := 0;
        ELSIF x =- 22253 THEN
            exp_f := 0;
        ELSIF x =- 22252 THEN
            exp_f := 0;
        ELSIF x =- 22251 THEN
            exp_f := 0;
        ELSIF x =- 22250 THEN
            exp_f := 0;
        ELSIF x =- 22249 THEN
            exp_f := 0;
        ELSIF x =- 22248 THEN
            exp_f := 0;
        ELSIF x =- 22247 THEN
            exp_f := 0;
        ELSIF x =- 22246 THEN
            exp_f := 0;
        ELSIF x =- 22245 THEN
            exp_f := 0;
        ELSIF x =- 22244 THEN
            exp_f := 0;
        ELSIF x =- 22243 THEN
            exp_f := 0;
        ELSIF x =- 22242 THEN
            exp_f := 0;
        ELSIF x =- 22241 THEN
            exp_f := 0;
        ELSIF x =- 22240 THEN
            exp_f := 0;
        ELSIF x =- 22239 THEN
            exp_f := 0;
        ELSIF x =- 22238 THEN
            exp_f := 0;
        ELSIF x =- 22237 THEN
            exp_f := 0;
        ELSIF x =- 22236 THEN
            exp_f := 0;
        ELSIF x =- 22235 THEN
            exp_f := 0;
        ELSIF x =- 22234 THEN
            exp_f := 0;
        ELSIF x =- 22233 THEN
            exp_f := 0;
        ELSIF x =- 22232 THEN
            exp_f := 0;
        ELSIF x =- 22231 THEN
            exp_f := 0;
        ELSIF x =- 22230 THEN
            exp_f := 0;
        ELSIF x =- 22229 THEN
            exp_f := 0;
        ELSIF x =- 22228 THEN
            exp_f := 0;
        ELSIF x =- 22227 THEN
            exp_f := 0;
        ELSIF x =- 22226 THEN
            exp_f := 0;
        ELSIF x =- 22225 THEN
            exp_f := 0;
        ELSIF x =- 22224 THEN
            exp_f := 0;
        ELSIF x =- 22223 THEN
            exp_f := 0;
        ELSIF x =- 22222 THEN
            exp_f := 0;
        ELSIF x =- 22221 THEN
            exp_f := 0;
        ELSIF x =- 22220 THEN
            exp_f := 0;
        ELSIF x =- 22219 THEN
            exp_f := 0;
        ELSIF x =- 22218 THEN
            exp_f := 0;
        ELSIF x =- 22217 THEN
            exp_f := 0;
        ELSIF x =- 22216 THEN
            exp_f := 0;
        ELSIF x =- 22215 THEN
            exp_f := 0;
        ELSIF x =- 22214 THEN
            exp_f := 0;
        ELSIF x =- 22213 THEN
            exp_f := 0;
        ELSIF x =- 22212 THEN
            exp_f := 0;
        ELSIF x =- 22211 THEN
            exp_f := 0;
        ELSIF x =- 22210 THEN
            exp_f := 0;
        ELSIF x =- 22209 THEN
            exp_f := 0;
        ELSIF x =- 22208 THEN
            exp_f := 0;
        ELSIF x =- 22207 THEN
            exp_f := 0;
        ELSIF x =- 22206 THEN
            exp_f := 0;
        ELSIF x =- 22205 THEN
            exp_f := 0;
        ELSIF x =- 22204 THEN
            exp_f := 0;
        ELSIF x =- 22203 THEN
            exp_f := 0;
        ELSIF x =- 22202 THEN
            exp_f := 0;
        ELSIF x =- 22201 THEN
            exp_f := 0;
        ELSIF x =- 22200 THEN
            exp_f := 0;
        ELSIF x =- 22199 THEN
            exp_f := 0;
        ELSIF x =- 22198 THEN
            exp_f := 0;
        ELSIF x =- 22197 THEN
            exp_f := 0;
        ELSIF x =- 22196 THEN
            exp_f := 0;
        ELSIF x =- 22195 THEN
            exp_f := 0;
        ELSIF x =- 22194 THEN
            exp_f := 0;
        ELSIF x =- 22193 THEN
            exp_f := 0;
        ELSIF x =- 22192 THEN
            exp_f := 0;
        ELSIF x =- 22191 THEN
            exp_f := 0;
        ELSIF x =- 22190 THEN
            exp_f := 0;
        ELSIF x =- 22189 THEN
            exp_f := 0;
        ELSIF x =- 22188 THEN
            exp_f := 0;
        ELSIF x =- 22187 THEN
            exp_f := 0;
        ELSIF x =- 22186 THEN
            exp_f := 0;
        ELSIF x =- 22185 THEN
            exp_f := 0;
        ELSIF x =- 22184 THEN
            exp_f := 0;
        ELSIF x =- 22183 THEN
            exp_f := 0;
        ELSIF x =- 22182 THEN
            exp_f := 0;
        ELSIF x =- 22181 THEN
            exp_f := 0;
        ELSIF x =- 22180 THEN
            exp_f := 0;
        ELSIF x =- 22179 THEN
            exp_f := 0;
        ELSIF x =- 22178 THEN
            exp_f := 0;
        ELSIF x =- 22177 THEN
            exp_f := 0;
        ELSIF x =- 22176 THEN
            exp_f := 0;
        ELSIF x =- 22175 THEN
            exp_f := 0;
        ELSIF x =- 22174 THEN
            exp_f := 0;
        ELSIF x =- 22173 THEN
            exp_f := 0;
        ELSIF x =- 22172 THEN
            exp_f := 0;
        ELSIF x =- 22171 THEN
            exp_f := 0;
        ELSIF x =- 22170 THEN
            exp_f := 0;
        ELSIF x =- 22169 THEN
            exp_f := 0;
        ELSIF x =- 22168 THEN
            exp_f := 0;
        ELSIF x =- 22167 THEN
            exp_f := 0;
        ELSIF x =- 22166 THEN
            exp_f := 0;
        ELSIF x =- 22165 THEN
            exp_f := 0;
        ELSIF x =- 22164 THEN
            exp_f := 0;
        ELSIF x =- 22163 THEN
            exp_f := 0;
        ELSIF x =- 22162 THEN
            exp_f := 0;
        ELSIF x =- 22161 THEN
            exp_f := 0;
        ELSIF x =- 22160 THEN
            exp_f := 0;
        ELSIF x =- 22159 THEN
            exp_f := 0;
        ELSIF x =- 22158 THEN
            exp_f := 0;
        ELSIF x =- 22157 THEN
            exp_f := 0;
        ELSIF x =- 22156 THEN
            exp_f := 0;
        ELSIF x =- 22155 THEN
            exp_f := 0;
        ELSIF x =- 22154 THEN
            exp_f := 0;
        ELSIF x =- 22153 THEN
            exp_f := 0;
        ELSIF x =- 22152 THEN
            exp_f := 0;
        ELSIF x =- 22151 THEN
            exp_f := 0;
        ELSIF x =- 22150 THEN
            exp_f := 0;
        ELSIF x =- 22149 THEN
            exp_f := 0;
        ELSIF x =- 22148 THEN
            exp_f := 0;
        ELSIF x =- 22147 THEN
            exp_f := 0;
        ELSIF x =- 22146 THEN
            exp_f := 0;
        ELSIF x =- 22145 THEN
            exp_f := 0;
        ELSIF x =- 22144 THEN
            exp_f := 0;
        ELSIF x =- 22143 THEN
            exp_f := 0;
        ELSIF x =- 22142 THEN
            exp_f := 0;
        ELSIF x =- 22141 THEN
            exp_f := 0;
        ELSIF x =- 22140 THEN
            exp_f := 0;
        ELSIF x =- 22139 THEN
            exp_f := 0;
        ELSIF x =- 22138 THEN
            exp_f := 0;
        ELSIF x =- 22137 THEN
            exp_f := 0;
        ELSIF x =- 22136 THEN
            exp_f := 0;
        ELSIF x =- 22135 THEN
            exp_f := 0;
        ELSIF x =- 22134 THEN
            exp_f := 0;
        ELSIF x =- 22133 THEN
            exp_f := 0;
        ELSIF x =- 22132 THEN
            exp_f := 0;
        ELSIF x =- 22131 THEN
            exp_f := 0;
        ELSIF x =- 22130 THEN
            exp_f := 0;
        ELSIF x =- 22129 THEN
            exp_f := 0;
        ELSIF x =- 22128 THEN
            exp_f := 0;
        ELSIF x =- 22127 THEN
            exp_f := 0;
        ELSIF x =- 22126 THEN
            exp_f := 0;
        ELSIF x =- 22125 THEN
            exp_f := 0;
        ELSIF x =- 22124 THEN
            exp_f := 0;
        ELSIF x =- 22123 THEN
            exp_f := 0;
        ELSIF x =- 22122 THEN
            exp_f := 0;
        ELSIF x =- 22121 THEN
            exp_f := 0;
        ELSIF x =- 22120 THEN
            exp_f := 0;
        ELSIF x =- 22119 THEN
            exp_f := 0;
        ELSIF x =- 22118 THEN
            exp_f := 0;
        ELSIF x =- 22117 THEN
            exp_f := 0;
        ELSIF x =- 22116 THEN
            exp_f := 0;
        ELSIF x =- 22115 THEN
            exp_f := 0;
        ELSIF x =- 22114 THEN
            exp_f := 0;
        ELSIF x =- 22113 THEN
            exp_f := 0;
        ELSIF x =- 22112 THEN
            exp_f := 0;
        ELSIF x =- 22111 THEN
            exp_f := 0;
        ELSIF x =- 22110 THEN
            exp_f := 0;
        ELSIF x =- 22109 THEN
            exp_f := 0;
        ELSIF x =- 22108 THEN
            exp_f := 0;
        ELSIF x =- 22107 THEN
            exp_f := 0;
        ELSIF x =- 22106 THEN
            exp_f := 0;
        ELSIF x =- 22105 THEN
            exp_f := 0;
        ELSIF x =- 22104 THEN
            exp_f := 0;
        ELSIF x =- 22103 THEN
            exp_f := 0;
        ELSIF x =- 22102 THEN
            exp_f := 0;
        ELSIF x =- 22101 THEN
            exp_f := 0;
        ELSIF x =- 22100 THEN
            exp_f := 0;
        ELSIF x =- 22099 THEN
            exp_f := 0;
        ELSIF x =- 22098 THEN
            exp_f := 0;
        ELSIF x =- 22097 THEN
            exp_f := 0;
        ELSIF x =- 22096 THEN
            exp_f := 0;
        ELSIF x =- 22095 THEN
            exp_f := 0;
        ELSIF x =- 22094 THEN
            exp_f := 0;
        ELSIF x =- 22093 THEN
            exp_f := 0;
        ELSIF x =- 22092 THEN
            exp_f := 0;
        ELSIF x =- 22091 THEN
            exp_f := 0;
        ELSIF x =- 22090 THEN
            exp_f := 0;
        ELSIF x =- 22089 THEN
            exp_f := 0;
        ELSIF x =- 22088 THEN
            exp_f := 0;
        ELSIF x =- 22087 THEN
            exp_f := 0;
        ELSIF x =- 22086 THEN
            exp_f := 0;
        ELSIF x =- 22085 THEN
            exp_f := 0;
        ELSIF x =- 22084 THEN
            exp_f := 0;
        ELSIF x =- 22083 THEN
            exp_f := 0;
        ELSIF x =- 22082 THEN
            exp_f := 0;
        ELSIF x =- 22081 THEN
            exp_f := 0;
        ELSIF x =- 22080 THEN
            exp_f := 0;
        ELSIF x =- 22079 THEN
            exp_f := 0;
        ELSIF x =- 22078 THEN
            exp_f := 0;
        ELSIF x =- 22077 THEN
            exp_f := 0;
        ELSIF x =- 22076 THEN
            exp_f := 0;
        ELSIF x =- 22075 THEN
            exp_f := 0;
        ELSIF x =- 22074 THEN
            exp_f := 0;
        ELSIF x =- 22073 THEN
            exp_f := 0;
        ELSIF x =- 22072 THEN
            exp_f := 0;
        ELSIF x =- 22071 THEN
            exp_f := 0;
        ELSIF x =- 22070 THEN
            exp_f := 0;
        ELSIF x =- 22069 THEN
            exp_f := 0;
        ELSIF x =- 22068 THEN
            exp_f := 0;
        ELSIF x =- 22067 THEN
            exp_f := 0;
        ELSIF x =- 22066 THEN
            exp_f := 0;
        ELSIF x =- 22065 THEN
            exp_f := 0;
        ELSIF x =- 22064 THEN
            exp_f := 0;
        ELSIF x =- 22063 THEN
            exp_f := 0;
        ELSIF x =- 22062 THEN
            exp_f := 0;
        ELSIF x =- 22061 THEN
            exp_f := 0;
        ELSIF x =- 22060 THEN
            exp_f := 0;
        ELSIF x =- 22059 THEN
            exp_f := 0;
        ELSIF x =- 22058 THEN
            exp_f := 0;
        ELSIF x =- 22057 THEN
            exp_f := 0;
        ELSIF x =- 22056 THEN
            exp_f := 0;
        ELSIF x =- 22055 THEN
            exp_f := 0;
        ELSIF x =- 22054 THEN
            exp_f := 0;
        ELSIF x =- 22053 THEN
            exp_f := 0;
        ELSIF x =- 22052 THEN
            exp_f := 0;
        ELSIF x =- 22051 THEN
            exp_f := 0;
        ELSIF x =- 22050 THEN
            exp_f := 0;
        ELSIF x =- 22049 THEN
            exp_f := 0;
        ELSIF x =- 22048 THEN
            exp_f := 0;
        ELSIF x =- 22047 THEN
            exp_f := 0;
        ELSIF x =- 22046 THEN
            exp_f := 0;
        ELSIF x =- 22045 THEN
            exp_f := 0;
        ELSIF x =- 22044 THEN
            exp_f := 0;
        ELSIF x =- 22043 THEN
            exp_f := 0;
        ELSIF x =- 22042 THEN
            exp_f := 0;
        ELSIF x =- 22041 THEN
            exp_f := 0;
        ELSIF x =- 22040 THEN
            exp_f := 0;
        ELSIF x =- 22039 THEN
            exp_f := 0;
        ELSIF x =- 22038 THEN
            exp_f := 0;
        ELSIF x =- 22037 THEN
            exp_f := 0;
        ELSIF x =- 22036 THEN
            exp_f := 0;
        ELSIF x =- 22035 THEN
            exp_f := 0;
        ELSIF x =- 22034 THEN
            exp_f := 0;
        ELSIF x =- 22033 THEN
            exp_f := 0;
        ELSIF x =- 22032 THEN
            exp_f := 0;
        ELSIF x =- 22031 THEN
            exp_f := 0;
        ELSIF x =- 22030 THEN
            exp_f := 0;
        ELSIF x =- 22029 THEN
            exp_f := 0;
        ELSIF x =- 22028 THEN
            exp_f := 0;
        ELSIF x =- 22027 THEN
            exp_f := 0;
        ELSIF x =- 22026 THEN
            exp_f := 0;
        ELSIF x =- 22025 THEN
            exp_f := 0;
        ELSIF x =- 22024 THEN
            exp_f := 0;
        ELSIF x =- 22023 THEN
            exp_f := 0;
        ELSIF x =- 22022 THEN
            exp_f := 0;
        ELSIF x =- 22021 THEN
            exp_f := 0;
        ELSIF x =- 22020 THEN
            exp_f := 0;
        ELSIF x =- 22019 THEN
            exp_f := 0;
        ELSIF x =- 22018 THEN
            exp_f := 0;
        ELSIF x =- 22017 THEN
            exp_f := 0;
        ELSIF x =- 22016 THEN
            exp_f := 0;
        ELSIF x =- 22015 THEN
            exp_f := 0;
        ELSIF x =- 22014 THEN
            exp_f := 0;
        ELSIF x =- 22013 THEN
            exp_f := 0;
        ELSIF x =- 22012 THEN
            exp_f := 0;
        ELSIF x =- 22011 THEN
            exp_f := 0;
        ELSIF x =- 22010 THEN
            exp_f := 0;
        ELSIF x =- 22009 THEN
            exp_f := 0;
        ELSIF x =- 22008 THEN
            exp_f := 0;
        ELSIF x =- 22007 THEN
            exp_f := 0;
        ELSIF x =- 22006 THEN
            exp_f := 0;
        ELSIF x =- 22005 THEN
            exp_f := 0;
        ELSIF x =- 22004 THEN
            exp_f := 0;
        ELSIF x =- 22003 THEN
            exp_f := 0;
        ELSIF x =- 22002 THEN
            exp_f := 0;
        ELSIF x =- 22001 THEN
            exp_f := 0;
        ELSIF x =- 22000 THEN
            exp_f := 0;
        ELSIF x =- 21999 THEN
            exp_f := 0;
        ELSIF x =- 21998 THEN
            exp_f := 0;
        ELSIF x =- 21997 THEN
            exp_f := 0;
        ELSIF x =- 21996 THEN
            exp_f := 0;
        ELSIF x =- 21995 THEN
            exp_f := 0;
        ELSIF x =- 21994 THEN
            exp_f := 0;
        ELSIF x =- 21993 THEN
            exp_f := 0;
        ELSIF x =- 21992 THEN
            exp_f := 0;
        ELSIF x =- 21991 THEN
            exp_f := 0;
        ELSIF x =- 21990 THEN
            exp_f := 0;
        ELSIF x =- 21989 THEN
            exp_f := 0;
        ELSIF x =- 21988 THEN
            exp_f := 0;
        ELSIF x =- 21987 THEN
            exp_f := 0;
        ELSIF x =- 21986 THEN
            exp_f := 0;
        ELSIF x =- 21985 THEN
            exp_f := 0;
        ELSIF x =- 21984 THEN
            exp_f := 0;
        ELSIF x =- 21983 THEN
            exp_f := 0;
        ELSIF x =- 21982 THEN
            exp_f := 0;
        ELSIF x =- 21981 THEN
            exp_f := 0;
        ELSIF x =- 21980 THEN
            exp_f := 0;
        ELSIF x =- 21979 THEN
            exp_f := 0;
        ELSIF x =- 21978 THEN
            exp_f := 0;
        ELSIF x =- 21977 THEN
            exp_f := 0;
        ELSIF x =- 21976 THEN
            exp_f := 0;
        ELSIF x =- 21975 THEN
            exp_f := 0;
        ELSIF x =- 21974 THEN
            exp_f := 0;
        ELSIF x =- 21973 THEN
            exp_f := 0;
        ELSIF x =- 21972 THEN
            exp_f := 0;
        ELSIF x =- 21971 THEN
            exp_f := 0;
        ELSIF x =- 21970 THEN
            exp_f := 0;
        ELSIF x =- 21969 THEN
            exp_f := 0;
        ELSIF x =- 21968 THEN
            exp_f := 0;
        ELSIF x =- 21967 THEN
            exp_f := 0;
        ELSIF x =- 21966 THEN
            exp_f := 0;
        ELSIF x =- 21965 THEN
            exp_f := 0;
        ELSIF x =- 21964 THEN
            exp_f := 0;
        ELSIF x =- 21963 THEN
            exp_f := 0;
        ELSIF x =- 21962 THEN
            exp_f := 0;
        ELSIF x =- 21961 THEN
            exp_f := 0;
        ELSIF x =- 21960 THEN
            exp_f := 0;
        ELSIF x =- 21959 THEN
            exp_f := 0;
        ELSIF x =- 21958 THEN
            exp_f := 0;
        ELSIF x =- 21957 THEN
            exp_f := 0;
        ELSIF x =- 21956 THEN
            exp_f := 0;
        ELSIF x =- 21955 THEN
            exp_f := 0;
        ELSIF x =- 21954 THEN
            exp_f := 0;
        ELSIF x =- 21953 THEN
            exp_f := 0;
        ELSIF x =- 21952 THEN
            exp_f := 0;
        ELSIF x =- 21951 THEN
            exp_f := 0;
        ELSIF x =- 21950 THEN
            exp_f := 0;
        ELSIF x =- 21949 THEN
            exp_f := 0;
        ELSIF x =- 21948 THEN
            exp_f := 0;
        ELSIF x =- 21947 THEN
            exp_f := 0;
        ELSIF x =- 21946 THEN
            exp_f := 0;
        ELSIF x =- 21945 THEN
            exp_f := 0;
        ELSIF x =- 21944 THEN
            exp_f := 0;
        ELSIF x =- 21943 THEN
            exp_f := 0;
        ELSIF x =- 21942 THEN
            exp_f := 0;
        ELSIF x =- 21941 THEN
            exp_f := 0;
        ELSIF x =- 21940 THEN
            exp_f := 0;
        ELSIF x =- 21939 THEN
            exp_f := 0;
        ELSIF x =- 21938 THEN
            exp_f := 0;
        ELSIF x =- 21937 THEN
            exp_f := 0;
        ELSIF x =- 21936 THEN
            exp_f := 0;
        ELSIF x =- 21935 THEN
            exp_f := 0;
        ELSIF x =- 21934 THEN
            exp_f := 0;
        ELSIF x =- 21933 THEN
            exp_f := 0;
        ELSIF x =- 21932 THEN
            exp_f := 0;
        ELSIF x =- 21931 THEN
            exp_f := 0;
        ELSIF x =- 21930 THEN
            exp_f := 0;
        ELSIF x =- 21929 THEN
            exp_f := 0;
        ELSIF x =- 21928 THEN
            exp_f := 0;
        ELSIF x =- 21927 THEN
            exp_f := 0;
        ELSIF x =- 21926 THEN
            exp_f := 0;
        ELSIF x =- 21925 THEN
            exp_f := 0;
        ELSIF x =- 21924 THEN
            exp_f := 0;
        ELSIF x =- 21923 THEN
            exp_f := 0;
        ELSIF x =- 21922 THEN
            exp_f := 0;
        ELSIF x =- 21921 THEN
            exp_f := 0;
        ELSIF x =- 21920 THEN
            exp_f := 0;
        ELSIF x =- 21919 THEN
            exp_f := 0;
        ELSIF x =- 21918 THEN
            exp_f := 0;
        ELSIF x =- 21917 THEN
            exp_f := 0;
        ELSIF x =- 21916 THEN
            exp_f := 0;
        ELSIF x =- 21915 THEN
            exp_f := 0;
        ELSIF x =- 21914 THEN
            exp_f := 0;
        ELSIF x =- 21913 THEN
            exp_f := 0;
        ELSIF x =- 21912 THEN
            exp_f := 0;
        ELSIF x =- 21911 THEN
            exp_f := 0;
        ELSIF x =- 21910 THEN
            exp_f := 0;
        ELSIF x =- 21909 THEN
            exp_f := 0;
        ELSIF x =- 21908 THEN
            exp_f := 0;
        ELSIF x =- 21907 THEN
            exp_f := 0;
        ELSIF x =- 21906 THEN
            exp_f := 0;
        ELSIF x =- 21905 THEN
            exp_f := 0;
        ELSIF x =- 21904 THEN
            exp_f := 0;
        ELSIF x =- 21903 THEN
            exp_f := 0;
        ELSIF x =- 21902 THEN
            exp_f := 0;
        ELSIF x =- 21901 THEN
            exp_f := 0;
        ELSIF x =- 21900 THEN
            exp_f := 0;
        ELSIF x =- 21899 THEN
            exp_f := 0;
        ELSIF x =- 21898 THEN
            exp_f := 0;
        ELSIF x =- 21897 THEN
            exp_f := 0;
        ELSIF x =- 21896 THEN
            exp_f := 0;
        ELSIF x =- 21895 THEN
            exp_f := 0;
        ELSIF x =- 21894 THEN
            exp_f := 0;
        ELSIF x =- 21893 THEN
            exp_f := 0;
        ELSIF x =- 21892 THEN
            exp_f := 0;
        ELSIF x =- 21891 THEN
            exp_f := 0;
        ELSIF x =- 21890 THEN
            exp_f := 0;
        ELSIF x =- 21889 THEN
            exp_f := 0;
        ELSIF x =- 21888 THEN
            exp_f := 0;
        ELSIF x =- 21887 THEN
            exp_f := 0;
        ELSIF x =- 21886 THEN
            exp_f := 0;
        ELSIF x =- 21885 THEN
            exp_f := 0;
        ELSIF x =- 21884 THEN
            exp_f := 0;
        ELSIF x =- 21883 THEN
            exp_f := 0;
        ELSIF x =- 21882 THEN
            exp_f := 0;
        ELSIF x =- 21881 THEN
            exp_f := 0;
        ELSIF x =- 21880 THEN
            exp_f := 0;
        ELSIF x =- 21879 THEN
            exp_f := 0;
        ELSIF x =- 21878 THEN
            exp_f := 0;
        ELSIF x =- 21877 THEN
            exp_f := 0;
        ELSIF x =- 21876 THEN
            exp_f := 0;
        ELSIF x =- 21875 THEN
            exp_f := 0;
        ELSIF x =- 21874 THEN
            exp_f := 0;
        ELSIF x =- 21873 THEN
            exp_f := 0;
        ELSIF x =- 21872 THEN
            exp_f := 0;
        ELSIF x =- 21871 THEN
            exp_f := 0;
        ELSIF x =- 21870 THEN
            exp_f := 0;
        ELSIF x =- 21869 THEN
            exp_f := 0;
        ELSIF x =- 21868 THEN
            exp_f := 0;
        ELSIF x =- 21867 THEN
            exp_f := 0;
        ELSIF x =- 21866 THEN
            exp_f := 0;
        ELSIF x =- 21865 THEN
            exp_f := 0;
        ELSIF x =- 21864 THEN
            exp_f := 0;
        ELSIF x =- 21863 THEN
            exp_f := 0;
        ELSIF x =- 21862 THEN
            exp_f := 0;
        ELSIF x =- 21861 THEN
            exp_f := 0;
        ELSIF x =- 21860 THEN
            exp_f := 0;
        ELSIF x =- 21859 THEN
            exp_f := 0;
        ELSIF x =- 21858 THEN
            exp_f := 0;
        ELSIF x =- 21857 THEN
            exp_f := 0;
        ELSIF x =- 21856 THEN
            exp_f := 0;
        ELSIF x =- 21855 THEN
            exp_f := 0;
        ELSIF x =- 21854 THEN
            exp_f := 0;
        ELSIF x =- 21853 THEN
            exp_f := 0;
        ELSIF x =- 21852 THEN
            exp_f := 0;
        ELSIF x =- 21851 THEN
            exp_f := 0;
        ELSIF x =- 21850 THEN
            exp_f := 0;
        ELSIF x =- 21849 THEN
            exp_f := 0;
        ELSIF x =- 21848 THEN
            exp_f := 0;
        ELSIF x =- 21847 THEN
            exp_f := 0;
        ELSIF x =- 21846 THEN
            exp_f := 0;
        ELSIF x =- 21845 THEN
            exp_f := 0;
        ELSIF x =- 21844 THEN
            exp_f := 0;
        ELSIF x =- 21843 THEN
            exp_f := 0;
        ELSIF x =- 21842 THEN
            exp_f := 0;
        ELSIF x =- 21841 THEN
            exp_f := 0;
        ELSIF x =- 21840 THEN
            exp_f := 0;
        ELSIF x =- 21839 THEN
            exp_f := 0;
        ELSIF x =- 21838 THEN
            exp_f := 0;
        ELSIF x =- 21837 THEN
            exp_f := 0;
        ELSIF x =- 21836 THEN
            exp_f := 0;
        ELSIF x =- 21835 THEN
            exp_f := 0;
        ELSIF x =- 21834 THEN
            exp_f := 0;
        ELSIF x =- 21833 THEN
            exp_f := 0;
        ELSIF x =- 21832 THEN
            exp_f := 0;
        ELSIF x =- 21831 THEN
            exp_f := 0;
        ELSIF x =- 21830 THEN
            exp_f := 0;
        ELSIF x =- 21829 THEN
            exp_f := 0;
        ELSIF x =- 21828 THEN
            exp_f := 0;
        ELSIF x =- 21827 THEN
            exp_f := 0;
        ELSIF x =- 21826 THEN
            exp_f := 0;
        ELSIF x =- 21825 THEN
            exp_f := 0;
        ELSIF x =- 21824 THEN
            exp_f := 0;
        ELSIF x =- 21823 THEN
            exp_f := 0;
        ELSIF x =- 21822 THEN
            exp_f := 0;
        ELSIF x =- 21821 THEN
            exp_f := 0;
        ELSIF x =- 21820 THEN
            exp_f := 0;
        ELSIF x =- 21819 THEN
            exp_f := 0;
        ELSIF x =- 21818 THEN
            exp_f := 0;
        ELSIF x =- 21817 THEN
            exp_f := 0;
        ELSIF x =- 21816 THEN
            exp_f := 0;
        ELSIF x =- 21815 THEN
            exp_f := 0;
        ELSIF x =- 21814 THEN
            exp_f := 0;
        ELSIF x =- 21813 THEN
            exp_f := 0;
        ELSIF x =- 21812 THEN
            exp_f := 0;
        ELSIF x =- 21811 THEN
            exp_f := 0;
        ELSIF x =- 21810 THEN
            exp_f := 0;
        ELSIF x =- 21809 THEN
            exp_f := 0;
        ELSIF x =- 21808 THEN
            exp_f := 0;
        ELSIF x =- 21807 THEN
            exp_f := 0;
        ELSIF x =- 21806 THEN
            exp_f := 0;
        ELSIF x =- 21805 THEN
            exp_f := 0;
        ELSIF x =- 21804 THEN
            exp_f := 0;
        ELSIF x =- 21803 THEN
            exp_f := 0;
        ELSIF x =- 21802 THEN
            exp_f := 0;
        ELSIF x =- 21801 THEN
            exp_f := 0;
        ELSIF x =- 21800 THEN
            exp_f := 0;
        ELSIF x =- 21799 THEN
            exp_f := 0;
        ELSIF x =- 21798 THEN
            exp_f := 0;
        ELSIF x =- 21797 THEN
            exp_f := 0;
        ELSIF x =- 21796 THEN
            exp_f := 0;
        ELSIF x =- 21795 THEN
            exp_f := 0;
        ELSIF x =- 21794 THEN
            exp_f := 0;
        ELSIF x =- 21793 THEN
            exp_f := 0;
        ELSIF x =- 21792 THEN
            exp_f := 0;
        ELSIF x =- 21791 THEN
            exp_f := 0;
        ELSIF x =- 21790 THEN
            exp_f := 0;
        ELSIF x =- 21789 THEN
            exp_f := 0;
        ELSIF x =- 21788 THEN
            exp_f := 0;
        ELSIF x =- 21787 THEN
            exp_f := 0;
        ELSIF x =- 21786 THEN
            exp_f := 0;
        ELSIF x =- 21785 THEN
            exp_f := 0;
        ELSIF x =- 21784 THEN
            exp_f := 0;
        ELSIF x =- 21783 THEN
            exp_f := 0;
        ELSIF x =- 21782 THEN
            exp_f := 0;
        ELSIF x =- 21781 THEN
            exp_f := 0;
        ELSIF x =- 21780 THEN
            exp_f := 0;
        ELSIF x =- 21779 THEN
            exp_f := 0;
        ELSIF x =- 21778 THEN
            exp_f := 0;
        ELSIF x =- 21777 THEN
            exp_f := 0;
        ELSIF x =- 21776 THEN
            exp_f := 0;
        ELSIF x =- 21775 THEN
            exp_f := 0;
        ELSIF x =- 21774 THEN
            exp_f := 0;
        ELSIF x =- 21773 THEN
            exp_f := 0;
        ELSIF x =- 21772 THEN
            exp_f := 0;
        ELSIF x =- 21771 THEN
            exp_f := 0;
        ELSIF x =- 21770 THEN
            exp_f := 0;
        ELSIF x =- 21769 THEN
            exp_f := 0;
        ELSIF x =- 21768 THEN
            exp_f := 0;
        ELSIF x =- 21767 THEN
            exp_f := 0;
        ELSIF x =- 21766 THEN
            exp_f := 0;
        ELSIF x =- 21765 THEN
            exp_f := 0;
        ELSIF x =- 21764 THEN
            exp_f := 0;
        ELSIF x =- 21763 THEN
            exp_f := 0;
        ELSIF x =- 21762 THEN
            exp_f := 0;
        ELSIF x =- 21761 THEN
            exp_f := 0;
        ELSIF x =- 21760 THEN
            exp_f := 0;
        ELSIF x =- 21759 THEN
            exp_f := 0;
        ELSIF x =- 21758 THEN
            exp_f := 0;
        ELSIF x =- 21757 THEN
            exp_f := 0;
        ELSIF x =- 21756 THEN
            exp_f := 0;
        ELSIF x =- 21755 THEN
            exp_f := 0;
        ELSIF x =- 21754 THEN
            exp_f := 0;
        ELSIF x =- 21753 THEN
            exp_f := 0;
        ELSIF x =- 21752 THEN
            exp_f := 0;
        ELSIF x =- 21751 THEN
            exp_f := 0;
        ELSIF x =- 21750 THEN
            exp_f := 0;
        ELSIF x =- 21749 THEN
            exp_f := 0;
        ELSIF x =- 21748 THEN
            exp_f := 0;
        ELSIF x =- 21747 THEN
            exp_f := 0;
        ELSIF x =- 21746 THEN
            exp_f := 0;
        ELSIF x =- 21745 THEN
            exp_f := 0;
        ELSIF x =- 21744 THEN
            exp_f := 0;
        ELSIF x =- 21743 THEN
            exp_f := 0;
        ELSIF x =- 21742 THEN
            exp_f := 0;
        ELSIF x =- 21741 THEN
            exp_f := 0;
        ELSIF x =- 21740 THEN
            exp_f := 0;
        ELSIF x =- 21739 THEN
            exp_f := 0;
        ELSIF x =- 21738 THEN
            exp_f := 0;
        ELSIF x =- 21737 THEN
            exp_f := 0;
        ELSIF x =- 21736 THEN
            exp_f := 0;
        ELSIF x =- 21735 THEN
            exp_f := 0;
        ELSIF x =- 21734 THEN
            exp_f := 0;
        ELSIF x =- 21733 THEN
            exp_f := 0;
        ELSIF x =- 21732 THEN
            exp_f := 0;
        ELSIF x =- 21731 THEN
            exp_f := 0;
        ELSIF x =- 21730 THEN
            exp_f := 0;
        ELSIF x =- 21729 THEN
            exp_f := 0;
        ELSIF x =- 21728 THEN
            exp_f := 0;
        ELSIF x =- 21727 THEN
            exp_f := 0;
        ELSIF x =- 21726 THEN
            exp_f := 0;
        ELSIF x =- 21725 THEN
            exp_f := 0;
        ELSIF x =- 21724 THEN
            exp_f := 0;
        ELSIF x =- 21723 THEN
            exp_f := 0;
        ELSIF x =- 21722 THEN
            exp_f := 0;
        ELSIF x =- 21721 THEN
            exp_f := 0;
        ELSIF x =- 21720 THEN
            exp_f := 0;
        ELSIF x =- 21719 THEN
            exp_f := 0;
        ELSIF x =- 21718 THEN
            exp_f := 0;
        ELSIF x =- 21717 THEN
            exp_f := 0;
        ELSIF x =- 21716 THEN
            exp_f := 0;
        ELSIF x =- 21715 THEN
            exp_f := 0;
        ELSIF x =- 21714 THEN
            exp_f := 0;
        ELSIF x =- 21713 THEN
            exp_f := 0;
        ELSIF x =- 21712 THEN
            exp_f := 0;
        ELSIF x =- 21711 THEN
            exp_f := 0;
        ELSIF x =- 21710 THEN
            exp_f := 0;
        ELSIF x =- 21709 THEN
            exp_f := 0;
        ELSIF x =- 21708 THEN
            exp_f := 0;
        ELSIF x =- 21707 THEN
            exp_f := 0;
        ELSIF x =- 21706 THEN
            exp_f := 0;
        ELSIF x =- 21705 THEN
            exp_f := 0;
        ELSIF x =- 21704 THEN
            exp_f := 0;
        ELSIF x =- 21703 THEN
            exp_f := 0;
        ELSIF x =- 21702 THEN
            exp_f := 0;
        ELSIF x =- 21701 THEN
            exp_f := 0;
        ELSIF x =- 21700 THEN
            exp_f := 0;
        ELSIF x =- 21699 THEN
            exp_f := 0;
        ELSIF x =- 21698 THEN
            exp_f := 0;
        ELSIF x =- 21697 THEN
            exp_f := 0;
        ELSIF x =- 21696 THEN
            exp_f := 0;
        ELSIF x =- 21695 THEN
            exp_f := 0;
        ELSIF x =- 21694 THEN
            exp_f := 0;
        ELSIF x =- 21693 THEN
            exp_f := 0;
        ELSIF x =- 21692 THEN
            exp_f := 0;
        ELSIF x =- 21691 THEN
            exp_f := 0;
        ELSIF x =- 21690 THEN
            exp_f := 0;
        ELSIF x =- 21689 THEN
            exp_f := 0;
        ELSIF x =- 21688 THEN
            exp_f := 0;
        ELSIF x =- 21687 THEN
            exp_f := 0;
        ELSIF x =- 21686 THEN
            exp_f := 0;
        ELSIF x =- 21685 THEN
            exp_f := 0;
        ELSIF x =- 21684 THEN
            exp_f := 0;
        ELSIF x =- 21683 THEN
            exp_f := 0;
        ELSIF x =- 21682 THEN
            exp_f := 0;
        ELSIF x =- 21681 THEN
            exp_f := 0;
        ELSIF x =- 21680 THEN
            exp_f := 0;
        ELSIF x =- 21679 THEN
            exp_f := 0;
        ELSIF x =- 21678 THEN
            exp_f := 0;
        ELSIF x =- 21677 THEN
            exp_f := 0;
        ELSIF x =- 21676 THEN
            exp_f := 0;
        ELSIF x =- 21675 THEN
            exp_f := 0;
        ELSIF x =- 21674 THEN
            exp_f := 0;
        ELSIF x =- 21673 THEN
            exp_f := 0;
        ELSIF x =- 21672 THEN
            exp_f := 0;
        ELSIF x =- 21671 THEN
            exp_f := 0;
        ELSIF x =- 21670 THEN
            exp_f := 0;
        ELSIF x =- 21669 THEN
            exp_f := 0;
        ELSIF x =- 21668 THEN
            exp_f := 0;
        ELSIF x =- 21667 THEN
            exp_f := 0;
        ELSIF x =- 21666 THEN
            exp_f := 0;
        ELSIF x =- 21665 THEN
            exp_f := 0;
        ELSIF x =- 21664 THEN
            exp_f := 0;
        ELSIF x =- 21663 THEN
            exp_f := 0;
        ELSIF x =- 21662 THEN
            exp_f := 0;
        ELSIF x =- 21661 THEN
            exp_f := 0;
        ELSIF x =- 21660 THEN
            exp_f := 0;
        ELSIF x =- 21659 THEN
            exp_f := 0;
        ELSIF x =- 21658 THEN
            exp_f := 0;
        ELSIF x =- 21657 THEN
            exp_f := 0;
        ELSIF x =- 21656 THEN
            exp_f := 0;
        ELSIF x =- 21655 THEN
            exp_f := 0;
        ELSIF x =- 21654 THEN
            exp_f := 0;
        ELSIF x =- 21653 THEN
            exp_f := 0;
        ELSIF x =- 21652 THEN
            exp_f := 0;
        ELSIF x =- 21651 THEN
            exp_f := 0;
        ELSIF x =- 21650 THEN
            exp_f := 0;
        ELSIF x =- 21649 THEN
            exp_f := 0;
        ELSIF x =- 21648 THEN
            exp_f := 0;
        ELSIF x =- 21647 THEN
            exp_f := 0;
        ELSIF x =- 21646 THEN
            exp_f := 0;
        ELSIF x =- 21645 THEN
            exp_f := 0;
        ELSIF x =- 21644 THEN
            exp_f := 0;
        ELSIF x =- 21643 THEN
            exp_f := 0;
        ELSIF x =- 21642 THEN
            exp_f := 0;
        ELSIF x =- 21641 THEN
            exp_f := 0;
        ELSIF x =- 21640 THEN
            exp_f := 0;
        ELSIF x =- 21639 THEN
            exp_f := 0;
        ELSIF x =- 21638 THEN
            exp_f := 0;
        ELSIF x =- 21637 THEN
            exp_f := 0;
        ELSIF x =- 21636 THEN
            exp_f := 0;
        ELSIF x =- 21635 THEN
            exp_f := 0;
        ELSIF x =- 21634 THEN
            exp_f := 0;
        ELSIF x =- 21633 THEN
            exp_f := 0;
        ELSIF x =- 21632 THEN
            exp_f := 0;
        ELSIF x =- 21631 THEN
            exp_f := 0;
        ELSIF x =- 21630 THEN
            exp_f := 0;
        ELSIF x =- 21629 THEN
            exp_f := 0;
        ELSIF x =- 21628 THEN
            exp_f := 0;
        ELSIF x =- 21627 THEN
            exp_f := 0;
        ELSIF x =- 21626 THEN
            exp_f := 0;
        ELSIF x =- 21625 THEN
            exp_f := 0;
        ELSIF x =- 21624 THEN
            exp_f := 0;
        ELSIF x =- 21623 THEN
            exp_f := 0;
        ELSIF x =- 21622 THEN
            exp_f := 0;
        ELSIF x =- 21621 THEN
            exp_f := 0;
        ELSIF x =- 21620 THEN
            exp_f := 0;
        ELSIF x =- 21619 THEN
            exp_f := 0;
        ELSIF x =- 21618 THEN
            exp_f := 0;
        ELSIF x =- 21617 THEN
            exp_f := 0;
        ELSIF x =- 21616 THEN
            exp_f := 0;
        ELSIF x =- 21615 THEN
            exp_f := 0;
        ELSIF x =- 21614 THEN
            exp_f := 0;
        ELSIF x =- 21613 THEN
            exp_f := 0;
        ELSIF x =- 21612 THEN
            exp_f := 0;
        ELSIF x =- 21611 THEN
            exp_f := 0;
        ELSIF x =- 21610 THEN
            exp_f := 0;
        ELSIF x =- 21609 THEN
            exp_f := 0;
        ELSIF x =- 21608 THEN
            exp_f := 0;
        ELSIF x =- 21607 THEN
            exp_f := 0;
        ELSIF x =- 21606 THEN
            exp_f := 0;
        ELSIF x =- 21605 THEN
            exp_f := 0;
        ELSIF x =- 21604 THEN
            exp_f := 0;
        ELSIF x =- 21603 THEN
            exp_f := 0;
        ELSIF x =- 21602 THEN
            exp_f := 0;
        ELSIF x =- 21601 THEN
            exp_f := 0;
        ELSIF x =- 21600 THEN
            exp_f := 0;
        ELSIF x =- 21599 THEN
            exp_f := 0;
        ELSIF x =- 21598 THEN
            exp_f := 0;
        ELSIF x =- 21597 THEN
            exp_f := 0;
        ELSIF x =- 21596 THEN
            exp_f := 0;
        ELSIF x =- 21595 THEN
            exp_f := 0;
        ELSIF x =- 21594 THEN
            exp_f := 0;
        ELSIF x =- 21593 THEN
            exp_f := 0;
        ELSIF x =- 21592 THEN
            exp_f := 0;
        ELSIF x =- 21591 THEN
            exp_f := 0;
        ELSIF x =- 21590 THEN
            exp_f := 0;
        ELSIF x =- 21589 THEN
            exp_f := 0;
        ELSIF x =- 21588 THEN
            exp_f := 0;
        ELSIF x =- 21587 THEN
            exp_f := 0;
        ELSIF x =- 21586 THEN
            exp_f := 0;
        ELSIF x =- 21585 THEN
            exp_f := 0;
        ELSIF x =- 21584 THEN
            exp_f := 0;
        ELSIF x =- 21583 THEN
            exp_f := 0;
        ELSIF x =- 21582 THEN
            exp_f := 0;
        ELSIF x =- 21581 THEN
            exp_f := 0;
        ELSIF x =- 21580 THEN
            exp_f := 0;
        ELSIF x =- 21579 THEN
            exp_f := 0;
        ELSIF x =- 21578 THEN
            exp_f := 0;
        ELSIF x =- 21577 THEN
            exp_f := 0;
        ELSIF x =- 21576 THEN
            exp_f := 0;
        ELSIF x =- 21575 THEN
            exp_f := 0;
        ELSIF x =- 21574 THEN
            exp_f := 0;
        ELSIF x =- 21573 THEN
            exp_f := 0;
        ELSIF x =- 21572 THEN
            exp_f := 0;
        ELSIF x =- 21571 THEN
            exp_f := 0;
        ELSIF x =- 21570 THEN
            exp_f := 0;
        ELSIF x =- 21569 THEN
            exp_f := 0;
        ELSIF x =- 21568 THEN
            exp_f := 0;
        ELSIF x =- 21567 THEN
            exp_f := 0;
        ELSIF x =- 21566 THEN
            exp_f := 0;
        ELSIF x =- 21565 THEN
            exp_f := 0;
        ELSIF x =- 21564 THEN
            exp_f := 0;
        ELSIF x =- 21563 THEN
            exp_f := 0;
        ELSIF x =- 21562 THEN
            exp_f := 0;
        ELSIF x =- 21561 THEN
            exp_f := 0;
        ELSIF x =- 21560 THEN
            exp_f := 0;
        ELSIF x =- 21559 THEN
            exp_f := 0;
        ELSIF x =- 21558 THEN
            exp_f := 0;
        ELSIF x =- 21557 THEN
            exp_f := 0;
        ELSIF x =- 21556 THEN
            exp_f := 0;
        ELSIF x =- 21555 THEN
            exp_f := 0;
        ELSIF x =- 21554 THEN
            exp_f := 0;
        ELSIF x =- 21553 THEN
            exp_f := 0;
        ELSIF x =- 21552 THEN
            exp_f := 0;
        ELSIF x =- 21551 THEN
            exp_f := 0;
        ELSIF x =- 21550 THEN
            exp_f := 0;
        ELSIF x =- 21549 THEN
            exp_f := 0;
        ELSIF x =- 21548 THEN
            exp_f := 0;
        ELSIF x =- 21547 THEN
            exp_f := 0;
        ELSIF x =- 21546 THEN
            exp_f := 0;
        ELSIF x =- 21545 THEN
            exp_f := 0;
        ELSIF x =- 21544 THEN
            exp_f := 0;
        ELSIF x =- 21543 THEN
            exp_f := 0;
        ELSIF x =- 21542 THEN
            exp_f := 0;
        ELSIF x =- 21541 THEN
            exp_f := 0;
        ELSIF x =- 21540 THEN
            exp_f := 0;
        ELSIF x =- 21539 THEN
            exp_f := 0;
        ELSIF x =- 21538 THEN
            exp_f := 0;
        ELSIF x =- 21537 THEN
            exp_f := 0;
        ELSIF x =- 21536 THEN
            exp_f := 0;
        ELSIF x =- 21535 THEN
            exp_f := 0;
        ELSIF x =- 21534 THEN
            exp_f := 0;
        ELSIF x =- 21533 THEN
            exp_f := 0;
        ELSIF x =- 21532 THEN
            exp_f := 0;
        ELSIF x =- 21531 THEN
            exp_f := 0;
        ELSIF x =- 21530 THEN
            exp_f := 0;
        ELSIF x =- 21529 THEN
            exp_f := 0;
        ELSIF x =- 21528 THEN
            exp_f := 0;
        ELSIF x =- 21527 THEN
            exp_f := 0;
        ELSIF x =- 21526 THEN
            exp_f := 0;
        ELSIF x =- 21525 THEN
            exp_f := 0;
        ELSIF x =- 21524 THEN
            exp_f := 0;
        ELSIF x =- 21523 THEN
            exp_f := 0;
        ELSIF x =- 21522 THEN
            exp_f := 0;
        ELSIF x =- 21521 THEN
            exp_f := 0;
        ELSIF x =- 21520 THEN
            exp_f := 0;
        ELSIF x =- 21519 THEN
            exp_f := 0;
        ELSIF x =- 21518 THEN
            exp_f := 0;
        ELSIF x =- 21517 THEN
            exp_f := 0;
        ELSIF x =- 21516 THEN
            exp_f := 0;
        ELSIF x =- 21515 THEN
            exp_f := 0;
        ELSIF x =- 21514 THEN
            exp_f := 0;
        ELSIF x =- 21513 THEN
            exp_f := 0;
        ELSIF x =- 21512 THEN
            exp_f := 0;
        ELSIF x =- 21511 THEN
            exp_f := 0;
        ELSIF x =- 21510 THEN
            exp_f := 0;
        ELSIF x =- 21509 THEN
            exp_f := 0;
        ELSIF x =- 21508 THEN
            exp_f := 0;
        ELSIF x =- 21507 THEN
            exp_f := 0;
        ELSIF x =- 21506 THEN
            exp_f := 0;
        ELSIF x =- 21505 THEN
            exp_f := 0;
        ELSIF x =- 21504 THEN
            exp_f := 0;
        ELSIF x =- 21503 THEN
            exp_f := 0;
        ELSIF x =- 21502 THEN
            exp_f := 0;
        ELSIF x =- 21501 THEN
            exp_f := 0;
        ELSIF x =- 21500 THEN
            exp_f := 0;
        ELSIF x =- 21499 THEN
            exp_f := 0;
        ELSIF x =- 21498 THEN
            exp_f := 0;
        ELSIF x =- 21497 THEN
            exp_f := 0;
        ELSIF x =- 21496 THEN
            exp_f := 0;
        ELSIF x =- 21495 THEN
            exp_f := 0;
        ELSIF x =- 21494 THEN
            exp_f := 0;
        ELSIF x =- 21493 THEN
            exp_f := 0;
        ELSIF x =- 21492 THEN
            exp_f := 0;
        ELSIF x =- 21491 THEN
            exp_f := 0;
        ELSIF x =- 21490 THEN
            exp_f := 0;
        ELSIF x =- 21489 THEN
            exp_f := 0;
        ELSIF x =- 21488 THEN
            exp_f := 0;
        ELSIF x =- 21487 THEN
            exp_f := 0;
        ELSIF x =- 21486 THEN
            exp_f := 0;
        ELSIF x =- 21485 THEN
            exp_f := 0;
        ELSIF x =- 21484 THEN
            exp_f := 0;
        ELSIF x =- 21483 THEN
            exp_f := 0;
        ELSIF x =- 21482 THEN
            exp_f := 0;
        ELSIF x =- 21481 THEN
            exp_f := 0;
        ELSIF x =- 21480 THEN
            exp_f := 0;
        ELSIF x =- 21479 THEN
            exp_f := 0;
        ELSIF x =- 21478 THEN
            exp_f := 0;
        ELSIF x =- 21477 THEN
            exp_f := 0;
        ELSIF x =- 21476 THEN
            exp_f := 0;
        ELSIF x =- 21475 THEN
            exp_f := 0;
        ELSIF x =- 21474 THEN
            exp_f := 0;
        ELSIF x =- 21473 THEN
            exp_f := 0;
        ELSIF x =- 21472 THEN
            exp_f := 0;
        ELSIF x =- 21471 THEN
            exp_f := 0;
        ELSIF x =- 21470 THEN
            exp_f := 0;
        ELSIF x =- 21469 THEN
            exp_f := 0;
        ELSIF x =- 21468 THEN
            exp_f := 0;
        ELSIF x =- 21467 THEN
            exp_f := 0;
        ELSIF x =- 21466 THEN
            exp_f := 0;
        ELSIF x =- 21465 THEN
            exp_f := 0;
        ELSIF x =- 21464 THEN
            exp_f := 0;
        ELSIF x =- 21463 THEN
            exp_f := 0;
        ELSIF x =- 21462 THEN
            exp_f := 0;
        ELSIF x =- 21461 THEN
            exp_f := 0;
        ELSIF x =- 21460 THEN
            exp_f := 0;
        ELSIF x =- 21459 THEN
            exp_f := 0;
        ELSIF x =- 21458 THEN
            exp_f := 0;
        ELSIF x =- 21457 THEN
            exp_f := 0;
        ELSIF x =- 21456 THEN
            exp_f := 0;
        ELSIF x =- 21455 THEN
            exp_f := 0;
        ELSIF x =- 21454 THEN
            exp_f := 0;
        ELSIF x =- 21453 THEN
            exp_f := 0;
        ELSIF x =- 21452 THEN
            exp_f := 0;
        ELSIF x =- 21451 THEN
            exp_f := 0;
        ELSIF x =- 21450 THEN
            exp_f := 0;
        ELSIF x =- 21449 THEN
            exp_f := 0;
        ELSIF x =- 21448 THEN
            exp_f := 0;
        ELSIF x =- 21447 THEN
            exp_f := 0;
        ELSIF x =- 21446 THEN
            exp_f := 0;
        ELSIF x =- 21445 THEN
            exp_f := 0;
        ELSIF x =- 21444 THEN
            exp_f := 0;
        ELSIF x =- 21443 THEN
            exp_f := 0;
        ELSIF x =- 21442 THEN
            exp_f := 0;
        ELSIF x =- 21441 THEN
            exp_f := 0;
        ELSIF x =- 21440 THEN
            exp_f := 0;
        ELSIF x =- 21439 THEN
            exp_f := 0;
        ELSIF x =- 21438 THEN
            exp_f := 0;
        ELSIF x =- 21437 THEN
            exp_f := 0;
        ELSIF x =- 21436 THEN
            exp_f := 0;
        ELSIF x =- 21435 THEN
            exp_f := 0;
        ELSIF x =- 21434 THEN
            exp_f := 0;
        ELSIF x =- 21433 THEN
            exp_f := 0;
        ELSIF x =- 21432 THEN
            exp_f := 0;
        ELSIF x =- 21431 THEN
            exp_f := 0;
        ELSIF x =- 21430 THEN
            exp_f := 0;
        ELSIF x =- 21429 THEN
            exp_f := 0;
        ELSIF x =- 21428 THEN
            exp_f := 0;
        ELSIF x =- 21427 THEN
            exp_f := 0;
        ELSIF x =- 21426 THEN
            exp_f := 0;
        ELSIF x =- 21425 THEN
            exp_f := 0;
        ELSIF x =- 21424 THEN
            exp_f := 0;
        ELSIF x =- 21423 THEN
            exp_f := 0;
        ELSIF x =- 21422 THEN
            exp_f := 0;
        ELSIF x =- 21421 THEN
            exp_f := 0;
        ELSIF x =- 21420 THEN
            exp_f := 0;
        ELSIF x =- 21419 THEN
            exp_f := 0;
        ELSIF x =- 21418 THEN
            exp_f := 0;
        ELSIF x =- 21417 THEN
            exp_f := 0;
        ELSIF x =- 21416 THEN
            exp_f := 0;
        ELSIF x =- 21415 THEN
            exp_f := 0;
        ELSIF x =- 21414 THEN
            exp_f := 0;
        ELSIF x =- 21413 THEN
            exp_f := 0;
        ELSIF x =- 21412 THEN
            exp_f := 0;
        ELSIF x =- 21411 THEN
            exp_f := 0;
        ELSIF x =- 21410 THEN
            exp_f := 0;
        ELSIF x =- 21409 THEN
            exp_f := 0;
        ELSIF x =- 21408 THEN
            exp_f := 0;
        ELSIF x =- 21407 THEN
            exp_f := 0;
        ELSIF x =- 21406 THEN
            exp_f := 0;
        ELSIF x =- 21405 THEN
            exp_f := 0;
        ELSIF x =- 21404 THEN
            exp_f := 0;
        ELSIF x =- 21403 THEN
            exp_f := 0;
        ELSIF x =- 21402 THEN
            exp_f := 0;
        ELSIF x =- 21401 THEN
            exp_f := 0;
        ELSIF x =- 21400 THEN
            exp_f := 0;
        ELSIF x =- 21399 THEN
            exp_f := 0;
        ELSIF x =- 21398 THEN
            exp_f := 0;
        ELSIF x =- 21397 THEN
            exp_f := 0;
        ELSIF x =- 21396 THEN
            exp_f := 0;
        ELSIF x =- 21395 THEN
            exp_f := 0;
        ELSIF x =- 21394 THEN
            exp_f := 0;
        ELSIF x =- 21393 THEN
            exp_f := 0;
        ELSIF x =- 21392 THEN
            exp_f := 0;
        ELSIF x =- 21391 THEN
            exp_f := 0;
        ELSIF x =- 21390 THEN
            exp_f := 0;
        ELSIF x =- 21389 THEN
            exp_f := 0;
        ELSIF x =- 21388 THEN
            exp_f := 0;
        ELSIF x =- 21387 THEN
            exp_f := 0;
        ELSIF x =- 21386 THEN
            exp_f := 0;
        ELSIF x =- 21385 THEN
            exp_f := 0;
        ELSIF x =- 21384 THEN
            exp_f := 0;
        ELSIF x =- 21383 THEN
            exp_f := 0;
        ELSIF x =- 21382 THEN
            exp_f := 0;
        ELSIF x =- 21381 THEN
            exp_f := 0;
        ELSIF x =- 21380 THEN
            exp_f := 0;
        ELSIF x =- 21379 THEN
            exp_f := 0;
        ELSIF x =- 21378 THEN
            exp_f := 0;
        ELSIF x =- 21377 THEN
            exp_f := 0;
        ELSIF x =- 21376 THEN
            exp_f := 0;
        ELSIF x =- 21375 THEN
            exp_f := 0;
        ELSIF x =- 21374 THEN
            exp_f := 0;
        ELSIF x =- 21373 THEN
            exp_f := 0;
        ELSIF x =- 21372 THEN
            exp_f := 0;
        ELSIF x =- 21371 THEN
            exp_f := 0;
        ELSIF x =- 21370 THEN
            exp_f := 0;
        ELSIF x =- 21369 THEN
            exp_f := 0;
        ELSIF x =- 21368 THEN
            exp_f := 0;
        ELSIF x =- 21367 THEN
            exp_f := 0;
        ELSIF x =- 21366 THEN
            exp_f := 0;
        ELSIF x =- 21365 THEN
            exp_f := 0;
        ELSIF x =- 21364 THEN
            exp_f := 0;
        ELSIF x =- 21363 THEN
            exp_f := 0;
        ELSIF x =- 21362 THEN
            exp_f := 0;
        ELSIF x =- 21361 THEN
            exp_f := 0;
        ELSIF x =- 21360 THEN
            exp_f := 0;
        ELSIF x =- 21359 THEN
            exp_f := 0;
        ELSIF x =- 21358 THEN
            exp_f := 0;
        ELSIF x =- 21357 THEN
            exp_f := 0;
        ELSIF x =- 21356 THEN
            exp_f := 0;
        ELSIF x =- 21355 THEN
            exp_f := 0;
        ELSIF x =- 21354 THEN
            exp_f := 0;
        ELSIF x =- 21353 THEN
            exp_f := 0;
        ELSIF x =- 21352 THEN
            exp_f := 0;
        ELSIF x =- 21351 THEN
            exp_f := 0;
        ELSIF x =- 21350 THEN
            exp_f := 0;
        ELSIF x =- 21349 THEN
            exp_f := 0;
        ELSIF x =- 21348 THEN
            exp_f := 0;
        ELSIF x =- 21347 THEN
            exp_f := 0;
        ELSIF x =- 21346 THEN
            exp_f := 0;
        ELSIF x =- 21345 THEN
            exp_f := 0;
        ELSIF x =- 21344 THEN
            exp_f := 0;
        ELSIF x =- 21343 THEN
            exp_f := 0;
        ELSIF x =- 21342 THEN
            exp_f := 0;
        ELSIF x =- 21341 THEN
            exp_f := 0;
        ELSIF x =- 21340 THEN
            exp_f := 0;
        ELSIF x =- 21339 THEN
            exp_f := 0;
        ELSIF x =- 21338 THEN
            exp_f := 0;
        ELSIF x =- 21337 THEN
            exp_f := 0;
        ELSIF x =- 21336 THEN
            exp_f := 0;
        ELSIF x =- 21335 THEN
            exp_f := 0;
        ELSIF x =- 21334 THEN
            exp_f := 0;
        ELSIF x =- 21333 THEN
            exp_f := 0;
        ELSIF x =- 21332 THEN
            exp_f := 0;
        ELSIF x =- 21331 THEN
            exp_f := 0;
        ELSIF x =- 21330 THEN
            exp_f := 0;
        ELSIF x =- 21329 THEN
            exp_f := 0;
        ELSIF x =- 21328 THEN
            exp_f := 0;
        ELSIF x =- 21327 THEN
            exp_f := 0;
        ELSIF x =- 21326 THEN
            exp_f := 0;
        ELSIF x =- 21325 THEN
            exp_f := 0;
        ELSIF x =- 21324 THEN
            exp_f := 0;
        ELSIF x =- 21323 THEN
            exp_f := 0;
        ELSIF x =- 21322 THEN
            exp_f := 0;
        ELSIF x =- 21321 THEN
            exp_f := 0;
        ELSIF x =- 21320 THEN
            exp_f := 0;
        ELSIF x =- 21319 THEN
            exp_f := 0;
        ELSIF x =- 21318 THEN
            exp_f := 0;
        ELSIF x =- 21317 THEN
            exp_f := 0;
        ELSIF x =- 21316 THEN
            exp_f := 0;
        ELSIF x =- 21315 THEN
            exp_f := 0;
        ELSIF x =- 21314 THEN
            exp_f := 0;
        ELSIF x =- 21313 THEN
            exp_f := 0;
        ELSIF x =- 21312 THEN
            exp_f := 0;
        ELSIF x =- 21311 THEN
            exp_f := 0;
        ELSIF x =- 21310 THEN
            exp_f := 0;
        ELSIF x =- 21309 THEN
            exp_f := 0;
        ELSIF x =- 21308 THEN
            exp_f := 0;
        ELSIF x =- 21307 THEN
            exp_f := 0;
        ELSIF x =- 21306 THEN
            exp_f := 0;
        ELSIF x =- 21305 THEN
            exp_f := 0;
        ELSIF x =- 21304 THEN
            exp_f := 0;
        ELSIF x =- 21303 THEN
            exp_f := 0;
        ELSIF x =- 21302 THEN
            exp_f := 0;
        ELSIF x =- 21301 THEN
            exp_f := 0;
        ELSIF x =- 21300 THEN
            exp_f := 0;
        ELSIF x =- 21299 THEN
            exp_f := 0;
        ELSIF x =- 21298 THEN
            exp_f := 0;
        ELSIF x =- 21297 THEN
            exp_f := 0;
        ELSIF x =- 21296 THEN
            exp_f := 0;
        ELSIF x =- 21295 THEN
            exp_f := 0;
        ELSIF x =- 21294 THEN
            exp_f := 0;
        ELSIF x =- 21293 THEN
            exp_f := 0;
        ELSIF x =- 21292 THEN
            exp_f := 0;
        ELSIF x =- 21291 THEN
            exp_f := 0;
        ELSIF x =- 21290 THEN
            exp_f := 0;
        ELSIF x =- 21289 THEN
            exp_f := 0;
        ELSIF x =- 21288 THEN
            exp_f := 0;
        ELSIF x =- 21287 THEN
            exp_f := 0;
        ELSIF x =- 21286 THEN
            exp_f := 0;
        ELSIF x =- 21285 THEN
            exp_f := 0;
        ELSIF x =- 21284 THEN
            exp_f := 0;
        ELSIF x =- 21283 THEN
            exp_f := 0;
        ELSIF x =- 21282 THEN
            exp_f := 0;
        ELSIF x =- 21281 THEN
            exp_f := 0;
        ELSIF x =- 21280 THEN
            exp_f := 0;
        ELSIF x =- 21279 THEN
            exp_f := 0;
        ELSIF x =- 21278 THEN
            exp_f := 0;
        ELSIF x =- 21277 THEN
            exp_f := 0;
        ELSIF x =- 21276 THEN
            exp_f := 0;
        ELSIF x =- 21275 THEN
            exp_f := 0;
        ELSIF x =- 21274 THEN
            exp_f := 0;
        ELSIF x =- 21273 THEN
            exp_f := 0;
        ELSIF x =- 21272 THEN
            exp_f := 0;
        ELSIF x =- 21271 THEN
            exp_f := 0;
        ELSIF x =- 21270 THEN
            exp_f := 0;
        ELSIF x =- 21269 THEN
            exp_f := 0;
        ELSIF x =- 21268 THEN
            exp_f := 0;
        ELSIF x =- 21267 THEN
            exp_f := 0;
        ELSIF x =- 21266 THEN
            exp_f := 0;
        ELSIF x =- 21265 THEN
            exp_f := 0;
        ELSIF x =- 21264 THEN
            exp_f := 0;
        ELSIF x =- 21263 THEN
            exp_f := 0;
        ELSIF x =- 21262 THEN
            exp_f := 0;
        ELSIF x =- 21261 THEN
            exp_f := 0;
        ELSIF x =- 21260 THEN
            exp_f := 0;
        ELSIF x =- 21259 THEN
            exp_f := 0;
        ELSIF x =- 21258 THEN
            exp_f := 0;
        ELSIF x =- 21257 THEN
            exp_f := 0;
        ELSIF x =- 21256 THEN
            exp_f := 0;
        ELSIF x =- 21255 THEN
            exp_f := 0;
        ELSIF x =- 21254 THEN
            exp_f := 0;
        ELSIF x =- 21253 THEN
            exp_f := 0;
        ELSIF x =- 21252 THEN
            exp_f := 0;
        ELSIF x =- 21251 THEN
            exp_f := 0;
        ELSIF x =- 21250 THEN
            exp_f := 0;
        ELSIF x =- 21249 THEN
            exp_f := 0;
        ELSIF x =- 21248 THEN
            exp_f := 0;
        ELSIF x =- 21247 THEN
            exp_f := 0;
        ELSIF x =- 21246 THEN
            exp_f := 0;
        ELSIF x =- 21245 THEN
            exp_f := 0;
        ELSIF x =- 21244 THEN
            exp_f := 0;
        ELSIF x =- 21243 THEN
            exp_f := 0;
        ELSIF x =- 21242 THEN
            exp_f := 0;
        ELSIF x =- 21241 THEN
            exp_f := 0;
        ELSIF x =- 21240 THEN
            exp_f := 0;
        ELSIF x =- 21239 THEN
            exp_f := 0;
        ELSIF x =- 21238 THEN
            exp_f := 0;
        ELSIF x =- 21237 THEN
            exp_f := 0;
        ELSIF x =- 21236 THEN
            exp_f := 0;
        ELSIF x =- 21235 THEN
            exp_f := 0;
        ELSIF x =- 21234 THEN
            exp_f := 0;
        ELSIF x =- 21233 THEN
            exp_f := 0;
        ELSIF x =- 21232 THEN
            exp_f := 0;
        ELSIF x =- 21231 THEN
            exp_f := 0;
        ELSIF x =- 21230 THEN
            exp_f := 0;
        ELSIF x =- 21229 THEN
            exp_f := 0;
        ELSIF x =- 21228 THEN
            exp_f := 0;
        ELSIF x =- 21227 THEN
            exp_f := 0;
        ELSIF x =- 21226 THEN
            exp_f := 0;
        ELSIF x =- 21225 THEN
            exp_f := 0;
        ELSIF x =- 21224 THEN
            exp_f := 0;
        ELSIF x =- 21223 THEN
            exp_f := 0;
        ELSIF x =- 21222 THEN
            exp_f := 0;
        ELSIF x =- 21221 THEN
            exp_f := 0;
        ELSIF x =- 21220 THEN
            exp_f := 0;
        ELSIF x =- 21219 THEN
            exp_f := 0;
        ELSIF x =- 21218 THEN
            exp_f := 0;
        ELSIF x =- 21217 THEN
            exp_f := 0;
        ELSIF x =- 21216 THEN
            exp_f := 0;
        ELSIF x =- 21215 THEN
            exp_f := 0;
        ELSIF x =- 21214 THEN
            exp_f := 0;
        ELSIF x =- 21213 THEN
            exp_f := 0;
        ELSIF x =- 21212 THEN
            exp_f := 0;
        ELSIF x =- 21211 THEN
            exp_f := 0;
        ELSIF x =- 21210 THEN
            exp_f := 0;
        ELSIF x =- 21209 THEN
            exp_f := 0;
        ELSIF x =- 21208 THEN
            exp_f := 0;
        ELSIF x =- 21207 THEN
            exp_f := 0;
        ELSIF x =- 21206 THEN
            exp_f := 0;
        ELSIF x =- 21205 THEN
            exp_f := 0;
        ELSIF x =- 21204 THEN
            exp_f := 0;
        ELSIF x =- 21203 THEN
            exp_f := 0;
        ELSIF x =- 21202 THEN
            exp_f := 0;
        ELSIF x =- 21201 THEN
            exp_f := 0;
        ELSIF x =- 21200 THEN
            exp_f := 0;
        ELSIF x =- 21199 THEN
            exp_f := 0;
        ELSIF x =- 21198 THEN
            exp_f := 0;
        ELSIF x =- 21197 THEN
            exp_f := 0;
        ELSIF x =- 21196 THEN
            exp_f := 0;
        ELSIF x =- 21195 THEN
            exp_f := 0;
        ELSIF x =- 21194 THEN
            exp_f := 0;
        ELSIF x =- 21193 THEN
            exp_f := 0;
        ELSIF x =- 21192 THEN
            exp_f := 0;
        ELSIF x =- 21191 THEN
            exp_f := 0;
        ELSIF x =- 21190 THEN
            exp_f := 0;
        ELSIF x =- 21189 THEN
            exp_f := 0;
        ELSIF x =- 21188 THEN
            exp_f := 0;
        ELSIF x =- 21187 THEN
            exp_f := 0;
        ELSIF x =- 21186 THEN
            exp_f := 0;
        ELSIF x =- 21185 THEN
            exp_f := 0;
        ELSIF x =- 21184 THEN
            exp_f := 0;
        ELSIF x =- 21183 THEN
            exp_f := 0;
        ELSIF x =- 21182 THEN
            exp_f := 0;
        ELSIF x =- 21181 THEN
            exp_f := 0;
        ELSIF x =- 21180 THEN
            exp_f := 0;
        ELSIF x =- 21179 THEN
            exp_f := 0;
        ELSIF x =- 21178 THEN
            exp_f := 0;
        ELSIF x =- 21177 THEN
            exp_f := 0;
        ELSIF x =- 21176 THEN
            exp_f := 0;
        ELSIF x =- 21175 THEN
            exp_f := 0;
        ELSIF x =- 21174 THEN
            exp_f := 0;
        ELSIF x =- 21173 THEN
            exp_f := 0;
        ELSIF x =- 21172 THEN
            exp_f := 0;
        ELSIF x =- 21171 THEN
            exp_f := 0;
        ELSIF x =- 21170 THEN
            exp_f := 0;
        ELSIF x =- 21169 THEN
            exp_f := 0;
        ELSIF x =- 21168 THEN
            exp_f := 0;
        ELSIF x =- 21167 THEN
            exp_f := 0;
        ELSIF x =- 21166 THEN
            exp_f := 0;
        ELSIF x =- 21165 THEN
            exp_f := 0;
        ELSIF x =- 21164 THEN
            exp_f := 0;
        ELSIF x =- 21163 THEN
            exp_f := 0;
        ELSIF x =- 21162 THEN
            exp_f := 0;
        ELSIF x =- 21161 THEN
            exp_f := 0;
        ELSIF x =- 21160 THEN
            exp_f := 0;
        ELSIF x =- 21159 THEN
            exp_f := 0;
        ELSIF x =- 21158 THEN
            exp_f := 0;
        ELSIF x =- 21157 THEN
            exp_f := 0;
        ELSIF x =- 21156 THEN
            exp_f := 0;
        ELSIF x =- 21155 THEN
            exp_f := 0;
        ELSIF x =- 21154 THEN
            exp_f := 0;
        ELSIF x =- 21153 THEN
            exp_f := 0;
        ELSIF x =- 21152 THEN
            exp_f := 0;
        ELSIF x =- 21151 THEN
            exp_f := 0;
        ELSIF x =- 21150 THEN
            exp_f := 0;
        ELSIF x =- 21149 THEN
            exp_f := 0;
        ELSIF x =- 21148 THEN
            exp_f := 0;
        ELSIF x =- 21147 THEN
            exp_f := 0;
        ELSIF x =- 21146 THEN
            exp_f := 0;
        ELSIF x =- 21145 THEN
            exp_f := 0;
        ELSIF x =- 21144 THEN
            exp_f := 0;
        ELSIF x =- 21143 THEN
            exp_f := 0;
        ELSIF x =- 21142 THEN
            exp_f := 0;
        ELSIF x =- 21141 THEN
            exp_f := 0;
        ELSIF x =- 21140 THEN
            exp_f := 0;
        ELSIF x =- 21139 THEN
            exp_f := 0;
        ELSIF x =- 21138 THEN
            exp_f := 0;
        ELSIF x =- 21137 THEN
            exp_f := 0;
        ELSIF x =- 21136 THEN
            exp_f := 0;
        ELSIF x =- 21135 THEN
            exp_f := 0;
        ELSIF x =- 21134 THEN
            exp_f := 0;
        ELSIF x =- 21133 THEN
            exp_f := 0;
        ELSIF x =- 21132 THEN
            exp_f := 0;
        ELSIF x =- 21131 THEN
            exp_f := 0;
        ELSIF x =- 21130 THEN
            exp_f := 0;
        ELSIF x =- 21129 THEN
            exp_f := 0;
        ELSIF x =- 21128 THEN
            exp_f := 0;
        ELSIF x =- 21127 THEN
            exp_f := 0;
        ELSIF x =- 21126 THEN
            exp_f := 0;
        ELSIF x =- 21125 THEN
            exp_f := 0;
        ELSIF x =- 21124 THEN
            exp_f := 0;
        ELSIF x =- 21123 THEN
            exp_f := 0;
        ELSIF x =- 21122 THEN
            exp_f := 0;
        ELSIF x =- 21121 THEN
            exp_f := 0;
        ELSIF x =- 21120 THEN
            exp_f := 0;
        ELSIF x =- 21119 THEN
            exp_f := 0;
        ELSIF x =- 21118 THEN
            exp_f := 0;
        ELSIF x =- 21117 THEN
            exp_f := 0;
        ELSIF x =- 21116 THEN
            exp_f := 0;
        ELSIF x =- 21115 THEN
            exp_f := 0;
        ELSIF x =- 21114 THEN
            exp_f := 0;
        ELSIF x =- 21113 THEN
            exp_f := 0;
        ELSIF x =- 21112 THEN
            exp_f := 0;
        ELSIF x =- 21111 THEN
            exp_f := 0;
        ELSIF x =- 21110 THEN
            exp_f := 0;
        ELSIF x =- 21109 THEN
            exp_f := 0;
        ELSIF x =- 21108 THEN
            exp_f := 0;
        ELSIF x =- 21107 THEN
            exp_f := 0;
        ELSIF x =- 21106 THEN
            exp_f := 0;
        ELSIF x =- 21105 THEN
            exp_f := 0;
        ELSIF x =- 21104 THEN
            exp_f := 0;
        ELSIF x =- 21103 THEN
            exp_f := 0;
        ELSIF x =- 21102 THEN
            exp_f := 0;
        ELSIF x =- 21101 THEN
            exp_f := 0;
        ELSIF x =- 21100 THEN
            exp_f := 0;
        ELSIF x =- 21099 THEN
            exp_f := 0;
        ELSIF x =- 21098 THEN
            exp_f := 0;
        ELSIF x =- 21097 THEN
            exp_f := 0;
        ELSIF x =- 21096 THEN
            exp_f := 0;
        ELSIF x =- 21095 THEN
            exp_f := 0;
        ELSIF x =- 21094 THEN
            exp_f := 0;
        ELSIF x =- 21093 THEN
            exp_f := 0;
        ELSIF x =- 21092 THEN
            exp_f := 0;
        ELSIF x =- 21091 THEN
            exp_f := 0;
        ELSIF x =- 21090 THEN
            exp_f := 0;
        ELSIF x =- 21089 THEN
            exp_f := 0;
        ELSIF x =- 21088 THEN
            exp_f := 0;
        ELSIF x =- 21087 THEN
            exp_f := 0;
        ELSIF x =- 21086 THEN
            exp_f := 0;
        ELSIF x =- 21085 THEN
            exp_f := 0;
        ELSIF x =- 21084 THEN
            exp_f := 0;
        ELSIF x =- 21083 THEN
            exp_f := 0;
        ELSIF x =- 21082 THEN
            exp_f := 0;
        ELSIF x =- 21081 THEN
            exp_f := 0;
        ELSIF x =- 21080 THEN
            exp_f := 0;
        ELSIF x =- 21079 THEN
            exp_f := 0;
        ELSIF x =- 21078 THEN
            exp_f := 0;
        ELSIF x =- 21077 THEN
            exp_f := 0;
        ELSIF x =- 21076 THEN
            exp_f := 0;
        ELSIF x =- 21075 THEN
            exp_f := 0;
        ELSIF x =- 21074 THEN
            exp_f := 0;
        ELSIF x =- 21073 THEN
            exp_f := 0;
        ELSIF x =- 21072 THEN
            exp_f := 0;
        ELSIF x =- 21071 THEN
            exp_f := 0;
        ELSIF x =- 21070 THEN
            exp_f := 0;
        ELSIF x =- 21069 THEN
            exp_f := 0;
        ELSIF x =- 21068 THEN
            exp_f := 0;
        ELSIF x =- 21067 THEN
            exp_f := 0;
        ELSIF x =- 21066 THEN
            exp_f := 0;
        ELSIF x =- 21065 THEN
            exp_f := 0;
        ELSIF x =- 21064 THEN
            exp_f := 0;
        ELSIF x =- 21063 THEN
            exp_f := 0;
        ELSIF x =- 21062 THEN
            exp_f := 0;
        ELSIF x =- 21061 THEN
            exp_f := 0;
        ELSIF x =- 21060 THEN
            exp_f := 0;
        ELSIF x =- 21059 THEN
            exp_f := 0;
        ELSIF x =- 21058 THEN
            exp_f := 0;
        ELSIF x =- 21057 THEN
            exp_f := 0;
        ELSIF x =- 21056 THEN
            exp_f := 0;
        ELSIF x =- 21055 THEN
            exp_f := 0;
        ELSIF x =- 21054 THEN
            exp_f := 0;
        ELSIF x =- 21053 THEN
            exp_f := 0;
        ELSIF x =- 21052 THEN
            exp_f := 0;
        ELSIF x =- 21051 THEN
            exp_f := 0;
        ELSIF x =- 21050 THEN
            exp_f := 0;
        ELSIF x =- 21049 THEN
            exp_f := 0;
        ELSIF x =- 21048 THEN
            exp_f := 0;
        ELSIF x =- 21047 THEN
            exp_f := 0;
        ELSIF x =- 21046 THEN
            exp_f := 0;
        ELSIF x =- 21045 THEN
            exp_f := 0;
        ELSIF x =- 21044 THEN
            exp_f := 0;
        ELSIF x =- 21043 THEN
            exp_f := 0;
        ELSIF x =- 21042 THEN
            exp_f := 0;
        ELSIF x =- 21041 THEN
            exp_f := 0;
        ELSIF x =- 21040 THEN
            exp_f := 0;
        ELSIF x =- 21039 THEN
            exp_f := 0;
        ELSIF x =- 21038 THEN
            exp_f := 0;
        ELSIF x =- 21037 THEN
            exp_f := 0;
        ELSIF x =- 21036 THEN
            exp_f := 0;
        ELSIF x =- 21035 THEN
            exp_f := 0;
        ELSIF x =- 21034 THEN
            exp_f := 0;
        ELSIF x =- 21033 THEN
            exp_f := 0;
        ELSIF x =- 21032 THEN
            exp_f := 0;
        ELSIF x =- 21031 THEN
            exp_f := 0;
        ELSIF x =- 21030 THEN
            exp_f := 0;
        ELSIF x =- 21029 THEN
            exp_f := 0;
        ELSIF x =- 21028 THEN
            exp_f := 0;
        ELSIF x =- 21027 THEN
            exp_f := 0;
        ELSIF x =- 21026 THEN
            exp_f := 0;
        ELSIF x =- 21025 THEN
            exp_f := 0;
        ELSIF x =- 21024 THEN
            exp_f := 0;
        ELSIF x =- 21023 THEN
            exp_f := 0;
        ELSIF x =- 21022 THEN
            exp_f := 0;
        ELSIF x =- 21021 THEN
            exp_f := 0;
        ELSIF x =- 21020 THEN
            exp_f := 0;
        ELSIF x =- 21019 THEN
            exp_f := 0;
        ELSIF x =- 21018 THEN
            exp_f := 0;
        ELSIF x =- 21017 THEN
            exp_f := 0;
        ELSIF x =- 21016 THEN
            exp_f := 0;
        ELSIF x =- 21015 THEN
            exp_f := 0;
        ELSIF x =- 21014 THEN
            exp_f := 0;
        ELSIF x =- 21013 THEN
            exp_f := 0;
        ELSIF x =- 21012 THEN
            exp_f := 0;
        ELSIF x =- 21011 THEN
            exp_f := 0;
        ELSIF x =- 21010 THEN
            exp_f := 0;
        ELSIF x =- 21009 THEN
            exp_f := 0;
        ELSIF x =- 21008 THEN
            exp_f := 0;
        ELSIF x =- 21007 THEN
            exp_f := 0;
        ELSIF x =- 21006 THEN
            exp_f := 0;
        ELSIF x =- 21005 THEN
            exp_f := 0;
        ELSIF x =- 21004 THEN
            exp_f := 0;
        ELSIF x =- 21003 THEN
            exp_f := 0;
        ELSIF x =- 21002 THEN
            exp_f := 0;
        ELSIF x =- 21001 THEN
            exp_f := 0;
        ELSIF x =- 21000 THEN
            exp_f := 0;
        ELSIF x =- 20999 THEN
            exp_f := 0;
        ELSIF x =- 20998 THEN
            exp_f := 0;
        ELSIF x =- 20997 THEN
            exp_f := 0;
        ELSIF x =- 20996 THEN
            exp_f := 0;
        ELSIF x =- 20995 THEN
            exp_f := 0;
        ELSIF x =- 20994 THEN
            exp_f := 0;
        ELSIF x =- 20993 THEN
            exp_f := 0;
        ELSIF x =- 20992 THEN
            exp_f := 0;
        ELSIF x =- 20991 THEN
            exp_f := 0;
        ELSIF x =- 20990 THEN
            exp_f := 0;
        ELSIF x =- 20989 THEN
            exp_f := 0;
        ELSIF x =- 20988 THEN
            exp_f := 0;
        ELSIF x =- 20987 THEN
            exp_f := 0;
        ELSIF x =- 20986 THEN
            exp_f := 0;
        ELSIF x =- 20985 THEN
            exp_f := 0;
        ELSIF x =- 20984 THEN
            exp_f := 0;
        ELSIF x =- 20983 THEN
            exp_f := 0;
        ELSIF x =- 20982 THEN
            exp_f := 0;
        ELSIF x =- 20981 THEN
            exp_f := 0;
        ELSIF x =- 20980 THEN
            exp_f := 0;
        ELSIF x =- 20979 THEN
            exp_f := 0;
        ELSIF x =- 20978 THEN
            exp_f := 0;
        ELSIF x =- 20977 THEN
            exp_f := 0;
        ELSIF x =- 20976 THEN
            exp_f := 0;
        ELSIF x =- 20975 THEN
            exp_f := 0;
        ELSIF x =- 20974 THEN
            exp_f := 0;
        ELSIF x =- 20973 THEN
            exp_f := 0;
        ELSIF x =- 20972 THEN
            exp_f := 0;
        ELSIF x =- 20971 THEN
            exp_f := 0;
        ELSIF x =- 20970 THEN
            exp_f := 0;
        ELSIF x =- 20969 THEN
            exp_f := 0;
        ELSIF x =- 20968 THEN
            exp_f := 0;
        ELSIF x =- 20967 THEN
            exp_f := 0;
        ELSIF x =- 20966 THEN
            exp_f := 0;
        ELSIF x =- 20965 THEN
            exp_f := 0;
        ELSIF x =- 20964 THEN
            exp_f := 0;
        ELSIF x =- 20963 THEN
            exp_f := 0;
        ELSIF x =- 20962 THEN
            exp_f := 0;
        ELSIF x =- 20961 THEN
            exp_f := 0;
        ELSIF x =- 20960 THEN
            exp_f := 0;
        ELSIF x =- 20959 THEN
            exp_f := 0;
        ELSIF x =- 20958 THEN
            exp_f := 0;
        ELSIF x =- 20957 THEN
            exp_f := 0;
        ELSIF x =- 20956 THEN
            exp_f := 0;
        ELSIF x =- 20955 THEN
            exp_f := 0;
        ELSIF x =- 20954 THEN
            exp_f := 0;
        ELSIF x =- 20953 THEN
            exp_f := 0;
        ELSIF x =- 20952 THEN
            exp_f := 0;
        ELSIF x =- 20951 THEN
            exp_f := 0;
        ELSIF x =- 20950 THEN
            exp_f := 0;
        ELSIF x =- 20949 THEN
            exp_f := 0;
        ELSIF x =- 20948 THEN
            exp_f := 0;
        ELSIF x =- 20947 THEN
            exp_f := 0;
        ELSIF x =- 20946 THEN
            exp_f := 0;
        ELSIF x =- 20945 THEN
            exp_f := 0;
        ELSIF x =- 20944 THEN
            exp_f := 0;
        ELSIF x =- 20943 THEN
            exp_f := 0;
        ELSIF x =- 20942 THEN
            exp_f := 0;
        ELSIF x =- 20941 THEN
            exp_f := 0;
        ELSIF x =- 20940 THEN
            exp_f := 0;
        ELSIF x =- 20939 THEN
            exp_f := 0;
        ELSIF x =- 20938 THEN
            exp_f := 0;
        ELSIF x =- 20937 THEN
            exp_f := 0;
        ELSIF x =- 20936 THEN
            exp_f := 0;
        ELSIF x =- 20935 THEN
            exp_f := 0;
        ELSIF x =- 20934 THEN
            exp_f := 0;
        ELSIF x =- 20933 THEN
            exp_f := 0;
        ELSIF x =- 20932 THEN
            exp_f := 0;
        ELSIF x =- 20931 THEN
            exp_f := 0;
        ELSIF x =- 20930 THEN
            exp_f := 0;
        ELSIF x =- 20929 THEN
            exp_f := 0;
        ELSIF x =- 20928 THEN
            exp_f := 0;
        ELSIF x =- 20927 THEN
            exp_f := 0;
        ELSIF x =- 20926 THEN
            exp_f := 0;
        ELSIF x =- 20925 THEN
            exp_f := 0;
        ELSIF x =- 20924 THEN
            exp_f := 0;
        ELSIF x =- 20923 THEN
            exp_f := 0;
        ELSIF x =- 20922 THEN
            exp_f := 0;
        ELSIF x =- 20921 THEN
            exp_f := 0;
        ELSIF x =- 20920 THEN
            exp_f := 0;
        ELSIF x =- 20919 THEN
            exp_f := 0;
        ELSIF x =- 20918 THEN
            exp_f := 0;
        ELSIF x =- 20917 THEN
            exp_f := 0;
        ELSIF x =- 20916 THEN
            exp_f := 0;
        ELSIF x =- 20915 THEN
            exp_f := 0;
        ELSIF x =- 20914 THEN
            exp_f := 0;
        ELSIF x =- 20913 THEN
            exp_f := 0;
        ELSIF x =- 20912 THEN
            exp_f := 0;
        ELSIF x =- 20911 THEN
            exp_f := 0;
        ELSIF x =- 20910 THEN
            exp_f := 0;
        ELSIF x =- 20909 THEN
            exp_f := 0;
        ELSIF x =- 20908 THEN
            exp_f := 0;
        ELSIF x =- 20907 THEN
            exp_f := 0;
        ELSIF x =- 20906 THEN
            exp_f := 0;
        ELSIF x =- 20905 THEN
            exp_f := 0;
        ELSIF x =- 20904 THEN
            exp_f := 0;
        ELSIF x =- 20903 THEN
            exp_f := 0;
        ELSIF x =- 20902 THEN
            exp_f := 0;
        ELSIF x =- 20901 THEN
            exp_f := 0;
        ELSIF x =- 20900 THEN
            exp_f := 0;
        ELSIF x =- 20899 THEN
            exp_f := 0;
        ELSIF x =- 20898 THEN
            exp_f := 0;
        ELSIF x =- 20897 THEN
            exp_f := 0;
        ELSIF x =- 20896 THEN
            exp_f := 0;
        ELSIF x =- 20895 THEN
            exp_f := 0;
        ELSIF x =- 20894 THEN
            exp_f := 0;
        ELSIF x =- 20893 THEN
            exp_f := 0;
        ELSIF x =- 20892 THEN
            exp_f := 0;
        ELSIF x =- 20891 THEN
            exp_f := 0;
        ELSIF x =- 20890 THEN
            exp_f := 0;
        ELSIF x =- 20889 THEN
            exp_f := 0;
        ELSIF x =- 20888 THEN
            exp_f := 0;
        ELSIF x =- 20887 THEN
            exp_f := 0;
        ELSIF x =- 20886 THEN
            exp_f := 0;
        ELSIF x =- 20885 THEN
            exp_f := 0;
        ELSIF x =- 20884 THEN
            exp_f := 0;
        ELSIF x =- 20883 THEN
            exp_f := 0;
        ELSIF x =- 20882 THEN
            exp_f := 0;
        ELSIF x =- 20881 THEN
            exp_f := 0;
        ELSIF x =- 20880 THEN
            exp_f := 0;
        ELSIF x =- 20879 THEN
            exp_f := 0;
        ELSIF x =- 20878 THEN
            exp_f := 0;
        ELSIF x =- 20877 THEN
            exp_f := 0;
        ELSIF x =- 20876 THEN
            exp_f := 0;
        ELSIF x =- 20875 THEN
            exp_f := 0;
        ELSIF x =- 20874 THEN
            exp_f := 0;
        ELSIF x =- 20873 THEN
            exp_f := 0;
        ELSIF x =- 20872 THEN
            exp_f := 0;
        ELSIF x =- 20871 THEN
            exp_f := 0;
        ELSIF x =- 20870 THEN
            exp_f := 0;
        ELSIF x =- 20869 THEN
            exp_f := 0;
        ELSIF x =- 20868 THEN
            exp_f := 0;
        ELSIF x =- 20867 THEN
            exp_f := 0;
        ELSIF x =- 20866 THEN
            exp_f := 0;
        ELSIF x =- 20865 THEN
            exp_f := 0;
        ELSIF x =- 20864 THEN
            exp_f := 0;
        ELSIF x =- 20863 THEN
            exp_f := 0;
        ELSIF x =- 20862 THEN
            exp_f := 0;
        ELSIF x =- 20861 THEN
            exp_f := 0;
        ELSIF x =- 20860 THEN
            exp_f := 0;
        ELSIF x =- 20859 THEN
            exp_f := 0;
        ELSIF x =- 20858 THEN
            exp_f := 0;
        ELSIF x =- 20857 THEN
            exp_f := 0;
        ELSIF x =- 20856 THEN
            exp_f := 0;
        ELSIF x =- 20855 THEN
            exp_f := 0;
        ELSIF x =- 20854 THEN
            exp_f := 0;
        ELSIF x =- 20853 THEN
            exp_f := 0;
        ELSIF x =- 20852 THEN
            exp_f := 0;
        ELSIF x =- 20851 THEN
            exp_f := 0;
        ELSIF x =- 20850 THEN
            exp_f := 0;
        ELSIF x =- 20849 THEN
            exp_f := 0;
        ELSIF x =- 20848 THEN
            exp_f := 0;
        ELSIF x =- 20847 THEN
            exp_f := 0;
        ELSIF x =- 20846 THEN
            exp_f := 0;
        ELSIF x =- 20845 THEN
            exp_f := 0;
        ELSIF x =- 20844 THEN
            exp_f := 0;
        ELSIF x =- 20843 THEN
            exp_f := 0;
        ELSIF x =- 20842 THEN
            exp_f := 0;
        ELSIF x =- 20841 THEN
            exp_f := 0;
        ELSIF x =- 20840 THEN
            exp_f := 0;
        ELSIF x =- 20839 THEN
            exp_f := 0;
        ELSIF x =- 20838 THEN
            exp_f := 0;
        ELSIF x =- 20837 THEN
            exp_f := 0;
        ELSIF x =- 20836 THEN
            exp_f := 0;
        ELSIF x =- 20835 THEN
            exp_f := 0;
        ELSIF x =- 20834 THEN
            exp_f := 0;
        ELSIF x =- 20833 THEN
            exp_f := 0;
        ELSIF x =- 20832 THEN
            exp_f := 0;
        ELSIF x =- 20831 THEN
            exp_f := 0;
        ELSIF x =- 20830 THEN
            exp_f := 0;
        ELSIF x =- 20829 THEN
            exp_f := 0;
        ELSIF x =- 20828 THEN
            exp_f := 0;
        ELSIF x =- 20827 THEN
            exp_f := 0;
        ELSIF x =- 20826 THEN
            exp_f := 0;
        ELSIF x =- 20825 THEN
            exp_f := 0;
        ELSIF x =- 20824 THEN
            exp_f := 0;
        ELSIF x =- 20823 THEN
            exp_f := 0;
        ELSIF x =- 20822 THEN
            exp_f := 0;
        ELSIF x =- 20821 THEN
            exp_f := 0;
        ELSIF x =- 20820 THEN
            exp_f := 0;
        ELSIF x =- 20819 THEN
            exp_f := 0;
        ELSIF x =- 20818 THEN
            exp_f := 0;
        ELSIF x =- 20817 THEN
            exp_f := 0;
        ELSIF x =- 20816 THEN
            exp_f := 0;
        ELSIF x =- 20815 THEN
            exp_f := 0;
        ELSIF x =- 20814 THEN
            exp_f := 0;
        ELSIF x =- 20813 THEN
            exp_f := 0;
        ELSIF x =- 20812 THEN
            exp_f := 0;
        ELSIF x =- 20811 THEN
            exp_f := 0;
        ELSIF x =- 20810 THEN
            exp_f := 0;
        ELSIF x =- 20809 THEN
            exp_f := 0;
        ELSIF x =- 20808 THEN
            exp_f := 0;
        ELSIF x =- 20807 THEN
            exp_f := 0;
        ELSIF x =- 20806 THEN
            exp_f := 0;
        ELSIF x =- 20805 THEN
            exp_f := 0;
        ELSIF x =- 20804 THEN
            exp_f := 0;
        ELSIF x =- 20803 THEN
            exp_f := 0;
        ELSIF x =- 20802 THEN
            exp_f := 0;
        ELSIF x =- 20801 THEN
            exp_f := 0;
        ELSIF x =- 20800 THEN
            exp_f := 0;
        ELSIF x =- 20799 THEN
            exp_f := 0;
        ELSIF x =- 20798 THEN
            exp_f := 0;
        ELSIF x =- 20797 THEN
            exp_f := 0;
        ELSIF x =- 20796 THEN
            exp_f := 0;
        ELSIF x =- 20795 THEN
            exp_f := 0;
        ELSIF x =- 20794 THEN
            exp_f := 0;
        ELSIF x =- 20793 THEN
            exp_f := 0;
        ELSIF x =- 20792 THEN
            exp_f := 0;
        ELSIF x =- 20791 THEN
            exp_f := 0;
        ELSIF x =- 20790 THEN
            exp_f := 0;
        ELSIF x =- 20789 THEN
            exp_f := 0;
        ELSIF x =- 20788 THEN
            exp_f := 0;
        ELSIF x =- 20787 THEN
            exp_f := 0;
        ELSIF x =- 20786 THEN
            exp_f := 0;
        ELSIF x =- 20785 THEN
            exp_f := 0;
        ELSIF x =- 20784 THEN
            exp_f := 0;
        ELSIF x =- 20783 THEN
            exp_f := 0;
        ELSIF x =- 20782 THEN
            exp_f := 0;
        ELSIF x =- 20781 THEN
            exp_f := 0;
        ELSIF x =- 20780 THEN
            exp_f := 0;
        ELSIF x =- 20779 THEN
            exp_f := 0;
        ELSIF x =- 20778 THEN
            exp_f := 0;
        ELSIF x =- 20777 THEN
            exp_f := 0;
        ELSIF x =- 20776 THEN
            exp_f := 0;
        ELSIF x =- 20775 THEN
            exp_f := 0;
        ELSIF x =- 20774 THEN
            exp_f := 0;
        ELSIF x =- 20773 THEN
            exp_f := 0;
        ELSIF x =- 20772 THEN
            exp_f := 0;
        ELSIF x =- 20771 THEN
            exp_f := 0;
        ELSIF x =- 20770 THEN
            exp_f := 0;
        ELSIF x =- 20769 THEN
            exp_f := 0;
        ELSIF x =- 20768 THEN
            exp_f := 0;
        ELSIF x =- 20767 THEN
            exp_f := 0;
        ELSIF x =- 20766 THEN
            exp_f := 0;
        ELSIF x =- 20765 THEN
            exp_f := 0;
        ELSIF x =- 20764 THEN
            exp_f := 0;
        ELSIF x =- 20763 THEN
            exp_f := 0;
        ELSIF x =- 20762 THEN
            exp_f := 0;
        ELSIF x =- 20761 THEN
            exp_f := 0;
        ELSIF x =- 20760 THEN
            exp_f := 0;
        ELSIF x =- 20759 THEN
            exp_f := 0;
        ELSIF x =- 20758 THEN
            exp_f := 0;
        ELSIF x =- 20757 THEN
            exp_f := 0;
        ELSIF x =- 20756 THEN
            exp_f := 0;
        ELSIF x =- 20755 THEN
            exp_f := 0;
        ELSIF x =- 20754 THEN
            exp_f := 0;
        ELSIF x =- 20753 THEN
            exp_f := 0;
        ELSIF x =- 20752 THEN
            exp_f := 0;
        ELSIF x =- 20751 THEN
            exp_f := 0;
        ELSIF x =- 20750 THEN
            exp_f := 0;
        ELSIF x =- 20749 THEN
            exp_f := 0;
        ELSIF x =- 20748 THEN
            exp_f := 0;
        ELSIF x =- 20747 THEN
            exp_f := 0;
        ELSIF x =- 20746 THEN
            exp_f := 0;
        ELSIF x =- 20745 THEN
            exp_f := 0;
        ELSIF x =- 20744 THEN
            exp_f := 0;
        ELSIF x =- 20743 THEN
            exp_f := 0;
        ELSIF x =- 20742 THEN
            exp_f := 0;
        ELSIF x =- 20741 THEN
            exp_f := 0;
        ELSIF x =- 20740 THEN
            exp_f := 0;
        ELSIF x =- 20739 THEN
            exp_f := 0;
        ELSIF x =- 20738 THEN
            exp_f := 0;
        ELSIF x =- 20737 THEN
            exp_f := 0;
        ELSIF x =- 20736 THEN
            exp_f := 0;
        ELSIF x =- 20735 THEN
            exp_f := 0;
        ELSIF x =- 20734 THEN
            exp_f := 0;
        ELSIF x =- 20733 THEN
            exp_f := 0;
        ELSIF x =- 20732 THEN
            exp_f := 0;
        ELSIF x =- 20731 THEN
            exp_f := 0;
        ELSIF x =- 20730 THEN
            exp_f := 0;
        ELSIF x =- 20729 THEN
            exp_f := 0;
        ELSIF x =- 20728 THEN
            exp_f := 0;
        ELSIF x =- 20727 THEN
            exp_f := 0;
        ELSIF x =- 20726 THEN
            exp_f := 0;
        ELSIF x =- 20725 THEN
            exp_f := 0;
        ELSIF x =- 20724 THEN
            exp_f := 0;
        ELSIF x =- 20723 THEN
            exp_f := 0;
        ELSIF x =- 20722 THEN
            exp_f := 0;
        ELSIF x =- 20721 THEN
            exp_f := 0;
        ELSIF x =- 20720 THEN
            exp_f := 0;
        ELSIF x =- 20719 THEN
            exp_f := 0;
        ELSIF x =- 20718 THEN
            exp_f := 0;
        ELSIF x =- 20717 THEN
            exp_f := 0;
        ELSIF x =- 20716 THEN
            exp_f := 0;
        ELSIF x =- 20715 THEN
            exp_f := 0;
        ELSIF x =- 20714 THEN
            exp_f := 0;
        ELSIF x =- 20713 THEN
            exp_f := 0;
        ELSIF x =- 20712 THEN
            exp_f := 0;
        ELSIF x =- 20711 THEN
            exp_f := 0;
        ELSIF x =- 20710 THEN
            exp_f := 0;
        ELSIF x =- 20709 THEN
            exp_f := 0;
        ELSIF x =- 20708 THEN
            exp_f := 0;
        ELSIF x =- 20707 THEN
            exp_f := 0;
        ELSIF x =- 20706 THEN
            exp_f := 0;
        ELSIF x =- 20705 THEN
            exp_f := 0;
        ELSIF x =- 20704 THEN
            exp_f := 0;
        ELSIF x =- 20703 THEN
            exp_f := 0;
        ELSIF x =- 20702 THEN
            exp_f := 0;
        ELSIF x =- 20701 THEN
            exp_f := 0;
        ELSIF x =- 20700 THEN
            exp_f := 0;
        ELSIF x =- 20699 THEN
            exp_f := 0;
        ELSIF x =- 20698 THEN
            exp_f := 0;
        ELSIF x =- 20697 THEN
            exp_f := 0;
        ELSIF x =- 20696 THEN
            exp_f := 0;
        ELSIF x =- 20695 THEN
            exp_f := 0;
        ELSIF x =- 20694 THEN
            exp_f := 0;
        ELSIF x =- 20693 THEN
            exp_f := 0;
        ELSIF x =- 20692 THEN
            exp_f := 0;
        ELSIF x =- 20691 THEN
            exp_f := 0;
        ELSIF x =- 20690 THEN
            exp_f := 0;
        ELSIF x =- 20689 THEN
            exp_f := 0;
        ELSIF x =- 20688 THEN
            exp_f := 0;
        ELSIF x =- 20687 THEN
            exp_f := 0;
        ELSIF x =- 20686 THEN
            exp_f := 0;
        ELSIF x =- 20685 THEN
            exp_f := 0;
        ELSIF x =- 20684 THEN
            exp_f := 0;
        ELSIF x =- 20683 THEN
            exp_f := 0;
        ELSIF x =- 20682 THEN
            exp_f := 0;
        ELSIF x =- 20681 THEN
            exp_f := 0;
        ELSIF x =- 20680 THEN
            exp_f := 0;
        ELSIF x =- 20679 THEN
            exp_f := 0;
        ELSIF x =- 20678 THEN
            exp_f := 0;
        ELSIF x =- 20677 THEN
            exp_f := 0;
        ELSIF x =- 20676 THEN
            exp_f := 0;
        ELSIF x =- 20675 THEN
            exp_f := 0;
        ELSIF x =- 20674 THEN
            exp_f := 0;
        ELSIF x =- 20673 THEN
            exp_f := 0;
        ELSIF x =- 20672 THEN
            exp_f := 0;
        ELSIF x =- 20671 THEN
            exp_f := 0;
        ELSIF x =- 20670 THEN
            exp_f := 0;
        ELSIF x =- 20669 THEN
            exp_f := 0;
        ELSIF x =- 20668 THEN
            exp_f := 0;
        ELSIF x =- 20667 THEN
            exp_f := 0;
        ELSIF x =- 20666 THEN
            exp_f := 0;
        ELSIF x =- 20665 THEN
            exp_f := 0;
        ELSIF x =- 20664 THEN
            exp_f := 0;
        ELSIF x =- 20663 THEN
            exp_f := 0;
        ELSIF x =- 20662 THEN
            exp_f := 0;
        ELSIF x =- 20661 THEN
            exp_f := 0;
        ELSIF x =- 20660 THEN
            exp_f := 0;
        ELSIF x =- 20659 THEN
            exp_f := 0;
        ELSIF x =- 20658 THEN
            exp_f := 0;
        ELSIF x =- 20657 THEN
            exp_f := 0;
        ELSIF x =- 20656 THEN
            exp_f := 0;
        ELSIF x =- 20655 THEN
            exp_f := 0;
        ELSIF x =- 20654 THEN
            exp_f := 0;
        ELSIF x =- 20653 THEN
            exp_f := 0;
        ELSIF x =- 20652 THEN
            exp_f := 0;
        ELSIF x =- 20651 THEN
            exp_f := 0;
        ELSIF x =- 20650 THEN
            exp_f := 0;
        ELSIF x =- 20649 THEN
            exp_f := 0;
        ELSIF x =- 20648 THEN
            exp_f := 0;
        ELSIF x =- 20647 THEN
            exp_f := 0;
        ELSIF x =- 20646 THEN
            exp_f := 0;
        ELSIF x =- 20645 THEN
            exp_f := 0;
        ELSIF x =- 20644 THEN
            exp_f := 0;
        ELSIF x =- 20643 THEN
            exp_f := 0;
        ELSIF x =- 20642 THEN
            exp_f := 0;
        ELSIF x =- 20641 THEN
            exp_f := 0;
        ELSIF x =- 20640 THEN
            exp_f := 0;
        ELSIF x =- 20639 THEN
            exp_f := 0;
        ELSIF x =- 20638 THEN
            exp_f := 0;
        ELSIF x =- 20637 THEN
            exp_f := 0;
        ELSIF x =- 20636 THEN
            exp_f := 0;
        ELSIF x =- 20635 THEN
            exp_f := 0;
        ELSIF x =- 20634 THEN
            exp_f := 0;
        ELSIF x =- 20633 THEN
            exp_f := 0;
        ELSIF x =- 20632 THEN
            exp_f := 0;
        ELSIF x =- 20631 THEN
            exp_f := 0;
        ELSIF x =- 20630 THEN
            exp_f := 0;
        ELSIF x =- 20629 THEN
            exp_f := 0;
        ELSIF x =- 20628 THEN
            exp_f := 0;
        ELSIF x =- 20627 THEN
            exp_f := 0;
        ELSIF x =- 20626 THEN
            exp_f := 0;
        ELSIF x =- 20625 THEN
            exp_f := 0;
        ELSIF x =- 20624 THEN
            exp_f := 0;
        ELSIF x =- 20623 THEN
            exp_f := 0;
        ELSIF x =- 20622 THEN
            exp_f := 0;
        ELSIF x =- 20621 THEN
            exp_f := 0;
        ELSIF x =- 20620 THEN
            exp_f := 0;
        ELSIF x =- 20619 THEN
            exp_f := 0;
        ELSIF x =- 20618 THEN
            exp_f := 0;
        ELSIF x =- 20617 THEN
            exp_f := 0;
        ELSIF x =- 20616 THEN
            exp_f := 0;
        ELSIF x =- 20615 THEN
            exp_f := 0;
        ELSIF x =- 20614 THEN
            exp_f := 0;
        ELSIF x =- 20613 THEN
            exp_f := 0;
        ELSIF x =- 20612 THEN
            exp_f := 0;
        ELSIF x =- 20611 THEN
            exp_f := 0;
        ELSIF x =- 20610 THEN
            exp_f := 0;
        ELSIF x =- 20609 THEN
            exp_f := 0;
        ELSIF x =- 20608 THEN
            exp_f := 0;
        ELSIF x =- 20607 THEN
            exp_f := 0;
        ELSIF x =- 20606 THEN
            exp_f := 0;
        ELSIF x =- 20605 THEN
            exp_f := 0;
        ELSIF x =- 20604 THEN
            exp_f := 0;
        ELSIF x =- 20603 THEN
            exp_f := 0;
        ELSIF x =- 20602 THEN
            exp_f := 0;
        ELSIF x =- 20601 THEN
            exp_f := 0;
        ELSIF x =- 20600 THEN
            exp_f := 0;
        ELSIF x =- 20599 THEN
            exp_f := 0;
        ELSIF x =- 20598 THEN
            exp_f := 0;
        ELSIF x =- 20597 THEN
            exp_f := 0;
        ELSIF x =- 20596 THEN
            exp_f := 0;
        ELSIF x =- 20595 THEN
            exp_f := 0;
        ELSIF x =- 20594 THEN
            exp_f := 0;
        ELSIF x =- 20593 THEN
            exp_f := 0;
        ELSIF x =- 20592 THEN
            exp_f := 0;
        ELSIF x =- 20591 THEN
            exp_f := 0;
        ELSIF x =- 20590 THEN
            exp_f := 0;
        ELSIF x =- 20589 THEN
            exp_f := 0;
        ELSIF x =- 20588 THEN
            exp_f := 0;
        ELSIF x =- 20587 THEN
            exp_f := 0;
        ELSIF x =- 20586 THEN
            exp_f := 0;
        ELSIF x =- 20585 THEN
            exp_f := 0;
        ELSIF x =- 20584 THEN
            exp_f := 0;
        ELSIF x =- 20583 THEN
            exp_f := 0;
        ELSIF x =- 20582 THEN
            exp_f := 0;
        ELSIF x =- 20581 THEN
            exp_f := 0;
        ELSIF x =- 20580 THEN
            exp_f := 0;
        ELSIF x =- 20579 THEN
            exp_f := 0;
        ELSIF x =- 20578 THEN
            exp_f := 0;
        ELSIF x =- 20577 THEN
            exp_f := 0;
        ELSIF x =- 20576 THEN
            exp_f := 0;
        ELSIF x =- 20575 THEN
            exp_f := 0;
        ELSIF x =- 20574 THEN
            exp_f := 0;
        ELSIF x =- 20573 THEN
            exp_f := 0;
        ELSIF x =- 20572 THEN
            exp_f := 0;
        ELSIF x =- 20571 THEN
            exp_f := 0;
        ELSIF x =- 20570 THEN
            exp_f := 0;
        ELSIF x =- 20569 THEN
            exp_f := 0;
        ELSIF x =- 20568 THEN
            exp_f := 0;
        ELSIF x =- 20567 THEN
            exp_f := 0;
        ELSIF x =- 20566 THEN
            exp_f := 0;
        ELSIF x =- 20565 THEN
            exp_f := 0;
        ELSIF x =- 20564 THEN
            exp_f := 0;
        ELSIF x =- 20563 THEN
            exp_f := 0;
        ELSIF x =- 20562 THEN
            exp_f := 0;
        ELSIF x =- 20561 THEN
            exp_f := 0;
        ELSIF x =- 20560 THEN
            exp_f := 0;
        ELSIF x =- 20559 THEN
            exp_f := 0;
        ELSIF x =- 20558 THEN
            exp_f := 0;
        ELSIF x =- 20557 THEN
            exp_f := 0;
        ELSIF x =- 20556 THEN
            exp_f := 0;
        ELSIF x =- 20555 THEN
            exp_f := 0;
        ELSIF x =- 20554 THEN
            exp_f := 0;
        ELSIF x =- 20553 THEN
            exp_f := 0;
        ELSIF x =- 20552 THEN
            exp_f := 0;
        ELSIF x =- 20551 THEN
            exp_f := 0;
        ELSIF x =- 20550 THEN
            exp_f := 0;
        ELSIF x =- 20549 THEN
            exp_f := 0;
        ELSIF x =- 20548 THEN
            exp_f := 0;
        ELSIF x =- 20547 THEN
            exp_f := 0;
        ELSIF x =- 20546 THEN
            exp_f := 0;
        ELSIF x =- 20545 THEN
            exp_f := 0;
        ELSIF x =- 20544 THEN
            exp_f := 0;
        ELSIF x =- 20543 THEN
            exp_f := 0;
        ELSIF x =- 20542 THEN
            exp_f := 0;
        ELSIF x =- 20541 THEN
            exp_f := 0;
        ELSIF x =- 20540 THEN
            exp_f := 0;
        ELSIF x =- 20539 THEN
            exp_f := 0;
        ELSIF x =- 20538 THEN
            exp_f := 0;
        ELSIF x =- 20537 THEN
            exp_f := 0;
        ELSIF x =- 20536 THEN
            exp_f := 0;
        ELSIF x =- 20535 THEN
            exp_f := 0;
        ELSIF x =- 20534 THEN
            exp_f := 0;
        ELSIF x =- 20533 THEN
            exp_f := 0;
        ELSIF x =- 20532 THEN
            exp_f := 0;
        ELSIF x =- 20531 THEN
            exp_f := 0;
        ELSIF x =- 20530 THEN
            exp_f := 0;
        ELSIF x =- 20529 THEN
            exp_f := 0;
        ELSIF x =- 20528 THEN
            exp_f := 0;
        ELSIF x =- 20527 THEN
            exp_f := 0;
        ELSIF x =- 20526 THEN
            exp_f := 0;
        ELSIF x =- 20525 THEN
            exp_f := 0;
        ELSIF x =- 20524 THEN
            exp_f := 0;
        ELSIF x =- 20523 THEN
            exp_f := 0;
        ELSIF x =- 20522 THEN
            exp_f := 0;
        ELSIF x =- 20521 THEN
            exp_f := 0;
        ELSIF x =- 20520 THEN
            exp_f := 0;
        ELSIF x =- 20519 THEN
            exp_f := 0;
        ELSIF x =- 20518 THEN
            exp_f := 0;
        ELSIF x =- 20517 THEN
            exp_f := 0;
        ELSIF x =- 20516 THEN
            exp_f := 0;
        ELSIF x =- 20515 THEN
            exp_f := 0;
        ELSIF x =- 20514 THEN
            exp_f := 0;
        ELSIF x =- 20513 THEN
            exp_f := 0;
        ELSIF x =- 20512 THEN
            exp_f := 0;
        ELSIF x =- 20511 THEN
            exp_f := 0;
        ELSIF x =- 20510 THEN
            exp_f := 0;
        ELSIF x =- 20509 THEN
            exp_f := 0;
        ELSIF x =- 20508 THEN
            exp_f := 0;
        ELSIF x =- 20507 THEN
            exp_f := 0;
        ELSIF x =- 20506 THEN
            exp_f := 0;
        ELSIF x =- 20505 THEN
            exp_f := 0;
        ELSIF x =- 20504 THEN
            exp_f := 0;
        ELSIF x =- 20503 THEN
            exp_f := 0;
        ELSIF x =- 20502 THEN
            exp_f := 0;
        ELSIF x =- 20501 THEN
            exp_f := 0;
        ELSIF x =- 20500 THEN
            exp_f := 0;
        ELSIF x =- 20499 THEN
            exp_f := 0;
        ELSIF x =- 20498 THEN
            exp_f := 0;
        ELSIF x =- 20497 THEN
            exp_f := 0;
        ELSIF x =- 20496 THEN
            exp_f := 0;
        ELSIF x =- 20495 THEN
            exp_f := 0;
        ELSIF x =- 20494 THEN
            exp_f := 0;
        ELSIF x =- 20493 THEN
            exp_f := 0;
        ELSIF x =- 20492 THEN
            exp_f := 0;
        ELSIF x =- 20491 THEN
            exp_f := 0;
        ELSIF x =- 20490 THEN
            exp_f := 0;
        ELSIF x =- 20489 THEN
            exp_f := 0;
        ELSIF x =- 20488 THEN
            exp_f := 0;
        ELSIF x =- 20487 THEN
            exp_f := 0;
        ELSIF x =- 20486 THEN
            exp_f := 0;
        ELSIF x =- 20485 THEN
            exp_f := 0;
        ELSIF x =- 20484 THEN
            exp_f := 0;
        ELSIF x =- 20483 THEN
            exp_f := 0;
        ELSIF x =- 20482 THEN
            exp_f := 0;
        ELSIF x =- 20481 THEN
            exp_f := 0;
        ELSIF x =- 20480 THEN
            exp_f := 0;
        ELSIF x =- 20479 THEN
            exp_f := 0;
        ELSIF x =- 20478 THEN
            exp_f := 0;
        ELSIF x =- 20477 THEN
            exp_f := 0;
        ELSIF x =- 20476 THEN
            exp_f := 0;
        ELSIF x =- 20475 THEN
            exp_f := 0;
        ELSIF x =- 20474 THEN
            exp_f := 0;
        ELSIF x =- 20473 THEN
            exp_f := 0;
        ELSIF x =- 20472 THEN
            exp_f := 0;
        ELSIF x =- 20471 THEN
            exp_f := 0;
        ELSIF x =- 20470 THEN
            exp_f := 0;
        ELSIF x =- 20469 THEN
            exp_f := 0;
        ELSIF x =- 20468 THEN
            exp_f := 0;
        ELSIF x =- 20467 THEN
            exp_f := 0;
        ELSIF x =- 20466 THEN
            exp_f := 0;
        ELSIF x =- 20465 THEN
            exp_f := 0;
        ELSIF x =- 20464 THEN
            exp_f := 0;
        ELSIF x =- 20463 THEN
            exp_f := 0;
        ELSIF x =- 20462 THEN
            exp_f := 0;
        ELSIF x =- 20461 THEN
            exp_f := 0;
        ELSIF x =- 20460 THEN
            exp_f := 0;
        ELSIF x =- 20459 THEN
            exp_f := 0;
        ELSIF x =- 20458 THEN
            exp_f := 0;
        ELSIF x =- 20457 THEN
            exp_f := 0;
        ELSIF x =- 20456 THEN
            exp_f := 0;
        ELSIF x =- 20455 THEN
            exp_f := 0;
        ELSIF x =- 20454 THEN
            exp_f := 0;
        ELSIF x =- 20453 THEN
            exp_f := 0;
        ELSIF x =- 20452 THEN
            exp_f := 0;
        ELSIF x =- 20451 THEN
            exp_f := 0;
        ELSIF x =- 20450 THEN
            exp_f := 0;
        ELSIF x =- 20449 THEN
            exp_f := 0;
        ELSIF x =- 20448 THEN
            exp_f := 0;
        ELSIF x =- 20447 THEN
            exp_f := 0;
        ELSIF x =- 20446 THEN
            exp_f := 0;
        ELSIF x =- 20445 THEN
            exp_f := 0;
        ELSIF x =- 20444 THEN
            exp_f := 0;
        ELSIF x =- 20443 THEN
            exp_f := 0;
        ELSIF x =- 20442 THEN
            exp_f := 0;
        ELSIF x =- 20441 THEN
            exp_f := 0;
        ELSIF x =- 20440 THEN
            exp_f := 0;
        ELSIF x =- 20439 THEN
            exp_f := 0;
        ELSIF x =- 20438 THEN
            exp_f := 0;
        ELSIF x =- 20437 THEN
            exp_f := 0;
        ELSIF x =- 20436 THEN
            exp_f := 0;
        ELSIF x =- 20435 THEN
            exp_f := 0;
        ELSIF x =- 20434 THEN
            exp_f := 0;
        ELSIF x =- 20433 THEN
            exp_f := 0;
        ELSIF x =- 20432 THEN
            exp_f := 0;
        ELSIF x =- 20431 THEN
            exp_f := 0;
        ELSIF x =- 20430 THEN
            exp_f := 0;
        ELSIF x =- 20429 THEN
            exp_f := 0;
        ELSIF x =- 20428 THEN
            exp_f := 0;
        ELSIF x =- 20427 THEN
            exp_f := 0;
        ELSIF x =- 20426 THEN
            exp_f := 0;
        ELSIF x =- 20425 THEN
            exp_f := 0;
        ELSIF x =- 20424 THEN
            exp_f := 0;
        ELSIF x =- 20423 THEN
            exp_f := 0;
        ELSIF x =- 20422 THEN
            exp_f := 0;
        ELSIF x =- 20421 THEN
            exp_f := 0;
        ELSIF x =- 20420 THEN
            exp_f := 0;
        ELSIF x =- 20419 THEN
            exp_f := 0;
        ELSIF x =- 20418 THEN
            exp_f := 0;
        ELSIF x =- 20417 THEN
            exp_f := 0;
        ELSIF x =- 20416 THEN
            exp_f := 0;
        ELSIF x =- 20415 THEN
            exp_f := 0;
        ELSIF x =- 20414 THEN
            exp_f := 0;
        ELSIF x =- 20413 THEN
            exp_f := 0;
        ELSIF x =- 20412 THEN
            exp_f := 0;
        ELSIF x =- 20411 THEN
            exp_f := 0;
        ELSIF x =- 20410 THEN
            exp_f := 0;
        ELSIF x =- 20409 THEN
            exp_f := 0;
        ELSIF x =- 20408 THEN
            exp_f := 0;
        ELSIF x =- 20407 THEN
            exp_f := 0;
        ELSIF x =- 20406 THEN
            exp_f := 0;
        ELSIF x =- 20405 THEN
            exp_f := 0;
        ELSIF x =- 20404 THEN
            exp_f := 0;
        ELSIF x =- 20403 THEN
            exp_f := 0;
        ELSIF x =- 20402 THEN
            exp_f := 0;
        ELSIF x =- 20401 THEN
            exp_f := 0;
        ELSIF x =- 20400 THEN
            exp_f := 0;
        ELSIF x =- 20399 THEN
            exp_f := 0;
        ELSIF x =- 20398 THEN
            exp_f := 0;
        ELSIF x =- 20397 THEN
            exp_f := 0;
        ELSIF x =- 20396 THEN
            exp_f := 0;
        ELSIF x =- 20395 THEN
            exp_f := 0;
        ELSIF x =- 20394 THEN
            exp_f := 0;
        ELSIF x =- 20393 THEN
            exp_f := 0;
        ELSIF x =- 20392 THEN
            exp_f := 0;
        ELSIF x =- 20391 THEN
            exp_f := 0;
        ELSIF x =- 20390 THEN
            exp_f := 0;
        ELSIF x =- 20389 THEN
            exp_f := 0;
        ELSIF x =- 20388 THEN
            exp_f := 0;
        ELSIF x =- 20387 THEN
            exp_f := 0;
        ELSIF x =- 20386 THEN
            exp_f := 0;
        ELSIF x =- 20385 THEN
            exp_f := 0;
        ELSIF x =- 20384 THEN
            exp_f := 0;
        ELSIF x =- 20383 THEN
            exp_f := 0;
        ELSIF x =- 20382 THEN
            exp_f := 0;
        ELSIF x =- 20381 THEN
            exp_f := 0;
        ELSIF x =- 20380 THEN
            exp_f := 0;
        ELSIF x =- 20379 THEN
            exp_f := 0;
        ELSIF x =- 20378 THEN
            exp_f := 0;
        ELSIF x =- 20377 THEN
            exp_f := 0;
        ELSIF x =- 20376 THEN
            exp_f := 0;
        ELSIF x =- 20375 THEN
            exp_f := 0;
        ELSIF x =- 20374 THEN
            exp_f := 0;
        ELSIF x =- 20373 THEN
            exp_f := 0;
        ELSIF x =- 20372 THEN
            exp_f := 0;
        ELSIF x =- 20371 THEN
            exp_f := 0;
        ELSIF x =- 20370 THEN
            exp_f := 0;
        ELSIF x =- 20369 THEN
            exp_f := 0;
        ELSIF x =- 20368 THEN
            exp_f := 0;
        ELSIF x =- 20367 THEN
            exp_f := 0;
        ELSIF x =- 20366 THEN
            exp_f := 0;
        ELSIF x =- 20365 THEN
            exp_f := 0;
        ELSIF x =- 20364 THEN
            exp_f := 0;
        ELSIF x =- 20363 THEN
            exp_f := 0;
        ELSIF x =- 20362 THEN
            exp_f := 0;
        ELSIF x =- 20361 THEN
            exp_f := 0;
        ELSIF x =- 20360 THEN
            exp_f := 0;
        ELSIF x =- 20359 THEN
            exp_f := 0;
        ELSIF x =- 20358 THEN
            exp_f := 0;
        ELSIF x =- 20357 THEN
            exp_f := 0;
        ELSIF x =- 20356 THEN
            exp_f := 0;
        ELSIF x =- 20355 THEN
            exp_f := 0;
        ELSIF x =- 20354 THEN
            exp_f := 0;
        ELSIF x =- 20353 THEN
            exp_f := 0;
        ELSIF x =- 20352 THEN
            exp_f := 0;
        ELSIF x =- 20351 THEN
            exp_f := 0;
        ELSIF x =- 20350 THEN
            exp_f := 0;
        ELSIF x =- 20349 THEN
            exp_f := 0;
        ELSIF x =- 20348 THEN
            exp_f := 0;
        ELSIF x =- 20347 THEN
            exp_f := 0;
        ELSIF x =- 20346 THEN
            exp_f := 0;
        ELSIF x =- 20345 THEN
            exp_f := 0;
        ELSIF x =- 20344 THEN
            exp_f := 0;
        ELSIF x =- 20343 THEN
            exp_f := 0;
        ELSIF x =- 20342 THEN
            exp_f := 0;
        ELSIF x =- 20341 THEN
            exp_f := 0;
        ELSIF x =- 20340 THEN
            exp_f := 0;
        ELSIF x =- 20339 THEN
            exp_f := 0;
        ELSIF x =- 20338 THEN
            exp_f := 0;
        ELSIF x =- 20337 THEN
            exp_f := 0;
        ELSIF x =- 20336 THEN
            exp_f := 0;
        ELSIF x =- 20335 THEN
            exp_f := 0;
        ELSIF x =- 20334 THEN
            exp_f := 0;
        ELSIF x =- 20333 THEN
            exp_f := 0;
        ELSIF x =- 20332 THEN
            exp_f := 0;
        ELSIF x =- 20331 THEN
            exp_f := 0;
        ELSIF x =- 20330 THEN
            exp_f := 0;
        ELSIF x =- 20329 THEN
            exp_f := 0;
        ELSIF x =- 20328 THEN
            exp_f := 0;
        ELSIF x =- 20327 THEN
            exp_f := 0;
        ELSIF x =- 20326 THEN
            exp_f := 0;
        ELSIF x =- 20325 THEN
            exp_f := 0;
        ELSIF x =- 20324 THEN
            exp_f := 0;
        ELSIF x =- 20323 THEN
            exp_f := 0;
        ELSIF x =- 20322 THEN
            exp_f := 0;
        ELSIF x =- 20321 THEN
            exp_f := 0;
        ELSIF x =- 20320 THEN
            exp_f := 0;
        ELSIF x =- 20319 THEN
            exp_f := 0;
        ELSIF x =- 20318 THEN
            exp_f := 0;
        ELSIF x =- 20317 THEN
            exp_f := 0;
        ELSIF x =- 20316 THEN
            exp_f := 0;
        ELSIF x =- 20315 THEN
            exp_f := 0;
        ELSIF x =- 20314 THEN
            exp_f := 0;
        ELSIF x =- 20313 THEN
            exp_f := 0;
        ELSIF x =- 20312 THEN
            exp_f := 0;
        ELSIF x =- 20311 THEN
            exp_f := 0;
        ELSIF x =- 20310 THEN
            exp_f := 0;
        ELSIF x =- 20309 THEN
            exp_f := 0;
        ELSIF x =- 20308 THEN
            exp_f := 0;
        ELSIF x =- 20307 THEN
            exp_f := 0;
        ELSIF x =- 20306 THEN
            exp_f := 0;
        ELSIF x =- 20305 THEN
            exp_f := 0;
        ELSIF x =- 20304 THEN
            exp_f := 0;
        ELSIF x =- 20303 THEN
            exp_f := 0;
        ELSIF x =- 20302 THEN
            exp_f := 0;
        ELSIF x =- 20301 THEN
            exp_f := 0;
        ELSIF x =- 20300 THEN
            exp_f := 0;
        ELSIF x =- 20299 THEN
            exp_f := 0;
        ELSIF x =- 20298 THEN
            exp_f := 0;
        ELSIF x =- 20297 THEN
            exp_f := 0;
        ELSIF x =- 20296 THEN
            exp_f := 0;
        ELSIF x =- 20295 THEN
            exp_f := 0;
        ELSIF x =- 20294 THEN
            exp_f := 0;
        ELSIF x =- 20293 THEN
            exp_f := 0;
        ELSIF x =- 20292 THEN
            exp_f := 0;
        ELSIF x =- 20291 THEN
            exp_f := 0;
        ELSIF x =- 20290 THEN
            exp_f := 0;
        ELSIF x =- 20289 THEN
            exp_f := 0;
        ELSIF x =- 20288 THEN
            exp_f := 0;
        ELSIF x =- 20287 THEN
            exp_f := 0;
        ELSIF x =- 20286 THEN
            exp_f := 0;
        ELSIF x =- 20285 THEN
            exp_f := 0;
        ELSIF x =- 20284 THEN
            exp_f := 0;
        ELSIF x =- 20283 THEN
            exp_f := 0;
        ELSIF x =- 20282 THEN
            exp_f := 0;
        ELSIF x =- 20281 THEN
            exp_f := 0;
        ELSIF x =- 20280 THEN
            exp_f := 0;
        ELSIF x =- 20279 THEN
            exp_f := 0;
        ELSIF x =- 20278 THEN
            exp_f := 0;
        ELSIF x =- 20277 THEN
            exp_f := 0;
        ELSIF x =- 20276 THEN
            exp_f := 0;
        ELSIF x =- 20275 THEN
            exp_f := 0;
        ELSIF x =- 20274 THEN
            exp_f := 0;
        ELSIF x =- 20273 THEN
            exp_f := 0;
        ELSIF x =- 20272 THEN
            exp_f := 0;
        ELSIF x =- 20271 THEN
            exp_f := 0;
        ELSIF x =- 20270 THEN
            exp_f := 0;
        ELSIF x =- 20269 THEN
            exp_f := 0;
        ELSIF x =- 20268 THEN
            exp_f := 0;
        ELSIF x =- 20267 THEN
            exp_f := 0;
        ELSIF x =- 20266 THEN
            exp_f := 0;
        ELSIF x =- 20265 THEN
            exp_f := 0;
        ELSIF x =- 20264 THEN
            exp_f := 0;
        ELSIF x =- 20263 THEN
            exp_f := 0;
        ELSIF x =- 20262 THEN
            exp_f := 0;
        ELSIF x =- 20261 THEN
            exp_f := 0;
        ELSIF x =- 20260 THEN
            exp_f := 0;
        ELSIF x =- 20259 THEN
            exp_f := 0;
        ELSIF x =- 20258 THEN
            exp_f := 0;
        ELSIF x =- 20257 THEN
            exp_f := 0;
        ELSIF x =- 20256 THEN
            exp_f := 0;
        ELSIF x =- 20255 THEN
            exp_f := 0;
        ELSIF x =- 20254 THEN
            exp_f := 0;
        ELSIF x =- 20253 THEN
            exp_f := 0;
        ELSIF x =- 20252 THEN
            exp_f := 0;
        ELSIF x =- 20251 THEN
            exp_f := 0;
        ELSIF x =- 20250 THEN
            exp_f := 0;
        ELSIF x =- 20249 THEN
            exp_f := 0;
        ELSIF x =- 20248 THEN
            exp_f := 0;
        ELSIF x =- 20247 THEN
            exp_f := 0;
        ELSIF x =- 20246 THEN
            exp_f := 0;
        ELSIF x =- 20245 THEN
            exp_f := 0;
        ELSIF x =- 20244 THEN
            exp_f := 0;
        ELSIF x =- 20243 THEN
            exp_f := 0;
        ELSIF x =- 20242 THEN
            exp_f := 0;
        ELSIF x =- 20241 THEN
            exp_f := 0;
        ELSIF x =- 20240 THEN
            exp_f := 0;
        ELSIF x =- 20239 THEN
            exp_f := 0;
        ELSIF x =- 20238 THEN
            exp_f := 0;
        ELSIF x =- 20237 THEN
            exp_f := 0;
        ELSIF x =- 20236 THEN
            exp_f := 0;
        ELSIF x =- 20235 THEN
            exp_f := 0;
        ELSIF x =- 20234 THEN
            exp_f := 0;
        ELSIF x =- 20233 THEN
            exp_f := 0;
        ELSIF x =- 20232 THEN
            exp_f := 0;
        ELSIF x =- 20231 THEN
            exp_f := 0;
        ELSIF x =- 20230 THEN
            exp_f := 0;
        ELSIF x =- 20229 THEN
            exp_f := 0;
        ELSIF x =- 20228 THEN
            exp_f := 0;
        ELSIF x =- 20227 THEN
            exp_f := 0;
        ELSIF x =- 20226 THEN
            exp_f := 0;
        ELSIF x =- 20225 THEN
            exp_f := 0;
        ELSIF x =- 20224 THEN
            exp_f := 0;
        ELSIF x =- 20223 THEN
            exp_f := 0;
        ELSIF x =- 20222 THEN
            exp_f := 0;
        ELSIF x =- 20221 THEN
            exp_f := 0;
        ELSIF x =- 20220 THEN
            exp_f := 0;
        ELSIF x =- 20219 THEN
            exp_f := 0;
        ELSIF x =- 20218 THEN
            exp_f := 0;
        ELSIF x =- 20217 THEN
            exp_f := 0;
        ELSIF x =- 20216 THEN
            exp_f := 0;
        ELSIF x =- 20215 THEN
            exp_f := 0;
        ELSIF x =- 20214 THEN
            exp_f := 0;
        ELSIF x =- 20213 THEN
            exp_f := 0;
        ELSIF x =- 20212 THEN
            exp_f := 0;
        ELSIF x =- 20211 THEN
            exp_f := 0;
        ELSIF x =- 20210 THEN
            exp_f := 0;
        ELSIF x =- 20209 THEN
            exp_f := 0;
        ELSIF x =- 20208 THEN
            exp_f := 0;
        ELSIF x =- 20207 THEN
            exp_f := 0;
        ELSIF x =- 20206 THEN
            exp_f := 0;
        ELSIF x =- 20205 THEN
            exp_f := 0;
        ELSIF x =- 20204 THEN
            exp_f := 0;
        ELSIF x =- 20203 THEN
            exp_f := 0;
        ELSIF x =- 20202 THEN
            exp_f := 0;
        ELSIF x =- 20201 THEN
            exp_f := 0;
        ELSIF x =- 20200 THEN
            exp_f := 0;
        ELSIF x =- 20199 THEN
            exp_f := 0;
        ELSIF x =- 20198 THEN
            exp_f := 0;
        ELSIF x =- 20197 THEN
            exp_f := 0;
        ELSIF x =- 20196 THEN
            exp_f := 0;
        ELSIF x =- 20195 THEN
            exp_f := 0;
        ELSIF x =- 20194 THEN
            exp_f := 0;
        ELSIF x =- 20193 THEN
            exp_f := 0;
        ELSIF x =- 20192 THEN
            exp_f := 0;
        ELSIF x =- 20191 THEN
            exp_f := 0;
        ELSIF x =- 20190 THEN
            exp_f := 0;
        ELSIF x =- 20189 THEN
            exp_f := 0;
        ELSIF x =- 20188 THEN
            exp_f := 0;
        ELSIF x =- 20187 THEN
            exp_f := 0;
        ELSIF x =- 20186 THEN
            exp_f := 0;
        ELSIF x =- 20185 THEN
            exp_f := 0;
        ELSIF x =- 20184 THEN
            exp_f := 0;
        ELSIF x =- 20183 THEN
            exp_f := 0;
        ELSIF x =- 20182 THEN
            exp_f := 0;
        ELSIF x =- 20181 THEN
            exp_f := 0;
        ELSIF x =- 20180 THEN
            exp_f := 0;
        ELSIF x =- 20179 THEN
            exp_f := 0;
        ELSIF x =- 20178 THEN
            exp_f := 0;
        ELSIF x =- 20177 THEN
            exp_f := 0;
        ELSIF x =- 20176 THEN
            exp_f := 0;
        ELSIF x =- 20175 THEN
            exp_f := 0;
        ELSIF x =- 20174 THEN
            exp_f := 0;
        ELSIF x =- 20173 THEN
            exp_f := 0;
        ELSIF x =- 20172 THEN
            exp_f := 0;
        ELSIF x =- 20171 THEN
            exp_f := 0;
        ELSIF x =- 20170 THEN
            exp_f := 0;
        ELSIF x =- 20169 THEN
            exp_f := 0;
        ELSIF x =- 20168 THEN
            exp_f := 0;
        ELSIF x =- 20167 THEN
            exp_f := 0;
        ELSIF x =- 20166 THEN
            exp_f := 0;
        ELSIF x =- 20165 THEN
            exp_f := 0;
        ELSIF x =- 20164 THEN
            exp_f := 0;
        ELSIF x =- 20163 THEN
            exp_f := 0;
        ELSIF x =- 20162 THEN
            exp_f := 0;
        ELSIF x =- 20161 THEN
            exp_f := 0;
        ELSIF x =- 20160 THEN
            exp_f := 0;
        ELSIF x =- 20159 THEN
            exp_f := 0;
        ELSIF x =- 20158 THEN
            exp_f := 0;
        ELSIF x =- 20157 THEN
            exp_f := 0;
        ELSIF x =- 20156 THEN
            exp_f := 0;
        ELSIF x =- 20155 THEN
            exp_f := 0;
        ELSIF x =- 20154 THEN
            exp_f := 0;
        ELSIF x =- 20153 THEN
            exp_f := 0;
        ELSIF x =- 20152 THEN
            exp_f := 0;
        ELSIF x =- 20151 THEN
            exp_f := 0;
        ELSIF x =- 20150 THEN
            exp_f := 0;
        ELSIF x =- 20149 THEN
            exp_f := 0;
        ELSIF x =- 20148 THEN
            exp_f := 0;
        ELSIF x =- 20147 THEN
            exp_f := 0;
        ELSIF x =- 20146 THEN
            exp_f := 0;
        ELSIF x =- 20145 THEN
            exp_f := 0;
        ELSIF x =- 20144 THEN
            exp_f := 0;
        ELSIF x =- 20143 THEN
            exp_f := 0;
        ELSIF x =- 20142 THEN
            exp_f := 0;
        ELSIF x =- 20141 THEN
            exp_f := 0;
        ELSIF x =- 20140 THEN
            exp_f := 0;
        ELSIF x =- 20139 THEN
            exp_f := 0;
        ELSIF x =- 20138 THEN
            exp_f := 0;
        ELSIF x =- 20137 THEN
            exp_f := 0;
        ELSIF x =- 20136 THEN
            exp_f := 0;
        ELSIF x =- 20135 THEN
            exp_f := 0;
        ELSIF x =- 20134 THEN
            exp_f := 0;
        ELSIF x =- 20133 THEN
            exp_f := 0;
        ELSIF x =- 20132 THEN
            exp_f := 0;
        ELSIF x =- 20131 THEN
            exp_f := 0;
        ELSIF x =- 20130 THEN
            exp_f := 0;
        ELSIF x =- 20129 THEN
            exp_f := 0;
        ELSIF x =- 20128 THEN
            exp_f := 0;
        ELSIF x =- 20127 THEN
            exp_f := 0;
        ELSIF x =- 20126 THEN
            exp_f := 0;
        ELSIF x =- 20125 THEN
            exp_f := 0;
        ELSIF x =- 20124 THEN
            exp_f := 0;
        ELSIF x =- 20123 THEN
            exp_f := 0;
        ELSIF x =- 20122 THEN
            exp_f := 0;
        ELSIF x =- 20121 THEN
            exp_f := 0;
        ELSIF x =- 20120 THEN
            exp_f := 0;
        ELSIF x =- 20119 THEN
            exp_f := 0;
        ELSIF x =- 20118 THEN
            exp_f := 0;
        ELSIF x =- 20117 THEN
            exp_f := 0;
        ELSIF x =- 20116 THEN
            exp_f := 0;
        ELSIF x =- 20115 THEN
            exp_f := 0;
        ELSIF x =- 20114 THEN
            exp_f := 0;
        ELSIF x =- 20113 THEN
            exp_f := 0;
        ELSIF x =- 20112 THEN
            exp_f := 0;
        ELSIF x =- 20111 THEN
            exp_f := 0;
        ELSIF x =- 20110 THEN
            exp_f := 0;
        ELSIF x =- 20109 THEN
            exp_f := 0;
        ELSIF x =- 20108 THEN
            exp_f := 0;
        ELSIF x =- 20107 THEN
            exp_f := 0;
        ELSIF x =- 20106 THEN
            exp_f := 0;
        ELSIF x =- 20105 THEN
            exp_f := 0;
        ELSIF x =- 20104 THEN
            exp_f := 0;
        ELSIF x =- 20103 THEN
            exp_f := 0;
        ELSIF x =- 20102 THEN
            exp_f := 0;
        ELSIF x =- 20101 THEN
            exp_f := 0;
        ELSIF x =- 20100 THEN
            exp_f := 0;
        ELSIF x =- 20099 THEN
            exp_f := 0;
        ELSIF x =- 20098 THEN
            exp_f := 0;
        ELSIF x =- 20097 THEN
            exp_f := 0;
        ELSIF x =- 20096 THEN
            exp_f := 0;
        ELSIF x =- 20095 THEN
            exp_f := 0;
        ELSIF x =- 20094 THEN
            exp_f := 0;
        ELSIF x =- 20093 THEN
            exp_f := 0;
        ELSIF x =- 20092 THEN
            exp_f := 0;
        ELSIF x =- 20091 THEN
            exp_f := 0;
        ELSIF x =- 20090 THEN
            exp_f := 0;
        ELSIF x =- 20089 THEN
            exp_f := 0;
        ELSIF x =- 20088 THEN
            exp_f := 0;
        ELSIF x =- 20087 THEN
            exp_f := 0;
        ELSIF x =- 20086 THEN
            exp_f := 0;
        ELSIF x =- 20085 THEN
            exp_f := 0;
        ELSIF x =- 20084 THEN
            exp_f := 0;
        ELSIF x =- 20083 THEN
            exp_f := 0;
        ELSIF x =- 20082 THEN
            exp_f := 0;
        ELSIF x =- 20081 THEN
            exp_f := 0;
        ELSIF x =- 20080 THEN
            exp_f := 0;
        ELSIF x =- 20079 THEN
            exp_f := 0;
        ELSIF x =- 20078 THEN
            exp_f := 0;
        ELSIF x =- 20077 THEN
            exp_f := 0;
        ELSIF x =- 20076 THEN
            exp_f := 0;
        ELSIF x =- 20075 THEN
            exp_f := 0;
        ELSIF x =- 20074 THEN
            exp_f := 0;
        ELSIF x =- 20073 THEN
            exp_f := 0;
        ELSIF x =- 20072 THEN
            exp_f := 0;
        ELSIF x =- 20071 THEN
            exp_f := 0;
        ELSIF x =- 20070 THEN
            exp_f := 0;
        ELSIF x =- 20069 THEN
            exp_f := 0;
        ELSIF x =- 20068 THEN
            exp_f := 0;
        ELSIF x =- 20067 THEN
            exp_f := 0;
        ELSIF x =- 20066 THEN
            exp_f := 0;
        ELSIF x =- 20065 THEN
            exp_f := 0;
        ELSIF x =- 20064 THEN
            exp_f := 0;
        ELSIF x =- 20063 THEN
            exp_f := 0;
        ELSIF x =- 20062 THEN
            exp_f := 0;
        ELSIF x =- 20061 THEN
            exp_f := 0;
        ELSIF x =- 20060 THEN
            exp_f := 0;
        ELSIF x =- 20059 THEN
            exp_f := 0;
        ELSIF x =- 20058 THEN
            exp_f := 0;
        ELSIF x =- 20057 THEN
            exp_f := 0;
        ELSIF x =- 20056 THEN
            exp_f := 0;
        ELSIF x =- 20055 THEN
            exp_f := 0;
        ELSIF x =- 20054 THEN
            exp_f := 0;
        ELSIF x =- 20053 THEN
            exp_f := 0;
        ELSIF x =- 20052 THEN
            exp_f := 0;
        ELSIF x =- 20051 THEN
            exp_f := 0;
        ELSIF x =- 20050 THEN
            exp_f := 0;
        ELSIF x =- 20049 THEN
            exp_f := 0;
        ELSIF x =- 20048 THEN
            exp_f := 0;
        ELSIF x =- 20047 THEN
            exp_f := 0;
        ELSIF x =- 20046 THEN
            exp_f := 0;
        ELSIF x =- 20045 THEN
            exp_f := 0;
        ELSIF x =- 20044 THEN
            exp_f := 0;
        ELSIF x =- 20043 THEN
            exp_f := 0;
        ELSIF x =- 20042 THEN
            exp_f := 0;
        ELSIF x =- 20041 THEN
            exp_f := 0;
        ELSIF x =- 20040 THEN
            exp_f := 0;
        ELSIF x =- 20039 THEN
            exp_f := 0;
        ELSIF x =- 20038 THEN
            exp_f := 0;
        ELSIF x =- 20037 THEN
            exp_f := 0;
        ELSIF x =- 20036 THEN
            exp_f := 0;
        ELSIF x =- 20035 THEN
            exp_f := 0;
        ELSIF x =- 20034 THEN
            exp_f := 0;
        ELSIF x =- 20033 THEN
            exp_f := 0;
        ELSIF x =- 20032 THEN
            exp_f := 0;
        ELSIF x =- 20031 THEN
            exp_f := 0;
        ELSIF x =- 20030 THEN
            exp_f := 0;
        ELSIF x =- 20029 THEN
            exp_f := 0;
        ELSIF x =- 20028 THEN
            exp_f := 0;
        ELSIF x =- 20027 THEN
            exp_f := 0;
        ELSIF x =- 20026 THEN
            exp_f := 0;
        ELSIF x =- 20025 THEN
            exp_f := 0;
        ELSIF x =- 20024 THEN
            exp_f := 0;
        ELSIF x =- 20023 THEN
            exp_f := 0;
        ELSIF x =- 20022 THEN
            exp_f := 0;
        ELSIF x =- 20021 THEN
            exp_f := 0;
        ELSIF x =- 20020 THEN
            exp_f := 0;
        ELSIF x =- 20019 THEN
            exp_f := 0;
        ELSIF x =- 20018 THEN
            exp_f := 0;
        ELSIF x =- 20017 THEN
            exp_f := 0;
        ELSIF x =- 20016 THEN
            exp_f := 0;
        ELSIF x =- 20015 THEN
            exp_f := 0;
        ELSIF x =- 20014 THEN
            exp_f := 0;
        ELSIF x =- 20013 THEN
            exp_f := 0;
        ELSIF x =- 20012 THEN
            exp_f := 0;
        ELSIF x =- 20011 THEN
            exp_f := 0;
        ELSIF x =- 20010 THEN
            exp_f := 0;
        ELSIF x =- 20009 THEN
            exp_f := 0;
        ELSIF x =- 20008 THEN
            exp_f := 0;
        ELSIF x =- 20007 THEN
            exp_f := 0;
        ELSIF x =- 20006 THEN
            exp_f := 0;
        ELSIF x =- 20005 THEN
            exp_f := 0;
        ELSIF x =- 20004 THEN
            exp_f := 0;
        ELSIF x =- 20003 THEN
            exp_f := 0;
        ELSIF x =- 20002 THEN
            exp_f := 0;
        ELSIF x =- 20001 THEN
            exp_f := 0;
        ELSIF x =- 20000 THEN
            exp_f := 0;
        ELSIF x =- 19999 THEN
            exp_f := 0;
        ELSIF x =- 19998 THEN
            exp_f := 0;
        ELSIF x =- 19997 THEN
            exp_f := 0;
        ELSIF x =- 19996 THEN
            exp_f := 0;
        ELSIF x =- 19995 THEN
            exp_f := 0;
        ELSIF x =- 19994 THEN
            exp_f := 0;
        ELSIF x =- 19993 THEN
            exp_f := 0;
        ELSIF x =- 19992 THEN
            exp_f := 0;
        ELSIF x =- 19991 THEN
            exp_f := 0;
        ELSIF x =- 19990 THEN
            exp_f := 0;
        ELSIF x =- 19989 THEN
            exp_f := 0;
        ELSIF x =- 19988 THEN
            exp_f := 0;
        ELSIF x =- 19987 THEN
            exp_f := 0;
        ELSIF x =- 19986 THEN
            exp_f := 0;
        ELSIF x =- 19985 THEN
            exp_f := 0;
        ELSIF x =- 19984 THEN
            exp_f := 0;
        ELSIF x =- 19983 THEN
            exp_f := 0;
        ELSIF x =- 19982 THEN
            exp_f := 0;
        ELSIF x =- 19981 THEN
            exp_f := 0;
        ELSIF x =- 19980 THEN
            exp_f := 0;
        ELSIF x =- 19979 THEN
            exp_f := 0;
        ELSIF x =- 19978 THEN
            exp_f := 0;
        ELSIF x =- 19977 THEN
            exp_f := 0;
        ELSIF x =- 19976 THEN
            exp_f := 0;
        ELSIF x =- 19975 THEN
            exp_f := 0;
        ELSIF x =- 19974 THEN
            exp_f := 0;
        ELSIF x =- 19973 THEN
            exp_f := 0;
        ELSIF x =- 19972 THEN
            exp_f := 0;
        ELSIF x =- 19971 THEN
            exp_f := 0;
        ELSIF x =- 19970 THEN
            exp_f := 0;
        ELSIF x =- 19969 THEN
            exp_f := 0;
        ELSIF x =- 19968 THEN
            exp_f := 0;
        ELSIF x =- 19967 THEN
            exp_f := 0;
        ELSIF x =- 19966 THEN
            exp_f := 0;
        ELSIF x =- 19965 THEN
            exp_f := 0;
        ELSIF x =- 19964 THEN
            exp_f := 0;
        ELSIF x =- 19963 THEN
            exp_f := 0;
        ELSIF x =- 19962 THEN
            exp_f := 0;
        ELSIF x =- 19961 THEN
            exp_f := 0;
        ELSIF x =- 19960 THEN
            exp_f := 0;
        ELSIF x =- 19959 THEN
            exp_f := 0;
        ELSIF x =- 19958 THEN
            exp_f := 0;
        ELSIF x =- 19957 THEN
            exp_f := 0;
        ELSIF x =- 19956 THEN
            exp_f := 0;
        ELSIF x =- 19955 THEN
            exp_f := 0;
        ELSIF x =- 19954 THEN
            exp_f := 0;
        ELSIF x =- 19953 THEN
            exp_f := 0;
        ELSIF x =- 19952 THEN
            exp_f := 0;
        ELSIF x =- 19951 THEN
            exp_f := 0;
        ELSIF x =- 19950 THEN
            exp_f := 0;
        ELSIF x =- 19949 THEN
            exp_f := 0;
        ELSIF x =- 19948 THEN
            exp_f := 0;
        ELSIF x =- 19947 THEN
            exp_f := 0;
        ELSIF x =- 19946 THEN
            exp_f := 0;
        ELSIF x =- 19945 THEN
            exp_f := 0;
        ELSIF x =- 19944 THEN
            exp_f := 0;
        ELSIF x =- 19943 THEN
            exp_f := 0;
        ELSIF x =- 19942 THEN
            exp_f := 0;
        ELSIF x =- 19941 THEN
            exp_f := 0;
        ELSIF x =- 19940 THEN
            exp_f := 0;
        ELSIF x =- 19939 THEN
            exp_f := 0;
        ELSIF x =- 19938 THEN
            exp_f := 0;
        ELSIF x =- 19937 THEN
            exp_f := 0;
        ELSIF x =- 19936 THEN
            exp_f := 0;
        ELSIF x =- 19935 THEN
            exp_f := 0;
        ELSIF x =- 19934 THEN
            exp_f := 0;
        ELSIF x =- 19933 THEN
            exp_f := 0;
        ELSIF x =- 19932 THEN
            exp_f := 0;
        ELSIF x =- 19931 THEN
            exp_f := 0;
        ELSIF x =- 19930 THEN
            exp_f := 0;
        ELSIF x =- 19929 THEN
            exp_f := 0;
        ELSIF x =- 19928 THEN
            exp_f := 0;
        ELSIF x =- 19927 THEN
            exp_f := 0;
        ELSIF x =- 19926 THEN
            exp_f := 0;
        ELSIF x =- 19925 THEN
            exp_f := 0;
        ELSIF x =- 19924 THEN
            exp_f := 0;
        ELSIF x =- 19923 THEN
            exp_f := 0;
        ELSIF x =- 19922 THEN
            exp_f := 0;
        ELSIF x =- 19921 THEN
            exp_f := 0;
        ELSIF x =- 19920 THEN
            exp_f := 0;
        ELSIF x =- 19919 THEN
            exp_f := 0;
        ELSIF x =- 19918 THEN
            exp_f := 0;
        ELSIF x =- 19917 THEN
            exp_f := 0;
        ELSIF x =- 19916 THEN
            exp_f := 0;
        ELSIF x =- 19915 THEN
            exp_f := 0;
        ELSIF x =- 19914 THEN
            exp_f := 0;
        ELSIF x =- 19913 THEN
            exp_f := 0;
        ELSIF x =- 19912 THEN
            exp_f := 0;
        ELSIF x =- 19911 THEN
            exp_f := 0;
        ELSIF x =- 19910 THEN
            exp_f := 0;
        ELSIF x =- 19909 THEN
            exp_f := 0;
        ELSIF x =- 19908 THEN
            exp_f := 0;
        ELSIF x =- 19907 THEN
            exp_f := 0;
        ELSIF x =- 19906 THEN
            exp_f := 0;
        ELSIF x =- 19905 THEN
            exp_f := 0;
        ELSIF x =- 19904 THEN
            exp_f := 0;
        ELSIF x =- 19903 THEN
            exp_f := 0;
        ELSIF x =- 19902 THEN
            exp_f := 0;
        ELSIF x =- 19901 THEN
            exp_f := 0;
        ELSIF x =- 19900 THEN
            exp_f := 0;
        ELSIF x =- 19899 THEN
            exp_f := 0;
        ELSIF x =- 19898 THEN
            exp_f := 0;
        ELSIF x =- 19897 THEN
            exp_f := 0;
        ELSIF x =- 19896 THEN
            exp_f := 0;
        ELSIF x =- 19895 THEN
            exp_f := 0;
        ELSIF x =- 19894 THEN
            exp_f := 0;
        ELSIF x =- 19893 THEN
            exp_f := 0;
        ELSIF x =- 19892 THEN
            exp_f := 0;
        ELSIF x =- 19891 THEN
            exp_f := 0;
        ELSIF x =- 19890 THEN
            exp_f := 0;
        ELSIF x =- 19889 THEN
            exp_f := 0;
        ELSIF x =- 19888 THEN
            exp_f := 0;
        ELSIF x =- 19887 THEN
            exp_f := 0;
        ELSIF x =- 19886 THEN
            exp_f := 0;
        ELSIF x =- 19885 THEN
            exp_f := 0;
        ELSIF x =- 19884 THEN
            exp_f := 0;
        ELSIF x =- 19883 THEN
            exp_f := 0;
        ELSIF x =- 19882 THEN
            exp_f := 0;
        ELSIF x =- 19881 THEN
            exp_f := 0;
        ELSIF x =- 19880 THEN
            exp_f := 0;
        ELSIF x =- 19879 THEN
            exp_f := 0;
        ELSIF x =- 19878 THEN
            exp_f := 0;
        ELSIF x =- 19877 THEN
            exp_f := 0;
        ELSIF x =- 19876 THEN
            exp_f := 0;
        ELSIF x =- 19875 THEN
            exp_f := 0;
        ELSIF x =- 19874 THEN
            exp_f := 0;
        ELSIF x =- 19873 THEN
            exp_f := 0;
        ELSIF x =- 19872 THEN
            exp_f := 0;
        ELSIF x =- 19871 THEN
            exp_f := 0;
        ELSIF x =- 19870 THEN
            exp_f := 0;
        ELSIF x =- 19869 THEN
            exp_f := 0;
        ELSIF x =- 19868 THEN
            exp_f := 0;
        ELSIF x =- 19867 THEN
            exp_f := 0;
        ELSIF x =- 19866 THEN
            exp_f := 0;
        ELSIF x =- 19865 THEN
            exp_f := 0;
        ELSIF x =- 19864 THEN
            exp_f := 0;
        ELSIF x =- 19863 THEN
            exp_f := 0;
        ELSIF x =- 19862 THEN
            exp_f := 0;
        ELSIF x =- 19861 THEN
            exp_f := 0;
        ELSIF x =- 19860 THEN
            exp_f := 0;
        ELSIF x =- 19859 THEN
            exp_f := 0;
        ELSIF x =- 19858 THEN
            exp_f := 0;
        ELSIF x =- 19857 THEN
            exp_f := 0;
        ELSIF x =- 19856 THEN
            exp_f := 0;
        ELSIF x =- 19855 THEN
            exp_f := 0;
        ELSIF x =- 19854 THEN
            exp_f := 0;
        ELSIF x =- 19853 THEN
            exp_f := 0;
        ELSIF x =- 19852 THEN
            exp_f := 0;
        ELSIF x =- 19851 THEN
            exp_f := 0;
        ELSIF x =- 19850 THEN
            exp_f := 0;
        ELSIF x =- 19849 THEN
            exp_f := 0;
        ELSIF x =- 19848 THEN
            exp_f := 0;
        ELSIF x =- 19847 THEN
            exp_f := 0;
        ELSIF x =- 19846 THEN
            exp_f := 0;
        ELSIF x =- 19845 THEN
            exp_f := 0;
        ELSIF x =- 19844 THEN
            exp_f := 0;
        ELSIF x =- 19843 THEN
            exp_f := 0;
        ELSIF x =- 19842 THEN
            exp_f := 0;
        ELSIF x =- 19841 THEN
            exp_f := 0;
        ELSIF x =- 19840 THEN
            exp_f := 0;
        ELSIF x =- 19839 THEN
            exp_f := 0;
        ELSIF x =- 19838 THEN
            exp_f := 0;
        ELSIF x =- 19837 THEN
            exp_f := 0;
        ELSIF x =- 19836 THEN
            exp_f := 0;
        ELSIF x =- 19835 THEN
            exp_f := 0;
        ELSIF x =- 19834 THEN
            exp_f := 0;
        ELSIF x =- 19833 THEN
            exp_f := 0;
        ELSIF x =- 19832 THEN
            exp_f := 0;
        ELSIF x =- 19831 THEN
            exp_f := 0;
        ELSIF x =- 19830 THEN
            exp_f := 0;
        ELSIF x =- 19829 THEN
            exp_f := 0;
        ELSIF x =- 19828 THEN
            exp_f := 0;
        ELSIF x =- 19827 THEN
            exp_f := 0;
        ELSIF x =- 19826 THEN
            exp_f := 0;
        ELSIF x =- 19825 THEN
            exp_f := 0;
        ELSIF x =- 19824 THEN
            exp_f := 0;
        ELSIF x =- 19823 THEN
            exp_f := 0;
        ELSIF x =- 19822 THEN
            exp_f := 0;
        ELSIF x =- 19821 THEN
            exp_f := 0;
        ELSIF x =- 19820 THEN
            exp_f := 0;
        ELSIF x =- 19819 THEN
            exp_f := 0;
        ELSIF x =- 19818 THEN
            exp_f := 0;
        ELSIF x =- 19817 THEN
            exp_f := 0;
        ELSIF x =- 19816 THEN
            exp_f := 0;
        ELSIF x =- 19815 THEN
            exp_f := 0;
        ELSIF x =- 19814 THEN
            exp_f := 0;
        ELSIF x =- 19813 THEN
            exp_f := 0;
        ELSIF x =- 19812 THEN
            exp_f := 0;
        ELSIF x =- 19811 THEN
            exp_f := 0;
        ELSIF x =- 19810 THEN
            exp_f := 0;
        ELSIF x =- 19809 THEN
            exp_f := 0;
        ELSIF x =- 19808 THEN
            exp_f := 0;
        ELSIF x =- 19807 THEN
            exp_f := 0;
        ELSIF x =- 19806 THEN
            exp_f := 0;
        ELSIF x =- 19805 THEN
            exp_f := 0;
        ELSIF x =- 19804 THEN
            exp_f := 0;
        ELSIF x =- 19803 THEN
            exp_f := 0;
        ELSIF x =- 19802 THEN
            exp_f := 0;
        ELSIF x =- 19801 THEN
            exp_f := 0;
        ELSIF x =- 19800 THEN
            exp_f := 0;
        ELSIF x =- 19799 THEN
            exp_f := 0;
        ELSIF x =- 19798 THEN
            exp_f := 0;
        ELSIF x =- 19797 THEN
            exp_f := 0;
        ELSIF x =- 19796 THEN
            exp_f := 0;
        ELSIF x =- 19795 THEN
            exp_f := 0;
        ELSIF x =- 19794 THEN
            exp_f := 0;
        ELSIF x =- 19793 THEN
            exp_f := 0;
        ELSIF x =- 19792 THEN
            exp_f := 0;
        ELSIF x =- 19791 THEN
            exp_f := 0;
        ELSIF x =- 19790 THEN
            exp_f := 0;
        ELSIF x =- 19789 THEN
            exp_f := 0;
        ELSIF x =- 19788 THEN
            exp_f := 0;
        ELSIF x =- 19787 THEN
            exp_f := 0;
        ELSIF x =- 19786 THEN
            exp_f := 0;
        ELSIF x =- 19785 THEN
            exp_f := 0;
        ELSIF x =- 19784 THEN
            exp_f := 0;
        ELSIF x =- 19783 THEN
            exp_f := 0;
        ELSIF x =- 19782 THEN
            exp_f := 0;
        ELSIF x =- 19781 THEN
            exp_f := 0;
        ELSIF x =- 19780 THEN
            exp_f := 0;
        ELSIF x =- 19779 THEN
            exp_f := 0;
        ELSIF x =- 19778 THEN
            exp_f := 0;
        ELSIF x =- 19777 THEN
            exp_f := 0;
        ELSIF x =- 19776 THEN
            exp_f := 0;
        ELSIF x =- 19775 THEN
            exp_f := 0;
        ELSIF x =- 19774 THEN
            exp_f := 0;
        ELSIF x =- 19773 THEN
            exp_f := 0;
        ELSIF x =- 19772 THEN
            exp_f := 0;
        ELSIF x =- 19771 THEN
            exp_f := 0;
        ELSIF x =- 19770 THEN
            exp_f := 0;
        ELSIF x =- 19769 THEN
            exp_f := 0;
        ELSIF x =- 19768 THEN
            exp_f := 0;
        ELSIF x =- 19767 THEN
            exp_f := 0;
        ELSIF x =- 19766 THEN
            exp_f := 0;
        ELSIF x =- 19765 THEN
            exp_f := 0;
        ELSIF x =- 19764 THEN
            exp_f := 0;
        ELSIF x =- 19763 THEN
            exp_f := 0;
        ELSIF x =- 19762 THEN
            exp_f := 0;
        ELSIF x =- 19761 THEN
            exp_f := 0;
        ELSIF x =- 19760 THEN
            exp_f := 0;
        ELSIF x =- 19759 THEN
            exp_f := 0;
        ELSIF x =- 19758 THEN
            exp_f := 0;
        ELSIF x =- 19757 THEN
            exp_f := 0;
        ELSIF x =- 19756 THEN
            exp_f := 0;
        ELSIF x =- 19755 THEN
            exp_f := 0;
        ELSIF x =- 19754 THEN
            exp_f := 0;
        ELSIF x =- 19753 THEN
            exp_f := 0;
        ELSIF x =- 19752 THEN
            exp_f := 0;
        ELSIF x =- 19751 THEN
            exp_f := 0;
        ELSIF x =- 19750 THEN
            exp_f := 0;
        ELSIF x =- 19749 THEN
            exp_f := 0;
        ELSIF x =- 19748 THEN
            exp_f := 0;
        ELSIF x =- 19747 THEN
            exp_f := 0;
        ELSIF x =- 19746 THEN
            exp_f := 0;
        ELSIF x =- 19745 THEN
            exp_f := 0;
        ELSIF x =- 19744 THEN
            exp_f := 0;
        ELSIF x =- 19743 THEN
            exp_f := 0;
        ELSIF x =- 19742 THEN
            exp_f := 0;
        ELSIF x =- 19741 THEN
            exp_f := 0;
        ELSIF x =- 19740 THEN
            exp_f := 0;
        ELSIF x =- 19739 THEN
            exp_f := 0;
        ELSIF x =- 19738 THEN
            exp_f := 0;
        ELSIF x =- 19737 THEN
            exp_f := 0;
        ELSIF x =- 19736 THEN
            exp_f := 0;
        ELSIF x =- 19735 THEN
            exp_f := 0;
        ELSIF x =- 19734 THEN
            exp_f := 0;
        ELSIF x =- 19733 THEN
            exp_f := 0;
        ELSIF x =- 19732 THEN
            exp_f := 0;
        ELSIF x =- 19731 THEN
            exp_f := 0;
        ELSIF x =- 19730 THEN
            exp_f := 0;
        ELSIF x =- 19729 THEN
            exp_f := 0;
        ELSIF x =- 19728 THEN
            exp_f := 0;
        ELSIF x =- 19727 THEN
            exp_f := 0;
        ELSIF x =- 19726 THEN
            exp_f := 0;
        ELSIF x =- 19725 THEN
            exp_f := 0;
        ELSIF x =- 19724 THEN
            exp_f := 0;
        ELSIF x =- 19723 THEN
            exp_f := 0;
        ELSIF x =- 19722 THEN
            exp_f := 0;
        ELSIF x =- 19721 THEN
            exp_f := 0;
        ELSIF x =- 19720 THEN
            exp_f := 0;
        ELSIF x =- 19719 THEN
            exp_f := 0;
        ELSIF x =- 19718 THEN
            exp_f := 0;
        ELSIF x =- 19717 THEN
            exp_f := 0;
        ELSIF x =- 19716 THEN
            exp_f := 0;
        ELSIF x =- 19715 THEN
            exp_f := 0;
        ELSIF x =- 19714 THEN
            exp_f := 0;
        ELSIF x =- 19713 THEN
            exp_f := 0;
        ELSIF x =- 19712 THEN
            exp_f := 0;
        ELSIF x =- 19711 THEN
            exp_f := 0;
        ELSIF x =- 19710 THEN
            exp_f := 0;
        ELSIF x =- 19709 THEN
            exp_f := 0;
        ELSIF x =- 19708 THEN
            exp_f := 0;
        ELSIF x =- 19707 THEN
            exp_f := 0;
        ELSIF x =- 19706 THEN
            exp_f := 0;
        ELSIF x =- 19705 THEN
            exp_f := 0;
        ELSIF x =- 19704 THEN
            exp_f := 0;
        ELSIF x =- 19703 THEN
            exp_f := 0;
        ELSIF x =- 19702 THEN
            exp_f := 0;
        ELSIF x =- 19701 THEN
            exp_f := 0;
        ELSIF x =- 19700 THEN
            exp_f := 0;
        ELSIF x =- 19699 THEN
            exp_f := 0;
        ELSIF x =- 19698 THEN
            exp_f := 0;
        ELSIF x =- 19697 THEN
            exp_f := 0;
        ELSIF x =- 19696 THEN
            exp_f := 0;
        ELSIF x =- 19695 THEN
            exp_f := 0;
        ELSIF x =- 19694 THEN
            exp_f := 0;
        ELSIF x =- 19693 THEN
            exp_f := 0;
        ELSIF x =- 19692 THEN
            exp_f := 0;
        ELSIF x =- 19691 THEN
            exp_f := 0;
        ELSIF x =- 19690 THEN
            exp_f := 0;
        ELSIF x =- 19689 THEN
            exp_f := 0;
        ELSIF x =- 19688 THEN
            exp_f := 0;
        ELSIF x =- 19687 THEN
            exp_f := 0;
        ELSIF x =- 19686 THEN
            exp_f := 0;
        ELSIF x =- 19685 THEN
            exp_f := 0;
        ELSIF x =- 19684 THEN
            exp_f := 0;
        ELSIF x =- 19683 THEN
            exp_f := 0;
        ELSIF x =- 19682 THEN
            exp_f := 0;
        ELSIF x =- 19681 THEN
            exp_f := 0;
        ELSIF x =- 19680 THEN
            exp_f := 0;
        ELSIF x =- 19679 THEN
            exp_f := 0;
        ELSIF x =- 19678 THEN
            exp_f := 0;
        ELSIF x =- 19677 THEN
            exp_f := 0;
        ELSIF x =- 19676 THEN
            exp_f := 0;
        ELSIF x =- 19675 THEN
            exp_f := 0;
        ELSIF x =- 19674 THEN
            exp_f := 0;
        ELSIF x =- 19673 THEN
            exp_f := 0;
        ELSIF x =- 19672 THEN
            exp_f := 0;
        ELSIF x =- 19671 THEN
            exp_f := 0;
        ELSIF x =- 19670 THEN
            exp_f := 0;
        ELSIF x =- 19669 THEN
            exp_f := 0;
        ELSIF x =- 19668 THEN
            exp_f := 0;
        ELSIF x =- 19667 THEN
            exp_f := 0;
        ELSIF x =- 19666 THEN
            exp_f := 0;
        ELSIF x =- 19665 THEN
            exp_f := 0;
        ELSIF x =- 19664 THEN
            exp_f := 0;
        ELSIF x =- 19663 THEN
            exp_f := 0;
        ELSIF x =- 19662 THEN
            exp_f := 0;
        ELSIF x =- 19661 THEN
            exp_f := 0;
        ELSIF x =- 19660 THEN
            exp_f := 0;
        ELSIF x =- 19659 THEN
            exp_f := 0;
        ELSIF x =- 19658 THEN
            exp_f := 0;
        ELSIF x =- 19657 THEN
            exp_f := 0;
        ELSIF x =- 19656 THEN
            exp_f := 0;
        ELSIF x =- 19655 THEN
            exp_f := 0;
        ELSIF x =- 19654 THEN
            exp_f := 0;
        ELSIF x =- 19653 THEN
            exp_f := 0;
        ELSIF x =- 19652 THEN
            exp_f := 0;
        ELSIF x =- 19651 THEN
            exp_f := 0;
        ELSIF x =- 19650 THEN
            exp_f := 0;
        ELSIF x =- 19649 THEN
            exp_f := 0;
        ELSIF x =- 19648 THEN
            exp_f := 0;
        ELSIF x =- 19647 THEN
            exp_f := 0;
        ELSIF x =- 19646 THEN
            exp_f := 0;
        ELSIF x =- 19645 THEN
            exp_f := 0;
        ELSIF x =- 19644 THEN
            exp_f := 0;
        ELSIF x =- 19643 THEN
            exp_f := 0;
        ELSIF x =- 19642 THEN
            exp_f := 0;
        ELSIF x =- 19641 THEN
            exp_f := 0;
        ELSIF x =- 19640 THEN
            exp_f := 0;
        ELSIF x =- 19639 THEN
            exp_f := 0;
        ELSIF x =- 19638 THEN
            exp_f := 0;
        ELSIF x =- 19637 THEN
            exp_f := 0;
        ELSIF x =- 19636 THEN
            exp_f := 0;
        ELSIF x =- 19635 THEN
            exp_f := 0;
        ELSIF x =- 19634 THEN
            exp_f := 0;
        ELSIF x =- 19633 THEN
            exp_f := 0;
        ELSIF x =- 19632 THEN
            exp_f := 0;
        ELSIF x =- 19631 THEN
            exp_f := 0;
        ELSIF x =- 19630 THEN
            exp_f := 0;
        ELSIF x =- 19629 THEN
            exp_f := 0;
        ELSIF x =- 19628 THEN
            exp_f := 0;
        ELSIF x =- 19627 THEN
            exp_f := 0;
        ELSIF x =- 19626 THEN
            exp_f := 0;
        ELSIF x =- 19625 THEN
            exp_f := 0;
        ELSIF x =- 19624 THEN
            exp_f := 0;
        ELSIF x =- 19623 THEN
            exp_f := 0;
        ELSIF x =- 19622 THEN
            exp_f := 0;
        ELSIF x =- 19621 THEN
            exp_f := 0;
        ELSIF x =- 19620 THEN
            exp_f := 0;
        ELSIF x =- 19619 THEN
            exp_f := 0;
        ELSIF x =- 19618 THEN
            exp_f := 0;
        ELSIF x =- 19617 THEN
            exp_f := 0;
        ELSIF x =- 19616 THEN
            exp_f := 0;
        ELSIF x =- 19615 THEN
            exp_f := 0;
        ELSIF x =- 19614 THEN
            exp_f := 0;
        ELSIF x =- 19613 THEN
            exp_f := 0;
        ELSIF x =- 19612 THEN
            exp_f := 0;
        ELSIF x =- 19611 THEN
            exp_f := 0;
        ELSIF x =- 19610 THEN
            exp_f := 0;
        ELSIF x =- 19609 THEN
            exp_f := 0;
        ELSIF x =- 19608 THEN
            exp_f := 0;
        ELSIF x =- 19607 THEN
            exp_f := 0;
        ELSIF x =- 19606 THEN
            exp_f := 0;
        ELSIF x =- 19605 THEN
            exp_f := 0;
        ELSIF x =- 19604 THEN
            exp_f := 0;
        ELSIF x =- 19603 THEN
            exp_f := 0;
        ELSIF x =- 19602 THEN
            exp_f := 0;
        ELSIF x =- 19601 THEN
            exp_f := 0;
        ELSIF x =- 19600 THEN
            exp_f := 0;
        ELSIF x =- 19599 THEN
            exp_f := 0;
        ELSIF x =- 19598 THEN
            exp_f := 0;
        ELSIF x =- 19597 THEN
            exp_f := 0;
        ELSIF x =- 19596 THEN
            exp_f := 0;
        ELSIF x =- 19595 THEN
            exp_f := 0;
        ELSIF x =- 19594 THEN
            exp_f := 0;
        ELSIF x =- 19593 THEN
            exp_f := 0;
        ELSIF x =- 19592 THEN
            exp_f := 0;
        ELSIF x =- 19591 THEN
            exp_f := 0;
        ELSIF x =- 19590 THEN
            exp_f := 0;
        ELSIF x =- 19589 THEN
            exp_f := 0;
        ELSIF x =- 19588 THEN
            exp_f := 0;
        ELSIF x =- 19587 THEN
            exp_f := 0;
        ELSIF x =- 19586 THEN
            exp_f := 0;
        ELSIF x =- 19585 THEN
            exp_f := 0;
        ELSIF x =- 19584 THEN
            exp_f := 0;
        ELSIF x =- 19583 THEN
            exp_f := 0;
        ELSIF x =- 19582 THEN
            exp_f := 0;
        ELSIF x =- 19581 THEN
            exp_f := 0;
        ELSIF x =- 19580 THEN
            exp_f := 0;
        ELSIF x =- 19579 THEN
            exp_f := 0;
        ELSIF x =- 19578 THEN
            exp_f := 0;
        ELSIF x =- 19577 THEN
            exp_f := 0;
        ELSIF x =- 19576 THEN
            exp_f := 0;
        ELSIF x =- 19575 THEN
            exp_f := 0;
        ELSIF x =- 19574 THEN
            exp_f := 0;
        ELSIF x =- 19573 THEN
            exp_f := 0;
        ELSIF x =- 19572 THEN
            exp_f := 0;
        ELSIF x =- 19571 THEN
            exp_f := 0;
        ELSIF x =- 19570 THEN
            exp_f := 0;
        ELSIF x =- 19569 THEN
            exp_f := 0;
        ELSIF x =- 19568 THEN
            exp_f := 0;
        ELSIF x =- 19567 THEN
            exp_f := 0;
        ELSIF x =- 19566 THEN
            exp_f := 0;
        ELSIF x =- 19565 THEN
            exp_f := 0;
        ELSIF x =- 19564 THEN
            exp_f := 0;
        ELSIF x =- 19563 THEN
            exp_f := 0;
        ELSIF x =- 19562 THEN
            exp_f := 0;
        ELSIF x =- 19561 THEN
            exp_f := 0;
        ELSIF x =- 19560 THEN
            exp_f := 0;
        ELSIF x =- 19559 THEN
            exp_f := 0;
        ELSIF x =- 19558 THEN
            exp_f := 0;
        ELSIF x =- 19557 THEN
            exp_f := 0;
        ELSIF x =- 19556 THEN
            exp_f := 0;
        ELSIF x =- 19555 THEN
            exp_f := 0;
        ELSIF x =- 19554 THEN
            exp_f := 0;
        ELSIF x =- 19553 THEN
            exp_f := 0;
        ELSIF x =- 19552 THEN
            exp_f := 0;
        ELSIF x =- 19551 THEN
            exp_f := 0;
        ELSIF x =- 19550 THEN
            exp_f := 0;
        ELSIF x =- 19549 THEN
            exp_f := 0;
        ELSIF x =- 19548 THEN
            exp_f := 0;
        ELSIF x =- 19547 THEN
            exp_f := 0;
        ELSIF x =- 19546 THEN
            exp_f := 0;
        ELSIF x =- 19545 THEN
            exp_f := 0;
        ELSIF x =- 19544 THEN
            exp_f := 0;
        ELSIF x =- 19543 THEN
            exp_f := 0;
        ELSIF x =- 19542 THEN
            exp_f := 0;
        ELSIF x =- 19541 THEN
            exp_f := 0;
        ELSIF x =- 19540 THEN
            exp_f := 0;
        ELSIF x =- 19539 THEN
            exp_f := 0;
        ELSIF x =- 19538 THEN
            exp_f := 0;
        ELSIF x =- 19537 THEN
            exp_f := 0;
        ELSIF x =- 19536 THEN
            exp_f := 0;
        ELSIF x =- 19535 THEN
            exp_f := 0;
        ELSIF x =- 19534 THEN
            exp_f := 0;
        ELSIF x =- 19533 THEN
            exp_f := 0;
        ELSIF x =- 19532 THEN
            exp_f := 0;
        ELSIF x =- 19531 THEN
            exp_f := 0;
        ELSIF x =- 19530 THEN
            exp_f := 0;
        ELSIF x =- 19529 THEN
            exp_f := 0;
        ELSIF x =- 19528 THEN
            exp_f := 0;
        ELSIF x =- 19527 THEN
            exp_f := 0;
        ELSIF x =- 19526 THEN
            exp_f := 0;
        ELSIF x =- 19525 THEN
            exp_f := 0;
        ELSIF x =- 19524 THEN
            exp_f := 0;
        ELSIF x =- 19523 THEN
            exp_f := 0;
        ELSIF x =- 19522 THEN
            exp_f := 0;
        ELSIF x =- 19521 THEN
            exp_f := 0;
        ELSIF x =- 19520 THEN
            exp_f := 0;
        ELSIF x =- 19519 THEN
            exp_f := 0;
        ELSIF x =- 19518 THEN
            exp_f := 0;
        ELSIF x =- 19517 THEN
            exp_f := 0;
        ELSIF x =- 19516 THEN
            exp_f := 0;
        ELSIF x =- 19515 THEN
            exp_f := 0;
        ELSIF x =- 19514 THEN
            exp_f := 0;
        ELSIF x =- 19513 THEN
            exp_f := 0;
        ELSIF x =- 19512 THEN
            exp_f := 0;
        ELSIF x =- 19511 THEN
            exp_f := 0;
        ELSIF x =- 19510 THEN
            exp_f := 0;
        ELSIF x =- 19509 THEN
            exp_f := 0;
        ELSIF x =- 19508 THEN
            exp_f := 0;
        ELSIF x =- 19507 THEN
            exp_f := 0;
        ELSIF x =- 19506 THEN
            exp_f := 0;
        ELSIF x =- 19505 THEN
            exp_f := 0;
        ELSIF x =- 19504 THEN
            exp_f := 0;
        ELSIF x =- 19503 THEN
            exp_f := 0;
        ELSIF x =- 19502 THEN
            exp_f := 0;
        ELSIF x =- 19501 THEN
            exp_f := 0;
        ELSIF x =- 19500 THEN
            exp_f := 0;
        ELSIF x =- 19499 THEN
            exp_f := 0;
        ELSIF x =- 19498 THEN
            exp_f := 0;
        ELSIF x =- 19497 THEN
            exp_f := 0;
        ELSIF x =- 19496 THEN
            exp_f := 0;
        ELSIF x =- 19495 THEN
            exp_f := 0;
        ELSIF x =- 19494 THEN
            exp_f := 0;
        ELSIF x =- 19493 THEN
            exp_f := 0;
        ELSIF x =- 19492 THEN
            exp_f := 0;
        ELSIF x =- 19491 THEN
            exp_f := 0;
        ELSIF x =- 19490 THEN
            exp_f := 0;
        ELSIF x =- 19489 THEN
            exp_f := 0;
        ELSIF x =- 19488 THEN
            exp_f := 0;
        ELSIF x =- 19487 THEN
            exp_f := 0;
        ELSIF x =- 19486 THEN
            exp_f := 0;
        ELSIF x =- 19485 THEN
            exp_f := 0;
        ELSIF x =- 19484 THEN
            exp_f := 0;
        ELSIF x =- 19483 THEN
            exp_f := 0;
        ELSIF x =- 19482 THEN
            exp_f := 0;
        ELSIF x =- 19481 THEN
            exp_f := 0;
        ELSIF x =- 19480 THEN
            exp_f := 0;
        ELSIF x =- 19479 THEN
            exp_f := 0;
        ELSIF x =- 19478 THEN
            exp_f := 0;
        ELSIF x =- 19477 THEN
            exp_f := 0;
        ELSIF x =- 19476 THEN
            exp_f := 0;
        ELSIF x =- 19475 THEN
            exp_f := 0;
        ELSIF x =- 19474 THEN
            exp_f := 0;
        ELSIF x =- 19473 THEN
            exp_f := 0;
        ELSIF x =- 19472 THEN
            exp_f := 0;
        ELSIF x =- 19471 THEN
            exp_f := 0;
        ELSIF x =- 19470 THEN
            exp_f := 0;
        ELSIF x =- 19469 THEN
            exp_f := 0;
        ELSIF x =- 19468 THEN
            exp_f := 0;
        ELSIF x =- 19467 THEN
            exp_f := 0;
        ELSIF x =- 19466 THEN
            exp_f := 0;
        ELSIF x =- 19465 THEN
            exp_f := 0;
        ELSIF x =- 19464 THEN
            exp_f := 0;
        ELSIF x =- 19463 THEN
            exp_f := 0;
        ELSIF x =- 19462 THEN
            exp_f := 0;
        ELSIF x =- 19461 THEN
            exp_f := 0;
        ELSIF x =- 19460 THEN
            exp_f := 0;
        ELSIF x =- 19459 THEN
            exp_f := 0;
        ELSIF x =- 19458 THEN
            exp_f := 0;
        ELSIF x =- 19457 THEN
            exp_f := 0;
        ELSIF x =- 19456 THEN
            exp_f := 0;
        ELSIF x =- 19455 THEN
            exp_f := 0;
        ELSIF x =- 19454 THEN
            exp_f := 0;
        ELSIF x =- 19453 THEN
            exp_f := 0;
        ELSIF x =- 19452 THEN
            exp_f := 0;
        ELSIF x =- 19451 THEN
            exp_f := 0;
        ELSIF x =- 19450 THEN
            exp_f := 0;
        ELSIF x =- 19449 THEN
            exp_f := 0;
        ELSIF x =- 19448 THEN
            exp_f := 0;
        ELSIF x =- 19447 THEN
            exp_f := 0;
        ELSIF x =- 19446 THEN
            exp_f := 0;
        ELSIF x =- 19445 THEN
            exp_f := 0;
        ELSIF x =- 19444 THEN
            exp_f := 0;
        ELSIF x =- 19443 THEN
            exp_f := 0;
        ELSIF x =- 19442 THEN
            exp_f := 0;
        ELSIF x =- 19441 THEN
            exp_f := 0;
        ELSIF x =- 19440 THEN
            exp_f := 0;
        ELSIF x =- 19439 THEN
            exp_f := 0;
        ELSIF x =- 19438 THEN
            exp_f := 0;
        ELSIF x =- 19437 THEN
            exp_f := 0;
        ELSIF x =- 19436 THEN
            exp_f := 0;
        ELSIF x =- 19435 THEN
            exp_f := 0;
        ELSIF x =- 19434 THEN
            exp_f := 0;
        ELSIF x =- 19433 THEN
            exp_f := 0;
        ELSIF x =- 19432 THEN
            exp_f := 0;
        ELSIF x =- 19431 THEN
            exp_f := 0;
        ELSIF x =- 19430 THEN
            exp_f := 0;
        ELSIF x =- 19429 THEN
            exp_f := 0;
        ELSIF x =- 19428 THEN
            exp_f := 0;
        ELSIF x =- 19427 THEN
            exp_f := 0;
        ELSIF x =- 19426 THEN
            exp_f := 0;
        ELSIF x =- 19425 THEN
            exp_f := 0;
        ELSIF x =- 19424 THEN
            exp_f := 0;
        ELSIF x =- 19423 THEN
            exp_f := 0;
        ELSIF x =- 19422 THEN
            exp_f := 0;
        ELSIF x =- 19421 THEN
            exp_f := 0;
        ELSIF x =- 19420 THEN
            exp_f := 0;
        ELSIF x =- 19419 THEN
            exp_f := 0;
        ELSIF x =- 19418 THEN
            exp_f := 0;
        ELSIF x =- 19417 THEN
            exp_f := 0;
        ELSIF x =- 19416 THEN
            exp_f := 0;
        ELSIF x =- 19415 THEN
            exp_f := 0;
        ELSIF x =- 19414 THEN
            exp_f := 0;
        ELSIF x =- 19413 THEN
            exp_f := 0;
        ELSIF x =- 19412 THEN
            exp_f := 0;
        ELSIF x =- 19411 THEN
            exp_f := 0;
        ELSIF x =- 19410 THEN
            exp_f := 0;
        ELSIF x =- 19409 THEN
            exp_f := 0;
        ELSIF x =- 19408 THEN
            exp_f := 0;
        ELSIF x =- 19407 THEN
            exp_f := 0;
        ELSIF x =- 19406 THEN
            exp_f := 0;
        ELSIF x =- 19405 THEN
            exp_f := 0;
        ELSIF x =- 19404 THEN
            exp_f := 0;
        ELSIF x =- 19403 THEN
            exp_f := 0;
        ELSIF x =- 19402 THEN
            exp_f := 0;
        ELSIF x =- 19401 THEN
            exp_f := 0;
        ELSIF x =- 19400 THEN
            exp_f := 0;
        ELSIF x =- 19399 THEN
            exp_f := 0;
        ELSIF x =- 19398 THEN
            exp_f := 0;
        ELSIF x =- 19397 THEN
            exp_f := 0;
        ELSIF x =- 19396 THEN
            exp_f := 0;
        ELSIF x =- 19395 THEN
            exp_f := 0;
        ELSIF x =- 19394 THEN
            exp_f := 0;
        ELSIF x =- 19393 THEN
            exp_f := 0;
        ELSIF x =- 19392 THEN
            exp_f := 0;
        ELSIF x =- 19391 THEN
            exp_f := 0;
        ELSIF x =- 19390 THEN
            exp_f := 0;
        ELSIF x =- 19389 THEN
            exp_f := 0;
        ELSIF x =- 19388 THEN
            exp_f := 0;
        ELSIF x =- 19387 THEN
            exp_f := 0;
        ELSIF x =- 19386 THEN
            exp_f := 0;
        ELSIF x =- 19385 THEN
            exp_f := 0;
        ELSIF x =- 19384 THEN
            exp_f := 0;
        ELSIF x =- 19383 THEN
            exp_f := 0;
        ELSIF x =- 19382 THEN
            exp_f := 0;
        ELSIF x =- 19381 THEN
            exp_f := 0;
        ELSIF x =- 19380 THEN
            exp_f := 0;
        ELSIF x =- 19379 THEN
            exp_f := 0;
        ELSIF x =- 19378 THEN
            exp_f := 0;
        ELSIF x =- 19377 THEN
            exp_f := 0;
        ELSIF x =- 19376 THEN
            exp_f := 0;
        ELSIF x =- 19375 THEN
            exp_f := 0;
        ELSIF x =- 19374 THEN
            exp_f := 0;
        ELSIF x =- 19373 THEN
            exp_f := 0;
        ELSIF x =- 19372 THEN
            exp_f := 0;
        ELSIF x =- 19371 THEN
            exp_f := 0;
        ELSIF x =- 19370 THEN
            exp_f := 0;
        ELSIF x =- 19369 THEN
            exp_f := 0;
        ELSIF x =- 19368 THEN
            exp_f := 0;
        ELSIF x =- 19367 THEN
            exp_f := 0;
        ELSIF x =- 19366 THEN
            exp_f := 0;
        ELSIF x =- 19365 THEN
            exp_f := 0;
        ELSIF x =- 19364 THEN
            exp_f := 0;
        ELSIF x =- 19363 THEN
            exp_f := 0;
        ELSIF x =- 19362 THEN
            exp_f := 0;
        ELSIF x =- 19361 THEN
            exp_f := 0;
        ELSIF x =- 19360 THEN
            exp_f := 0;
        ELSIF x =- 19359 THEN
            exp_f := 0;
        ELSIF x =- 19358 THEN
            exp_f := 0;
        ELSIF x =- 19357 THEN
            exp_f := 0;
        ELSIF x =- 19356 THEN
            exp_f := 0;
        ELSIF x =- 19355 THEN
            exp_f := 0;
        ELSIF x =- 19354 THEN
            exp_f := 0;
        ELSIF x =- 19353 THEN
            exp_f := 0;
        ELSIF x =- 19352 THEN
            exp_f := 0;
        ELSIF x =- 19351 THEN
            exp_f := 0;
        ELSIF x =- 19350 THEN
            exp_f := 0;
        ELSIF x =- 19349 THEN
            exp_f := 0;
        ELSIF x =- 19348 THEN
            exp_f := 0;
        ELSIF x =- 19347 THEN
            exp_f := 0;
        ELSIF x =- 19346 THEN
            exp_f := 0;
        ELSIF x =- 19345 THEN
            exp_f := 0;
        ELSIF x =- 19344 THEN
            exp_f := 0;
        ELSIF x =- 19343 THEN
            exp_f := 0;
        ELSIF x =- 19342 THEN
            exp_f := 0;
        ELSIF x =- 19341 THEN
            exp_f := 0;
        ELSIF x =- 19340 THEN
            exp_f := 0;
        ELSIF x =- 19339 THEN
            exp_f := 0;
        ELSIF x =- 19338 THEN
            exp_f := 0;
        ELSIF x =- 19337 THEN
            exp_f := 0;
        ELSIF x =- 19336 THEN
            exp_f := 0;
        ELSIF x =- 19335 THEN
            exp_f := 0;
        ELSIF x =- 19334 THEN
            exp_f := 0;
        ELSIF x =- 19333 THEN
            exp_f := 0;
        ELSIF x =- 19332 THEN
            exp_f := 0;
        ELSIF x =- 19331 THEN
            exp_f := 0;
        ELSIF x =- 19330 THEN
            exp_f := 0;
        ELSIF x =- 19329 THEN
            exp_f := 0;
        ELSIF x =- 19328 THEN
            exp_f := 0;
        ELSIF x =- 19327 THEN
            exp_f := 0;
        ELSIF x =- 19326 THEN
            exp_f := 0;
        ELSIF x =- 19325 THEN
            exp_f := 0;
        ELSIF x =- 19324 THEN
            exp_f := 0;
        ELSIF x =- 19323 THEN
            exp_f := 0;
        ELSIF x =- 19322 THEN
            exp_f := 0;
        ELSIF x =- 19321 THEN
            exp_f := 0;
        ELSIF x =- 19320 THEN
            exp_f := 0;
        ELSIF x =- 19319 THEN
            exp_f := 0;
        ELSIF x =- 19318 THEN
            exp_f := 0;
        ELSIF x =- 19317 THEN
            exp_f := 0;
        ELSIF x =- 19316 THEN
            exp_f := 0;
        ELSIF x =- 19315 THEN
            exp_f := 0;
        ELSIF x =- 19314 THEN
            exp_f := 0;
        ELSIF x =- 19313 THEN
            exp_f := 0;
        ELSIF x =- 19312 THEN
            exp_f := 0;
        ELSIF x =- 19311 THEN
            exp_f := 0;
        ELSIF x =- 19310 THEN
            exp_f := 0;
        ELSIF x =- 19309 THEN
            exp_f := 0;
        ELSIF x =- 19308 THEN
            exp_f := 0;
        ELSIF x =- 19307 THEN
            exp_f := 0;
        ELSIF x =- 19306 THEN
            exp_f := 0;
        ELSIF x =- 19305 THEN
            exp_f := 0;
        ELSIF x =- 19304 THEN
            exp_f := 0;
        ELSIF x =- 19303 THEN
            exp_f := 0;
        ELSIF x =- 19302 THEN
            exp_f := 0;
        ELSIF x =- 19301 THEN
            exp_f := 0;
        ELSIF x =- 19300 THEN
            exp_f := 0;
        ELSIF x =- 19299 THEN
            exp_f := 0;
        ELSIF x =- 19298 THEN
            exp_f := 0;
        ELSIF x =- 19297 THEN
            exp_f := 0;
        ELSIF x =- 19296 THEN
            exp_f := 0;
        ELSIF x =- 19295 THEN
            exp_f := 0;
        ELSIF x =- 19294 THEN
            exp_f := 0;
        ELSIF x =- 19293 THEN
            exp_f := 0;
        ELSIF x =- 19292 THEN
            exp_f := 0;
        ELSIF x =- 19291 THEN
            exp_f := 0;
        ELSIF x =- 19290 THEN
            exp_f := 0;
        ELSIF x =- 19289 THEN
            exp_f := 0;
        ELSIF x =- 19288 THEN
            exp_f := 0;
        ELSIF x =- 19287 THEN
            exp_f := 0;
        ELSIF x =- 19286 THEN
            exp_f := 0;
        ELSIF x =- 19285 THEN
            exp_f := 0;
        ELSIF x =- 19284 THEN
            exp_f := 0;
        ELSIF x =- 19283 THEN
            exp_f := 0;
        ELSIF x =- 19282 THEN
            exp_f := 0;
        ELSIF x =- 19281 THEN
            exp_f := 0;
        ELSIF x =- 19280 THEN
            exp_f := 0;
        ELSIF x =- 19279 THEN
            exp_f := 0;
        ELSIF x =- 19278 THEN
            exp_f := 0;
        ELSIF x =- 19277 THEN
            exp_f := 0;
        ELSIF x =- 19276 THEN
            exp_f := 0;
        ELSIF x =- 19275 THEN
            exp_f := 0;
        ELSIF x =- 19274 THEN
            exp_f := 0;
        ELSIF x =- 19273 THEN
            exp_f := 0;
        ELSIF x =- 19272 THEN
            exp_f := 0;
        ELSIF x =- 19271 THEN
            exp_f := 0;
        ELSIF x =- 19270 THEN
            exp_f := 0;
        ELSIF x =- 19269 THEN
            exp_f := 0;
        ELSIF x =- 19268 THEN
            exp_f := 0;
        ELSIF x =- 19267 THEN
            exp_f := 0;
        ELSIF x =- 19266 THEN
            exp_f := 0;
        ELSIF x =- 19265 THEN
            exp_f := 0;
        ELSIF x =- 19264 THEN
            exp_f := 0;
        ELSIF x =- 19263 THEN
            exp_f := 0;
        ELSIF x =- 19262 THEN
            exp_f := 0;
        ELSIF x =- 19261 THEN
            exp_f := 0;
        ELSIF x =- 19260 THEN
            exp_f := 0;
        ELSIF x =- 19259 THEN
            exp_f := 0;
        ELSIF x =- 19258 THEN
            exp_f := 0;
        ELSIF x =- 19257 THEN
            exp_f := 0;
        ELSIF x =- 19256 THEN
            exp_f := 0;
        ELSIF x =- 19255 THEN
            exp_f := 0;
        ELSIF x =- 19254 THEN
            exp_f := 0;
        ELSIF x =- 19253 THEN
            exp_f := 0;
        ELSIF x =- 19252 THEN
            exp_f := 0;
        ELSIF x =- 19251 THEN
            exp_f := 0;
        ELSIF x =- 19250 THEN
            exp_f := 0;
        ELSIF x =- 19249 THEN
            exp_f := 0;
        ELSIF x =- 19248 THEN
            exp_f := 0;
        ELSIF x =- 19247 THEN
            exp_f := 0;
        ELSIF x =- 19246 THEN
            exp_f := 0;
        ELSIF x =- 19245 THEN
            exp_f := 0;
        ELSIF x =- 19244 THEN
            exp_f := 0;
        ELSIF x =- 19243 THEN
            exp_f := 0;
        ELSIF x =- 19242 THEN
            exp_f := 0;
        ELSIF x =- 19241 THEN
            exp_f := 0;
        ELSIF x =- 19240 THEN
            exp_f := 0;
        ELSIF x =- 19239 THEN
            exp_f := 0;
        ELSIF x =- 19238 THEN
            exp_f := 0;
        ELSIF x =- 19237 THEN
            exp_f := 0;
        ELSIF x =- 19236 THEN
            exp_f := 0;
        ELSIF x =- 19235 THEN
            exp_f := 0;
        ELSIF x =- 19234 THEN
            exp_f := 0;
        ELSIF x =- 19233 THEN
            exp_f := 0;
        ELSIF x =- 19232 THEN
            exp_f := 0;
        ELSIF x =- 19231 THEN
            exp_f := 0;
        ELSIF x =- 19230 THEN
            exp_f := 0;
        ELSIF x =- 19229 THEN
            exp_f := 0;
        ELSIF x =- 19228 THEN
            exp_f := 0;
        ELSIF x =- 19227 THEN
            exp_f := 0;
        ELSIF x =- 19226 THEN
            exp_f := 0;
        ELSIF x =- 19225 THEN
            exp_f := 0;
        ELSIF x =- 19224 THEN
            exp_f := 0;
        ELSIF x =- 19223 THEN
            exp_f := 0;
        ELSIF x =- 19222 THEN
            exp_f := 0;
        ELSIF x =- 19221 THEN
            exp_f := 0;
        ELSIF x =- 19220 THEN
            exp_f := 0;
        ELSIF x =- 19219 THEN
            exp_f := 0;
        ELSIF x =- 19218 THEN
            exp_f := 0;
        ELSIF x =- 19217 THEN
            exp_f := 0;
        ELSIF x =- 19216 THEN
            exp_f := 0;
        ELSIF x =- 19215 THEN
            exp_f := 0;
        ELSIF x =- 19214 THEN
            exp_f := 0;
        ELSIF x =- 19213 THEN
            exp_f := 0;
        ELSIF x =- 19212 THEN
            exp_f := 0;
        ELSIF x =- 19211 THEN
            exp_f := 0;
        ELSIF x =- 19210 THEN
            exp_f := 0;
        ELSIF x =- 19209 THEN
            exp_f := 0;
        ELSIF x =- 19208 THEN
            exp_f := 0;
        ELSIF x =- 19207 THEN
            exp_f := 0;
        ELSIF x =- 19206 THEN
            exp_f := 0;
        ELSIF x =- 19205 THEN
            exp_f := 0;
        ELSIF x =- 19204 THEN
            exp_f := 0;
        ELSIF x =- 19203 THEN
            exp_f := 0;
        ELSIF x =- 19202 THEN
            exp_f := 0;
        ELSIF x =- 19201 THEN
            exp_f := 0;
        ELSIF x =- 19200 THEN
            exp_f := 0;
        ELSIF x =- 19199 THEN
            exp_f := 0;
        ELSIF x =- 19198 THEN
            exp_f := 0;
        ELSIF x =- 19197 THEN
            exp_f := 0;
        ELSIF x =- 19196 THEN
            exp_f := 0;
        ELSIF x =- 19195 THEN
            exp_f := 0;
        ELSIF x =- 19194 THEN
            exp_f := 0;
        ELSIF x =- 19193 THEN
            exp_f := 0;
        ELSIF x =- 19192 THEN
            exp_f := 0;
        ELSIF x =- 19191 THEN
            exp_f := 0;
        ELSIF x =- 19190 THEN
            exp_f := 0;
        ELSIF x =- 19189 THEN
            exp_f := 0;
        ELSIF x =- 19188 THEN
            exp_f := 0;
        ELSIF x =- 19187 THEN
            exp_f := 0;
        ELSIF x =- 19186 THEN
            exp_f := 0;
        ELSIF x =- 19185 THEN
            exp_f := 0;
        ELSIF x =- 19184 THEN
            exp_f := 0;
        ELSIF x =- 19183 THEN
            exp_f := 0;
        ELSIF x =- 19182 THEN
            exp_f := 0;
        ELSIF x =- 19181 THEN
            exp_f := 0;
        ELSIF x =- 19180 THEN
            exp_f := 0;
        ELSIF x =- 19179 THEN
            exp_f := 0;
        ELSIF x =- 19178 THEN
            exp_f := 0;
        ELSIF x =- 19177 THEN
            exp_f := 0;
        ELSIF x =- 19176 THEN
            exp_f := 0;
        ELSIF x =- 19175 THEN
            exp_f := 0;
        ELSIF x =- 19174 THEN
            exp_f := 0;
        ELSIF x =- 19173 THEN
            exp_f := 0;
        ELSIF x =- 19172 THEN
            exp_f := 0;
        ELSIF x =- 19171 THEN
            exp_f := 0;
        ELSIF x =- 19170 THEN
            exp_f := 0;
        ELSIF x =- 19169 THEN
            exp_f := 0;
        ELSIF x =- 19168 THEN
            exp_f := 0;
        ELSIF x =- 19167 THEN
            exp_f := 0;
        ELSIF x =- 19166 THEN
            exp_f := 0;
        ELSIF x =- 19165 THEN
            exp_f := 0;
        ELSIF x =- 19164 THEN
            exp_f := 0;
        ELSIF x =- 19163 THEN
            exp_f := 0;
        ELSIF x =- 19162 THEN
            exp_f := 0;
        ELSIF x =- 19161 THEN
            exp_f := 0;
        ELSIF x =- 19160 THEN
            exp_f := 0;
        ELSIF x =- 19159 THEN
            exp_f := 0;
        ELSIF x =- 19158 THEN
            exp_f := 0;
        ELSIF x =- 19157 THEN
            exp_f := 0;
        ELSIF x =- 19156 THEN
            exp_f := 0;
        ELSIF x =- 19155 THEN
            exp_f := 0;
        ELSIF x =- 19154 THEN
            exp_f := 0;
        ELSIF x =- 19153 THEN
            exp_f := 0;
        ELSIF x =- 19152 THEN
            exp_f := 0;
        ELSIF x =- 19151 THEN
            exp_f := 0;
        ELSIF x =- 19150 THEN
            exp_f := 0;
        ELSIF x =- 19149 THEN
            exp_f := 0;
        ELSIF x =- 19148 THEN
            exp_f := 0;
        ELSIF x =- 19147 THEN
            exp_f := 0;
        ELSIF x =- 19146 THEN
            exp_f := 0;
        ELSIF x =- 19145 THEN
            exp_f := 0;
        ELSIF x =- 19144 THEN
            exp_f := 0;
        ELSIF x =- 19143 THEN
            exp_f := 0;
        ELSIF x =- 19142 THEN
            exp_f := 0;
        ELSIF x =- 19141 THEN
            exp_f := 0;
        ELSIF x =- 19140 THEN
            exp_f := 0;
        ELSIF x =- 19139 THEN
            exp_f := 0;
        ELSIF x =- 19138 THEN
            exp_f := 0;
        ELSIF x =- 19137 THEN
            exp_f := 0;
        ELSIF x =- 19136 THEN
            exp_f := 0;
        ELSIF x =- 19135 THEN
            exp_f := 0;
        ELSIF x =- 19134 THEN
            exp_f := 0;
        ELSIF x =- 19133 THEN
            exp_f := 0;
        ELSIF x =- 19132 THEN
            exp_f := 0;
        ELSIF x =- 19131 THEN
            exp_f := 0;
        ELSIF x =- 19130 THEN
            exp_f := 0;
        ELSIF x =- 19129 THEN
            exp_f := 0;
        ELSIF x =- 19128 THEN
            exp_f := 0;
        ELSIF x =- 19127 THEN
            exp_f := 0;
        ELSIF x =- 19126 THEN
            exp_f := 0;
        ELSIF x =- 19125 THEN
            exp_f := 0;
        ELSIF x =- 19124 THEN
            exp_f := 0;
        ELSIF x =- 19123 THEN
            exp_f := 0;
        ELSIF x =- 19122 THEN
            exp_f := 0;
        ELSIF x =- 19121 THEN
            exp_f := 0;
        ELSIF x =- 19120 THEN
            exp_f := 0;
        ELSIF x =- 19119 THEN
            exp_f := 0;
        ELSIF x =- 19118 THEN
            exp_f := 0;
        ELSIF x =- 19117 THEN
            exp_f := 0;
        ELSIF x =- 19116 THEN
            exp_f := 0;
        ELSIF x =- 19115 THEN
            exp_f := 0;
        ELSIF x =- 19114 THEN
            exp_f := 0;
        ELSIF x =- 19113 THEN
            exp_f := 0;
        ELSIF x =- 19112 THEN
            exp_f := 0;
        ELSIF x =- 19111 THEN
            exp_f := 0;
        ELSIF x =- 19110 THEN
            exp_f := 0;
        ELSIF x =- 19109 THEN
            exp_f := 0;
        ELSIF x =- 19108 THEN
            exp_f := 0;
        ELSIF x =- 19107 THEN
            exp_f := 0;
        ELSIF x =- 19106 THEN
            exp_f := 0;
        ELSIF x =- 19105 THEN
            exp_f := 0;
        ELSIF x =- 19104 THEN
            exp_f := 0;
        ELSIF x =- 19103 THEN
            exp_f := 0;
        ELSIF x =- 19102 THEN
            exp_f := 0;
        ELSIF x =- 19101 THEN
            exp_f := 0;
        ELSIF x =- 19100 THEN
            exp_f := 0;
        ELSIF x =- 19099 THEN
            exp_f := 0;
        ELSIF x =- 19098 THEN
            exp_f := 0;
        ELSIF x =- 19097 THEN
            exp_f := 0;
        ELSIF x =- 19096 THEN
            exp_f := 0;
        ELSIF x =- 19095 THEN
            exp_f := 0;
        ELSIF x =- 19094 THEN
            exp_f := 0;
        ELSIF x =- 19093 THEN
            exp_f := 0;
        ELSIF x =- 19092 THEN
            exp_f := 0;
        ELSIF x =- 19091 THEN
            exp_f := 0;
        ELSIF x =- 19090 THEN
            exp_f := 0;
        ELSIF x =- 19089 THEN
            exp_f := 0;
        ELSIF x =- 19088 THEN
            exp_f := 0;
        ELSIF x =- 19087 THEN
            exp_f := 0;
        ELSIF x =- 19086 THEN
            exp_f := 0;
        ELSIF x =- 19085 THEN
            exp_f := 0;
        ELSIF x =- 19084 THEN
            exp_f := 0;
        ELSIF x =- 19083 THEN
            exp_f := 0;
        ELSIF x =- 19082 THEN
            exp_f := 0;
        ELSIF x =- 19081 THEN
            exp_f := 0;
        ELSIF x =- 19080 THEN
            exp_f := 0;
        ELSIF x =- 19079 THEN
            exp_f := 0;
        ELSIF x =- 19078 THEN
            exp_f := 0;
        ELSIF x =- 19077 THEN
            exp_f := 0;
        ELSIF x =- 19076 THEN
            exp_f := 0;
        ELSIF x =- 19075 THEN
            exp_f := 0;
        ELSIF x =- 19074 THEN
            exp_f := 0;
        ELSIF x =- 19073 THEN
            exp_f := 0;
        ELSIF x =- 19072 THEN
            exp_f := 0;
        ELSIF x =- 19071 THEN
            exp_f := 0;
        ELSIF x =- 19070 THEN
            exp_f := 0;
        ELSIF x =- 19069 THEN
            exp_f := 0;
        ELSIF x =- 19068 THEN
            exp_f := 0;
        ELSIF x =- 19067 THEN
            exp_f := 0;
        ELSIF x =- 19066 THEN
            exp_f := 0;
        ELSIF x =- 19065 THEN
            exp_f := 0;
        ELSIF x =- 19064 THEN
            exp_f := 0;
        ELSIF x =- 19063 THEN
            exp_f := 0;
        ELSIF x =- 19062 THEN
            exp_f := 0;
        ELSIF x =- 19061 THEN
            exp_f := 0;
        ELSIF x =- 19060 THEN
            exp_f := 0;
        ELSIF x =- 19059 THEN
            exp_f := 0;
        ELSIF x =- 19058 THEN
            exp_f := 0;
        ELSIF x =- 19057 THEN
            exp_f := 0;
        ELSIF x =- 19056 THEN
            exp_f := 0;
        ELSIF x =- 19055 THEN
            exp_f := 0;
        ELSIF x =- 19054 THEN
            exp_f := 0;
        ELSIF x =- 19053 THEN
            exp_f := 0;
        ELSIF x =- 19052 THEN
            exp_f := 0;
        ELSIF x =- 19051 THEN
            exp_f := 0;
        ELSIF x =- 19050 THEN
            exp_f := 0;
        ELSIF x =- 19049 THEN
            exp_f := 0;
        ELSIF x =- 19048 THEN
            exp_f := 0;
        ELSIF x =- 19047 THEN
            exp_f := 0;
        ELSIF x =- 19046 THEN
            exp_f := 0;
        ELSIF x =- 19045 THEN
            exp_f := 0;
        ELSIF x =- 19044 THEN
            exp_f := 0;
        ELSIF x =- 19043 THEN
            exp_f := 0;
        ELSIF x =- 19042 THEN
            exp_f := 0;
        ELSIF x =- 19041 THEN
            exp_f := 0;
        ELSIF x =- 19040 THEN
            exp_f := 0;
        ELSIF x =- 19039 THEN
            exp_f := 0;
        ELSIF x =- 19038 THEN
            exp_f := 0;
        ELSIF x =- 19037 THEN
            exp_f := 0;
        ELSIF x =- 19036 THEN
            exp_f := 0;
        ELSIF x =- 19035 THEN
            exp_f := 0;
        ELSIF x =- 19034 THEN
            exp_f := 0;
        ELSIF x =- 19033 THEN
            exp_f := 0;
        ELSIF x =- 19032 THEN
            exp_f := 0;
        ELSIF x =- 19031 THEN
            exp_f := 0;
        ELSIF x =- 19030 THEN
            exp_f := 0;
        ELSIF x =- 19029 THEN
            exp_f := 0;
        ELSIF x =- 19028 THEN
            exp_f := 0;
        ELSIF x =- 19027 THEN
            exp_f := 0;
        ELSIF x =- 19026 THEN
            exp_f := 0;
        ELSIF x =- 19025 THEN
            exp_f := 0;
        ELSIF x =- 19024 THEN
            exp_f := 0;
        ELSIF x =- 19023 THEN
            exp_f := 0;
        ELSIF x =- 19022 THEN
            exp_f := 0;
        ELSIF x =- 19021 THEN
            exp_f := 0;
        ELSIF x =- 19020 THEN
            exp_f := 0;
        ELSIF x =- 19019 THEN
            exp_f := 0;
        ELSIF x =- 19018 THEN
            exp_f := 0;
        ELSIF x =- 19017 THEN
            exp_f := 0;
        ELSIF x =- 19016 THEN
            exp_f := 0;
        ELSIF x =- 19015 THEN
            exp_f := 0;
        ELSIF x =- 19014 THEN
            exp_f := 0;
        ELSIF x =- 19013 THEN
            exp_f := 0;
        ELSIF x =- 19012 THEN
            exp_f := 0;
        ELSIF x =- 19011 THEN
            exp_f := 0;
        ELSIF x =- 19010 THEN
            exp_f := 0;
        ELSIF x =- 19009 THEN
            exp_f := 0;
        ELSIF x =- 19008 THEN
            exp_f := 0;
        ELSIF x =- 19007 THEN
            exp_f := 0;
        ELSIF x =- 19006 THEN
            exp_f := 0;
        ELSIF x =- 19005 THEN
            exp_f := 0;
        ELSIF x =- 19004 THEN
            exp_f := 0;
        ELSIF x =- 19003 THEN
            exp_f := 0;
        ELSIF x =- 19002 THEN
            exp_f := 0;
        ELSIF x =- 19001 THEN
            exp_f := 0;
        ELSIF x =- 19000 THEN
            exp_f := 0;
        ELSIF x =- 18999 THEN
            exp_f := 0;
        ELSIF x =- 18998 THEN
            exp_f := 0;
        ELSIF x =- 18997 THEN
            exp_f := 0;
        ELSIF x =- 18996 THEN
            exp_f := 0;
        ELSIF x =- 18995 THEN
            exp_f := 0;
        ELSIF x =- 18994 THEN
            exp_f := 0;
        ELSIF x =- 18993 THEN
            exp_f := 0;
        ELSIF x =- 18992 THEN
            exp_f := 0;
        ELSIF x =- 18991 THEN
            exp_f := 0;
        ELSIF x =- 18990 THEN
            exp_f := 0;
        ELSIF x =- 18989 THEN
            exp_f := 0;
        ELSIF x =- 18988 THEN
            exp_f := 0;
        ELSIF x =- 18987 THEN
            exp_f := 0;
        ELSIF x =- 18986 THEN
            exp_f := 0;
        ELSIF x =- 18985 THEN
            exp_f := 0;
        ELSIF x =- 18984 THEN
            exp_f := 0;
        ELSIF x =- 18983 THEN
            exp_f := 0;
        ELSIF x =- 18982 THEN
            exp_f := 0;
        ELSIF x =- 18981 THEN
            exp_f := 0;
        ELSIF x =- 18980 THEN
            exp_f := 0;
        ELSIF x =- 18979 THEN
            exp_f := 0;
        ELSIF x =- 18978 THEN
            exp_f := 0;
        ELSIF x =- 18977 THEN
            exp_f := 0;
        ELSIF x =- 18976 THEN
            exp_f := 0;
        ELSIF x =- 18975 THEN
            exp_f := 0;
        ELSIF x =- 18974 THEN
            exp_f := 0;
        ELSIF x =- 18973 THEN
            exp_f := 0;
        ELSIF x =- 18972 THEN
            exp_f := 0;
        ELSIF x =- 18971 THEN
            exp_f := 0;
        ELSIF x =- 18970 THEN
            exp_f := 0;
        ELSIF x =- 18969 THEN
            exp_f := 0;
        ELSIF x =- 18968 THEN
            exp_f := 0;
        ELSIF x =- 18967 THEN
            exp_f := 0;
        ELSIF x =- 18966 THEN
            exp_f := 0;
        ELSIF x =- 18965 THEN
            exp_f := 0;
        ELSIF x =- 18964 THEN
            exp_f := 0;
        ELSIF x =- 18963 THEN
            exp_f := 0;
        ELSIF x =- 18962 THEN
            exp_f := 0;
        ELSIF x =- 18961 THEN
            exp_f := 0;
        ELSIF x =- 18960 THEN
            exp_f := 0;
        ELSIF x =- 18959 THEN
            exp_f := 0;
        ELSIF x =- 18958 THEN
            exp_f := 0;
        ELSIF x =- 18957 THEN
            exp_f := 0;
        ELSIF x =- 18956 THEN
            exp_f := 0;
        ELSIF x =- 18955 THEN
            exp_f := 0;
        ELSIF x =- 18954 THEN
            exp_f := 0;
        ELSIF x =- 18953 THEN
            exp_f := 0;
        ELSIF x =- 18952 THEN
            exp_f := 0;
        ELSIF x =- 18951 THEN
            exp_f := 0;
        ELSIF x =- 18950 THEN
            exp_f := 0;
        ELSIF x =- 18949 THEN
            exp_f := 0;
        ELSIF x =- 18948 THEN
            exp_f := 0;
        ELSIF x =- 18947 THEN
            exp_f := 0;
        ELSIF x =- 18946 THEN
            exp_f := 0;
        ELSIF x =- 18945 THEN
            exp_f := 0;
        ELSIF x =- 18944 THEN
            exp_f := 0;
        ELSIF x =- 18943 THEN
            exp_f := 0;
        ELSIF x =- 18942 THEN
            exp_f := 0;
        ELSIF x =- 18941 THEN
            exp_f := 0;
        ELSIF x =- 18940 THEN
            exp_f := 0;
        ELSIF x =- 18939 THEN
            exp_f := 0;
        ELSIF x =- 18938 THEN
            exp_f := 0;
        ELSIF x =- 18937 THEN
            exp_f := 0;
        ELSIF x =- 18936 THEN
            exp_f := 0;
        ELSIF x =- 18935 THEN
            exp_f := 0;
        ELSIF x =- 18934 THEN
            exp_f := 0;
        ELSIF x =- 18933 THEN
            exp_f := 0;
        ELSIF x =- 18932 THEN
            exp_f := 0;
        ELSIF x =- 18931 THEN
            exp_f := 0;
        ELSIF x =- 18930 THEN
            exp_f := 0;
        ELSIF x =- 18929 THEN
            exp_f := 0;
        ELSIF x =- 18928 THEN
            exp_f := 0;
        ELSIF x =- 18927 THEN
            exp_f := 0;
        ELSIF x =- 18926 THEN
            exp_f := 0;
        ELSIF x =- 18925 THEN
            exp_f := 0;
        ELSIF x =- 18924 THEN
            exp_f := 0;
        ELSIF x =- 18923 THEN
            exp_f := 0;
        ELSIF x =- 18922 THEN
            exp_f := 0;
        ELSIF x =- 18921 THEN
            exp_f := 0;
        ELSIF x =- 18920 THEN
            exp_f := 0;
        ELSIF x =- 18919 THEN
            exp_f := 0;
        ELSIF x =- 18918 THEN
            exp_f := 0;
        ELSIF x =- 18917 THEN
            exp_f := 0;
        ELSIF x =- 18916 THEN
            exp_f := 0;
        ELSIF x =- 18915 THEN
            exp_f := 0;
        ELSIF x =- 18914 THEN
            exp_f := 0;
        ELSIF x =- 18913 THEN
            exp_f := 0;
        ELSIF x =- 18912 THEN
            exp_f := 0;
        ELSIF x =- 18911 THEN
            exp_f := 0;
        ELSIF x =- 18910 THEN
            exp_f := 0;
        ELSIF x =- 18909 THEN
            exp_f := 0;
        ELSIF x =- 18908 THEN
            exp_f := 0;
        ELSIF x =- 18907 THEN
            exp_f := 0;
        ELSIF x =- 18906 THEN
            exp_f := 0;
        ELSIF x =- 18905 THEN
            exp_f := 0;
        ELSIF x =- 18904 THEN
            exp_f := 0;
        ELSIF x =- 18903 THEN
            exp_f := 0;
        ELSIF x =- 18902 THEN
            exp_f := 0;
        ELSIF x =- 18901 THEN
            exp_f := 0;
        ELSIF x =- 18900 THEN
            exp_f := 0;
        ELSIF x =- 18899 THEN
            exp_f := 0;
        ELSIF x =- 18898 THEN
            exp_f := 0;
        ELSIF x =- 18897 THEN
            exp_f := 0;
        ELSIF x =- 18896 THEN
            exp_f := 0;
        ELSIF x =- 18895 THEN
            exp_f := 0;
        ELSIF x =- 18894 THEN
            exp_f := 0;
        ELSIF x =- 18893 THEN
            exp_f := 0;
        ELSIF x =- 18892 THEN
            exp_f := 0;
        ELSIF x =- 18891 THEN
            exp_f := 0;
        ELSIF x =- 18890 THEN
            exp_f := 0;
        ELSIF x =- 18889 THEN
            exp_f := 0;
        ELSIF x =- 18888 THEN
            exp_f := 0;
        ELSIF x =- 18887 THEN
            exp_f := 0;
        ELSIF x =- 18886 THEN
            exp_f := 0;
        ELSIF x =- 18885 THEN
            exp_f := 0;
        ELSIF x =- 18884 THEN
            exp_f := 0;
        ELSIF x =- 18883 THEN
            exp_f := 0;
        ELSIF x =- 18882 THEN
            exp_f := 0;
        ELSIF x =- 18881 THEN
            exp_f := 0;
        ELSIF x =- 18880 THEN
            exp_f := 0;
        ELSIF x =- 18879 THEN
            exp_f := 0;
        ELSIF x =- 18878 THEN
            exp_f := 0;
        ELSIF x =- 18877 THEN
            exp_f := 0;
        ELSIF x =- 18876 THEN
            exp_f := 0;
        ELSIF x =- 18875 THEN
            exp_f := 0;
        ELSIF x =- 18874 THEN
            exp_f := 0;
        ELSIF x =- 18873 THEN
            exp_f := 0;
        ELSIF x =- 18872 THEN
            exp_f := 0;
        ELSIF x =- 18871 THEN
            exp_f := 0;
        ELSIF x =- 18870 THEN
            exp_f := 0;
        ELSIF x =- 18869 THEN
            exp_f := 0;
        ELSIF x =- 18868 THEN
            exp_f := 0;
        ELSIF x =- 18867 THEN
            exp_f := 0;
        ELSIF x =- 18866 THEN
            exp_f := 0;
        ELSIF x =- 18865 THEN
            exp_f := 0;
        ELSIF x =- 18864 THEN
            exp_f := 0;
        ELSIF x =- 18863 THEN
            exp_f := 0;
        ELSIF x =- 18862 THEN
            exp_f := 0;
        ELSIF x =- 18861 THEN
            exp_f := 0;
        ELSIF x =- 18860 THEN
            exp_f := 0;
        ELSIF x =- 18859 THEN
            exp_f := 0;
        ELSIF x =- 18858 THEN
            exp_f := 0;
        ELSIF x =- 18857 THEN
            exp_f := 0;
        ELSIF x =- 18856 THEN
            exp_f := 0;
        ELSIF x =- 18855 THEN
            exp_f := 0;
        ELSIF x =- 18854 THEN
            exp_f := 0;
        ELSIF x =- 18853 THEN
            exp_f := 0;
        ELSIF x =- 18852 THEN
            exp_f := 0;
        ELSIF x =- 18851 THEN
            exp_f := 0;
        ELSIF x =- 18850 THEN
            exp_f := 0;
        ELSIF x =- 18849 THEN
            exp_f := 0;
        ELSIF x =- 18848 THEN
            exp_f := 0;
        ELSIF x =- 18847 THEN
            exp_f := 0;
        ELSIF x =- 18846 THEN
            exp_f := 0;
        ELSIF x =- 18845 THEN
            exp_f := 0;
        ELSIF x =- 18844 THEN
            exp_f := 0;
        ELSIF x =- 18843 THEN
            exp_f := 0;
        ELSIF x =- 18842 THEN
            exp_f := 0;
        ELSIF x =- 18841 THEN
            exp_f := 0;
        ELSIF x =- 18840 THEN
            exp_f := 0;
        ELSIF x =- 18839 THEN
            exp_f := 0;
        ELSIF x =- 18838 THEN
            exp_f := 0;
        ELSIF x =- 18837 THEN
            exp_f := 0;
        ELSIF x =- 18836 THEN
            exp_f := 0;
        ELSIF x =- 18835 THEN
            exp_f := 0;
        ELSIF x =- 18834 THEN
            exp_f := 0;
        ELSIF x =- 18833 THEN
            exp_f := 0;
        ELSIF x =- 18832 THEN
            exp_f := 0;
        ELSIF x =- 18831 THEN
            exp_f := 0;
        ELSIF x =- 18830 THEN
            exp_f := 0;
        ELSIF x =- 18829 THEN
            exp_f := 0;
        ELSIF x =- 18828 THEN
            exp_f := 0;
        ELSIF x =- 18827 THEN
            exp_f := 0;
        ELSIF x =- 18826 THEN
            exp_f := 0;
        ELSIF x =- 18825 THEN
            exp_f := 0;
        ELSIF x =- 18824 THEN
            exp_f := 0;
        ELSIF x =- 18823 THEN
            exp_f := 0;
        ELSIF x =- 18822 THEN
            exp_f := 0;
        ELSIF x =- 18821 THEN
            exp_f := 0;
        ELSIF x =- 18820 THEN
            exp_f := 0;
        ELSIF x =- 18819 THEN
            exp_f := 0;
        ELSIF x =- 18818 THEN
            exp_f := 0;
        ELSIF x =- 18817 THEN
            exp_f := 0;
        ELSIF x =- 18816 THEN
            exp_f := 0;
        ELSIF x =- 18815 THEN
            exp_f := 0;
        ELSIF x =- 18814 THEN
            exp_f := 0;
        ELSIF x =- 18813 THEN
            exp_f := 0;
        ELSIF x =- 18812 THEN
            exp_f := 0;
        ELSIF x =- 18811 THEN
            exp_f := 0;
        ELSIF x =- 18810 THEN
            exp_f := 0;
        ELSIF x =- 18809 THEN
            exp_f := 0;
        ELSIF x =- 18808 THEN
            exp_f := 0;
        ELSIF x =- 18807 THEN
            exp_f := 0;
        ELSIF x =- 18806 THEN
            exp_f := 0;
        ELSIF x =- 18805 THEN
            exp_f := 0;
        ELSIF x =- 18804 THEN
            exp_f := 0;
        ELSIF x =- 18803 THEN
            exp_f := 0;
        ELSIF x =- 18802 THEN
            exp_f := 0;
        ELSIF x =- 18801 THEN
            exp_f := 0;
        ELSIF x =- 18800 THEN
            exp_f := 0;
        ELSIF x =- 18799 THEN
            exp_f := 0;
        ELSIF x =- 18798 THEN
            exp_f := 0;
        ELSIF x =- 18797 THEN
            exp_f := 0;
        ELSIF x =- 18796 THEN
            exp_f := 0;
        ELSIF x =- 18795 THEN
            exp_f := 0;
        ELSIF x =- 18794 THEN
            exp_f := 0;
        ELSIF x =- 18793 THEN
            exp_f := 0;
        ELSIF x =- 18792 THEN
            exp_f := 0;
        ELSIF x =- 18791 THEN
            exp_f := 0;
        ELSIF x =- 18790 THEN
            exp_f := 0;
        ELSIF x =- 18789 THEN
            exp_f := 0;
        ELSIF x =- 18788 THEN
            exp_f := 0;
        ELSIF x =- 18787 THEN
            exp_f := 0;
        ELSIF x =- 18786 THEN
            exp_f := 0;
        ELSIF x =- 18785 THEN
            exp_f := 0;
        ELSIF x =- 18784 THEN
            exp_f := 0;
        ELSIF x =- 18783 THEN
            exp_f := 0;
        ELSIF x =- 18782 THEN
            exp_f := 0;
        ELSIF x =- 18781 THEN
            exp_f := 0;
        ELSIF x =- 18780 THEN
            exp_f := 0;
        ELSIF x =- 18779 THEN
            exp_f := 0;
        ELSIF x =- 18778 THEN
            exp_f := 0;
        ELSIF x =- 18777 THEN
            exp_f := 0;
        ELSIF x =- 18776 THEN
            exp_f := 0;
        ELSIF x =- 18775 THEN
            exp_f := 0;
        ELSIF x =- 18774 THEN
            exp_f := 0;
        ELSIF x =- 18773 THEN
            exp_f := 0;
        ELSIF x =- 18772 THEN
            exp_f := 0;
        ELSIF x =- 18771 THEN
            exp_f := 0;
        ELSIF x =- 18770 THEN
            exp_f := 0;
        ELSIF x =- 18769 THEN
            exp_f := 0;
        ELSIF x =- 18768 THEN
            exp_f := 0;
        ELSIF x =- 18767 THEN
            exp_f := 0;
        ELSIF x =- 18766 THEN
            exp_f := 0;
        ELSIF x =- 18765 THEN
            exp_f := 0;
        ELSIF x =- 18764 THEN
            exp_f := 0;
        ELSIF x =- 18763 THEN
            exp_f := 0;
        ELSIF x =- 18762 THEN
            exp_f := 0;
        ELSIF x =- 18761 THEN
            exp_f := 0;
        ELSIF x =- 18760 THEN
            exp_f := 0;
        ELSIF x =- 18759 THEN
            exp_f := 0;
        ELSIF x =- 18758 THEN
            exp_f := 0;
        ELSIF x =- 18757 THEN
            exp_f := 0;
        ELSIF x =- 18756 THEN
            exp_f := 0;
        ELSIF x =- 18755 THEN
            exp_f := 0;
        ELSIF x =- 18754 THEN
            exp_f := 0;
        ELSIF x =- 18753 THEN
            exp_f := 0;
        ELSIF x =- 18752 THEN
            exp_f := 0;
        ELSIF x =- 18751 THEN
            exp_f := 0;
        ELSIF x =- 18750 THEN
            exp_f := 0;
        ELSIF x =- 18749 THEN
            exp_f := 0;
        ELSIF x =- 18748 THEN
            exp_f := 0;
        ELSIF x =- 18747 THEN
            exp_f := 0;
        ELSIF x =- 18746 THEN
            exp_f := 0;
        ELSIF x =- 18745 THEN
            exp_f := 0;
        ELSIF x =- 18744 THEN
            exp_f := 0;
        ELSIF x =- 18743 THEN
            exp_f := 0;
        ELSIF x =- 18742 THEN
            exp_f := 0;
        ELSIF x =- 18741 THEN
            exp_f := 0;
        ELSIF x =- 18740 THEN
            exp_f := 0;
        ELSIF x =- 18739 THEN
            exp_f := 0;
        ELSIF x =- 18738 THEN
            exp_f := 0;
        ELSIF x =- 18737 THEN
            exp_f := 0;
        ELSIF x =- 18736 THEN
            exp_f := 0;
        ELSIF x =- 18735 THEN
            exp_f := 0;
        ELSIF x =- 18734 THEN
            exp_f := 0;
        ELSIF x =- 18733 THEN
            exp_f := 0;
        ELSIF x =- 18732 THEN
            exp_f := 0;
        ELSIF x =- 18731 THEN
            exp_f := 0;
        ELSIF x =- 18730 THEN
            exp_f := 0;
        ELSIF x =- 18729 THEN
            exp_f := 0;
        ELSIF x =- 18728 THEN
            exp_f := 0;
        ELSIF x =- 18727 THEN
            exp_f := 0;
        ELSIF x =- 18726 THEN
            exp_f := 0;
        ELSIF x =- 18725 THEN
            exp_f := 0;
        ELSIF x =- 18724 THEN
            exp_f := 0;
        ELSIF x =- 18723 THEN
            exp_f := 0;
        ELSIF x =- 18722 THEN
            exp_f := 0;
        ELSIF x =- 18721 THEN
            exp_f := 0;
        ELSIF x =- 18720 THEN
            exp_f := 0;
        ELSIF x =- 18719 THEN
            exp_f := 0;
        ELSIF x =- 18718 THEN
            exp_f := 0;
        ELSIF x =- 18717 THEN
            exp_f := 0;
        ELSIF x =- 18716 THEN
            exp_f := 0;
        ELSIF x =- 18715 THEN
            exp_f := 0;
        ELSIF x =- 18714 THEN
            exp_f := 0;
        ELSIF x =- 18713 THEN
            exp_f := 0;
        ELSIF x =- 18712 THEN
            exp_f := 0;
        ELSIF x =- 18711 THEN
            exp_f := 0;
        ELSIF x =- 18710 THEN
            exp_f := 0;
        ELSIF x =- 18709 THEN
            exp_f := 0;
        ELSIF x =- 18708 THEN
            exp_f := 0;
        ELSIF x =- 18707 THEN
            exp_f := 0;
        ELSIF x =- 18706 THEN
            exp_f := 0;
        ELSIF x =- 18705 THEN
            exp_f := 0;
        ELSIF x =- 18704 THEN
            exp_f := 0;
        ELSIF x =- 18703 THEN
            exp_f := 0;
        ELSIF x =- 18702 THEN
            exp_f := 0;
        ELSIF x =- 18701 THEN
            exp_f := 0;
        ELSIF x =- 18700 THEN
            exp_f := 0;
        ELSIF x =- 18699 THEN
            exp_f := 0;
        ELSIF x =- 18698 THEN
            exp_f := 0;
        ELSIF x =- 18697 THEN
            exp_f := 0;
        ELSIF x =- 18696 THEN
            exp_f := 0;
        ELSIF x =- 18695 THEN
            exp_f := 0;
        ELSIF x =- 18694 THEN
            exp_f := 0;
        ELSIF x =- 18693 THEN
            exp_f := 0;
        ELSIF x =- 18692 THEN
            exp_f := 0;
        ELSIF x =- 18691 THEN
            exp_f := 0;
        ELSIF x =- 18690 THEN
            exp_f := 0;
        ELSIF x =- 18689 THEN
            exp_f := 0;
        ELSIF x =- 18688 THEN
            exp_f := 0;
        ELSIF x =- 18687 THEN
            exp_f := 0;
        ELSIF x =- 18686 THEN
            exp_f := 0;
        ELSIF x =- 18685 THEN
            exp_f := 0;
        ELSIF x =- 18684 THEN
            exp_f := 0;
        ELSIF x =- 18683 THEN
            exp_f := 0;
        ELSIF x =- 18682 THEN
            exp_f := 0;
        ELSIF x =- 18681 THEN
            exp_f := 0;
        ELSIF x =- 18680 THEN
            exp_f := 0;
        ELSIF x =- 18679 THEN
            exp_f := 0;
        ELSIF x =- 18678 THEN
            exp_f := 0;
        ELSIF x =- 18677 THEN
            exp_f := 0;
        ELSIF x =- 18676 THEN
            exp_f := 0;
        ELSIF x =- 18675 THEN
            exp_f := 0;
        ELSIF x =- 18674 THEN
            exp_f := 0;
        ELSIF x =- 18673 THEN
            exp_f := 0;
        ELSIF x =- 18672 THEN
            exp_f := 0;
        ELSIF x =- 18671 THEN
            exp_f := 0;
        ELSIF x =- 18670 THEN
            exp_f := 0;
        ELSIF x =- 18669 THEN
            exp_f := 0;
        ELSIF x =- 18668 THEN
            exp_f := 0;
        ELSIF x =- 18667 THEN
            exp_f := 0;
        ELSIF x =- 18666 THEN
            exp_f := 0;
        ELSIF x =- 18665 THEN
            exp_f := 0;
        ELSIF x =- 18664 THEN
            exp_f := 0;
        ELSIF x =- 18663 THEN
            exp_f := 0;
        ELSIF x =- 18662 THEN
            exp_f := 0;
        ELSIF x =- 18661 THEN
            exp_f := 0;
        ELSIF x =- 18660 THEN
            exp_f := 0;
        ELSIF x =- 18659 THEN
            exp_f := 0;
        ELSIF x =- 18658 THEN
            exp_f := 0;
        ELSIF x =- 18657 THEN
            exp_f := 0;
        ELSIF x =- 18656 THEN
            exp_f := 0;
        ELSIF x =- 18655 THEN
            exp_f := 0;
        ELSIF x =- 18654 THEN
            exp_f := 0;
        ELSIF x =- 18653 THEN
            exp_f := 0;
        ELSIF x =- 18652 THEN
            exp_f := 0;
        ELSIF x =- 18651 THEN
            exp_f := 0;
        ELSIF x =- 18650 THEN
            exp_f := 0;
        ELSIF x =- 18649 THEN
            exp_f := 0;
        ELSIF x =- 18648 THEN
            exp_f := 0;
        ELSIF x =- 18647 THEN
            exp_f := 0;
        ELSIF x =- 18646 THEN
            exp_f := 0;
        ELSIF x =- 18645 THEN
            exp_f := 0;
        ELSIF x =- 18644 THEN
            exp_f := 0;
        ELSIF x =- 18643 THEN
            exp_f := 0;
        ELSIF x =- 18642 THEN
            exp_f := 0;
        ELSIF x =- 18641 THEN
            exp_f := 0;
        ELSIF x =- 18640 THEN
            exp_f := 0;
        ELSIF x =- 18639 THEN
            exp_f := 0;
        ELSIF x =- 18638 THEN
            exp_f := 0;
        ELSIF x =- 18637 THEN
            exp_f := 0;
        ELSIF x =- 18636 THEN
            exp_f := 0;
        ELSIF x =- 18635 THEN
            exp_f := 0;
        ELSIF x =- 18634 THEN
            exp_f := 0;
        ELSIF x =- 18633 THEN
            exp_f := 0;
        ELSIF x =- 18632 THEN
            exp_f := 0;
        ELSIF x =- 18631 THEN
            exp_f := 0;
        ELSIF x =- 18630 THEN
            exp_f := 0;
        ELSIF x =- 18629 THEN
            exp_f := 0;
        ELSIF x =- 18628 THEN
            exp_f := 0;
        ELSIF x =- 18627 THEN
            exp_f := 0;
        ELSIF x =- 18626 THEN
            exp_f := 0;
        ELSIF x =- 18625 THEN
            exp_f := 0;
        ELSIF x =- 18624 THEN
            exp_f := 0;
        ELSIF x =- 18623 THEN
            exp_f := 0;
        ELSIF x =- 18622 THEN
            exp_f := 0;
        ELSIF x =- 18621 THEN
            exp_f := 0;
        ELSIF x =- 18620 THEN
            exp_f := 0;
        ELSIF x =- 18619 THEN
            exp_f := 0;
        ELSIF x =- 18618 THEN
            exp_f := 0;
        ELSIF x =- 18617 THEN
            exp_f := 0;
        ELSIF x =- 18616 THEN
            exp_f := 0;
        ELSIF x =- 18615 THEN
            exp_f := 0;
        ELSIF x =- 18614 THEN
            exp_f := 0;
        ELSIF x =- 18613 THEN
            exp_f := 0;
        ELSIF x =- 18612 THEN
            exp_f := 0;
        ELSIF x =- 18611 THEN
            exp_f := 0;
        ELSIF x =- 18610 THEN
            exp_f := 0;
        ELSIF x =- 18609 THEN
            exp_f := 0;
        ELSIF x =- 18608 THEN
            exp_f := 0;
        ELSIF x =- 18607 THEN
            exp_f := 0;
        ELSIF x =- 18606 THEN
            exp_f := 0;
        ELSIF x =- 18605 THEN
            exp_f := 0;
        ELSIF x =- 18604 THEN
            exp_f := 0;
        ELSIF x =- 18603 THEN
            exp_f := 0;
        ELSIF x =- 18602 THEN
            exp_f := 0;
        ELSIF x =- 18601 THEN
            exp_f := 0;
        ELSIF x =- 18600 THEN
            exp_f := 0;
        ELSIF x =- 18599 THEN
            exp_f := 0;
        ELSIF x =- 18598 THEN
            exp_f := 0;
        ELSIF x =- 18597 THEN
            exp_f := 0;
        ELSIF x =- 18596 THEN
            exp_f := 0;
        ELSIF x =- 18595 THEN
            exp_f := 0;
        ELSIF x =- 18594 THEN
            exp_f := 0;
        ELSIF x =- 18593 THEN
            exp_f := 0;
        ELSIF x =- 18592 THEN
            exp_f := 0;
        ELSIF x =- 18591 THEN
            exp_f := 0;
        ELSIF x =- 18590 THEN
            exp_f := 0;
        ELSIF x =- 18589 THEN
            exp_f := 0;
        ELSIF x =- 18588 THEN
            exp_f := 0;
        ELSIF x =- 18587 THEN
            exp_f := 0;
        ELSIF x =- 18586 THEN
            exp_f := 0;
        ELSIF x =- 18585 THEN
            exp_f := 0;
        ELSIF x =- 18584 THEN
            exp_f := 0;
        ELSIF x =- 18583 THEN
            exp_f := 0;
        ELSIF x =- 18582 THEN
            exp_f := 0;
        ELSIF x =- 18581 THEN
            exp_f := 0;
        ELSIF x =- 18580 THEN
            exp_f := 0;
        ELSIF x =- 18579 THEN
            exp_f := 0;
        ELSIF x =- 18578 THEN
            exp_f := 0;
        ELSIF x =- 18577 THEN
            exp_f := 0;
        ELSIF x =- 18576 THEN
            exp_f := 0;
        ELSIF x =- 18575 THEN
            exp_f := 0;
        ELSIF x =- 18574 THEN
            exp_f := 0;
        ELSIF x =- 18573 THEN
            exp_f := 0;
        ELSIF x =- 18572 THEN
            exp_f := 0;
        ELSIF x =- 18571 THEN
            exp_f := 0;
        ELSIF x =- 18570 THEN
            exp_f := 0;
        ELSIF x =- 18569 THEN
            exp_f := 0;
        ELSIF x =- 18568 THEN
            exp_f := 0;
        ELSIF x =- 18567 THEN
            exp_f := 0;
        ELSIF x =- 18566 THEN
            exp_f := 0;
        ELSIF x =- 18565 THEN
            exp_f := 0;
        ELSIF x =- 18564 THEN
            exp_f := 0;
        ELSIF x =- 18563 THEN
            exp_f := 0;
        ELSIF x =- 18562 THEN
            exp_f := 0;
        ELSIF x =- 18561 THEN
            exp_f := 0;
        ELSIF x =- 18560 THEN
            exp_f := 0;
        ELSIF x =- 18559 THEN
            exp_f := 0;
        ELSIF x =- 18558 THEN
            exp_f := 0;
        ELSIF x =- 18557 THEN
            exp_f := 0;
        ELSIF x =- 18556 THEN
            exp_f := 0;
        ELSIF x =- 18555 THEN
            exp_f := 0;
        ELSIF x =- 18554 THEN
            exp_f := 0;
        ELSIF x =- 18553 THEN
            exp_f := 0;
        ELSIF x =- 18552 THEN
            exp_f := 0;
        ELSIF x =- 18551 THEN
            exp_f := 0;
        ELSIF x =- 18550 THEN
            exp_f := 0;
        ELSIF x =- 18549 THEN
            exp_f := 0;
        ELSIF x =- 18548 THEN
            exp_f := 0;
        ELSIF x =- 18547 THEN
            exp_f := 0;
        ELSIF x =- 18546 THEN
            exp_f := 0;
        ELSIF x =- 18545 THEN
            exp_f := 0;
        ELSIF x =- 18544 THEN
            exp_f := 0;
        ELSIF x =- 18543 THEN
            exp_f := 0;
        ELSIF x =- 18542 THEN
            exp_f := 0;
        ELSIF x =- 18541 THEN
            exp_f := 0;
        ELSIF x =- 18540 THEN
            exp_f := 0;
        ELSIF x =- 18539 THEN
            exp_f := 0;
        ELSIF x =- 18538 THEN
            exp_f := 0;
        ELSIF x =- 18537 THEN
            exp_f := 0;
        ELSIF x =- 18536 THEN
            exp_f := 0;
        ELSIF x =- 18535 THEN
            exp_f := 0;
        ELSIF x =- 18534 THEN
            exp_f := 0;
        ELSIF x =- 18533 THEN
            exp_f := 0;
        ELSIF x =- 18532 THEN
            exp_f := 0;
        ELSIF x =- 18531 THEN
            exp_f := 0;
        ELSIF x =- 18530 THEN
            exp_f := 0;
        ELSIF x =- 18529 THEN
            exp_f := 0;
        ELSIF x =- 18528 THEN
            exp_f := 0;
        ELSIF x =- 18527 THEN
            exp_f := 0;
        ELSIF x =- 18526 THEN
            exp_f := 0;
        ELSIF x =- 18525 THEN
            exp_f := 0;
        ELSIF x =- 18524 THEN
            exp_f := 0;
        ELSIF x =- 18523 THEN
            exp_f := 0;
        ELSIF x =- 18522 THEN
            exp_f := 0;
        ELSIF x =- 18521 THEN
            exp_f := 0;
        ELSIF x =- 18520 THEN
            exp_f := 0;
        ELSIF x =- 18519 THEN
            exp_f := 0;
        ELSIF x =- 18518 THEN
            exp_f := 0;
        ELSIF x =- 18517 THEN
            exp_f := 0;
        ELSIF x =- 18516 THEN
            exp_f := 0;
        ELSIF x =- 18515 THEN
            exp_f := 0;
        ELSIF x =- 18514 THEN
            exp_f := 0;
        ELSIF x =- 18513 THEN
            exp_f := 0;
        ELSIF x =- 18512 THEN
            exp_f := 0;
        ELSIF x =- 18511 THEN
            exp_f := 0;
        ELSIF x =- 18510 THEN
            exp_f := 0;
        ELSIF x =- 18509 THEN
            exp_f := 0;
        ELSIF x =- 18508 THEN
            exp_f := 0;
        ELSIF x =- 18507 THEN
            exp_f := 0;
        ELSIF x =- 18506 THEN
            exp_f := 0;
        ELSIF x =- 18505 THEN
            exp_f := 0;
        ELSIF x =- 18504 THEN
            exp_f := 0;
        ELSIF x =- 18503 THEN
            exp_f := 0;
        ELSIF x =- 18502 THEN
            exp_f := 0;
        ELSIF x =- 18501 THEN
            exp_f := 0;
        ELSIF x =- 18500 THEN
            exp_f := 0;
        ELSIF x =- 18499 THEN
            exp_f := 0;
        ELSIF x =- 18498 THEN
            exp_f := 0;
        ELSIF x =- 18497 THEN
            exp_f := 0;
        ELSIF x =- 18496 THEN
            exp_f := 0;
        ELSIF x =- 18495 THEN
            exp_f := 0;
        ELSIF x =- 18494 THEN
            exp_f := 0;
        ELSIF x =- 18493 THEN
            exp_f := 0;
        ELSIF x =- 18492 THEN
            exp_f := 0;
        ELSIF x =- 18491 THEN
            exp_f := 0;
        ELSIF x =- 18490 THEN
            exp_f := 0;
        ELSIF x =- 18489 THEN
            exp_f := 0;
        ELSIF x =- 18488 THEN
            exp_f := 0;
        ELSIF x =- 18487 THEN
            exp_f := 0;
        ELSIF x =- 18486 THEN
            exp_f := 0;
        ELSIF x =- 18485 THEN
            exp_f := 0;
        ELSIF x =- 18484 THEN
            exp_f := 0;
        ELSIF x =- 18483 THEN
            exp_f := 0;
        ELSIF x =- 18482 THEN
            exp_f := 0;
        ELSIF x =- 18481 THEN
            exp_f := 0;
        ELSIF x =- 18480 THEN
            exp_f := 0;
        ELSIF x =- 18479 THEN
            exp_f := 0;
        ELSIF x =- 18478 THEN
            exp_f := 0;
        ELSIF x =- 18477 THEN
            exp_f := 0;
        ELSIF x =- 18476 THEN
            exp_f := 0;
        ELSIF x =- 18475 THEN
            exp_f := 0;
        ELSIF x =- 18474 THEN
            exp_f := 0;
        ELSIF x =- 18473 THEN
            exp_f := 0;
        ELSIF x =- 18472 THEN
            exp_f := 0;
        ELSIF x =- 18471 THEN
            exp_f := 0;
        ELSIF x =- 18470 THEN
            exp_f := 0;
        ELSIF x =- 18469 THEN
            exp_f := 0;
        ELSIF x =- 18468 THEN
            exp_f := 0;
        ELSIF x =- 18467 THEN
            exp_f := 0;
        ELSIF x =- 18466 THEN
            exp_f := 0;
        ELSIF x =- 18465 THEN
            exp_f := 0;
        ELSIF x =- 18464 THEN
            exp_f := 0;
        ELSIF x =- 18463 THEN
            exp_f := 0;
        ELSIF x =- 18462 THEN
            exp_f := 0;
        ELSIF x =- 18461 THEN
            exp_f := 0;
        ELSIF x =- 18460 THEN
            exp_f := 0;
        ELSIF x =- 18459 THEN
            exp_f := 0;
        ELSIF x =- 18458 THEN
            exp_f := 0;
        ELSIF x =- 18457 THEN
            exp_f := 0;
        ELSIF x =- 18456 THEN
            exp_f := 0;
        ELSIF x =- 18455 THEN
            exp_f := 0;
        ELSIF x =- 18454 THEN
            exp_f := 0;
        ELSIF x =- 18453 THEN
            exp_f := 0;
        ELSIF x =- 18452 THEN
            exp_f := 0;
        ELSIF x =- 18451 THEN
            exp_f := 0;
        ELSIF x =- 18450 THEN
            exp_f := 0;
        ELSIF x =- 18449 THEN
            exp_f := 0;
        ELSIF x =- 18448 THEN
            exp_f := 0;
        ELSIF x =- 18447 THEN
            exp_f := 0;
        ELSIF x =- 18446 THEN
            exp_f := 0;
        ELSIF x =- 18445 THEN
            exp_f := 0;
        ELSIF x =- 18444 THEN
            exp_f := 0;
        ELSIF x =- 18443 THEN
            exp_f := 0;
        ELSIF x =- 18442 THEN
            exp_f := 0;
        ELSIF x =- 18441 THEN
            exp_f := 0;
        ELSIF x =- 18440 THEN
            exp_f := 0;
        ELSIF x =- 18439 THEN
            exp_f := 0;
        ELSIF x =- 18438 THEN
            exp_f := 0;
        ELSIF x =- 18437 THEN
            exp_f := 0;
        ELSIF x =- 18436 THEN
            exp_f := 0;
        ELSIF x =- 18435 THEN
            exp_f := 0;
        ELSIF x =- 18434 THEN
            exp_f := 0;
        ELSIF x =- 18433 THEN
            exp_f := 0;
        ELSIF x =- 18432 THEN
            exp_f := 0;
        ELSIF x =- 18431 THEN
            exp_f := 0;
        ELSIF x =- 18430 THEN
            exp_f := 0;
        ELSIF x =- 18429 THEN
            exp_f := 0;
        ELSIF x =- 18428 THEN
            exp_f := 0;
        ELSIF x =- 18427 THEN
            exp_f := 0;
        ELSIF x =- 18426 THEN
            exp_f := 0;
        ELSIF x =- 18425 THEN
            exp_f := 0;
        ELSIF x =- 18424 THEN
            exp_f := 0;
        ELSIF x =- 18423 THEN
            exp_f := 0;
        ELSIF x =- 18422 THEN
            exp_f := 0;
        ELSIF x =- 18421 THEN
            exp_f := 0;
        ELSIF x =- 18420 THEN
            exp_f := 0;
        ELSIF x =- 18419 THEN
            exp_f := 0;
        ELSIF x =- 18418 THEN
            exp_f := 0;
        ELSIF x =- 18417 THEN
            exp_f := 0;
        ELSIF x =- 18416 THEN
            exp_f := 0;
        ELSIF x =- 18415 THEN
            exp_f := 0;
        ELSIF x =- 18414 THEN
            exp_f := 0;
        ELSIF x =- 18413 THEN
            exp_f := 0;
        ELSIF x =- 18412 THEN
            exp_f := 0;
        ELSIF x =- 18411 THEN
            exp_f := 0;
        ELSIF x =- 18410 THEN
            exp_f := 0;
        ELSIF x =- 18409 THEN
            exp_f := 0;
        ELSIF x =- 18408 THEN
            exp_f := 0;
        ELSIF x =- 18407 THEN
            exp_f := 0;
        ELSIF x =- 18406 THEN
            exp_f := 0;
        ELSIF x =- 18405 THEN
            exp_f := 0;
        ELSIF x =- 18404 THEN
            exp_f := 0;
        ELSIF x =- 18403 THEN
            exp_f := 0;
        ELSIF x =- 18402 THEN
            exp_f := 0;
        ELSIF x =- 18401 THEN
            exp_f := 0;
        ELSIF x =- 18400 THEN
            exp_f := 0;
        ELSIF x =- 18399 THEN
            exp_f := 0;
        ELSIF x =- 18398 THEN
            exp_f := 0;
        ELSIF x =- 18397 THEN
            exp_f := 0;
        ELSIF x =- 18396 THEN
            exp_f := 0;
        ELSIF x =- 18395 THEN
            exp_f := 0;
        ELSIF x =- 18394 THEN
            exp_f := 0;
        ELSIF x =- 18393 THEN
            exp_f := 0;
        ELSIF x =- 18392 THEN
            exp_f := 0;
        ELSIF x =- 18391 THEN
            exp_f := 0;
        ELSIF x =- 18390 THEN
            exp_f := 0;
        ELSIF x =- 18389 THEN
            exp_f := 0;
        ELSIF x =- 18388 THEN
            exp_f := 0;
        ELSIF x =- 18387 THEN
            exp_f := 0;
        ELSIF x =- 18386 THEN
            exp_f := 0;
        ELSIF x =- 18385 THEN
            exp_f := 0;
        ELSIF x =- 18384 THEN
            exp_f := 0;
        ELSIF x =- 18383 THEN
            exp_f := 0;
        ELSIF x =- 18382 THEN
            exp_f := 0;
        ELSIF x =- 18381 THEN
            exp_f := 0;
        ELSIF x =- 18380 THEN
            exp_f := 0;
        ELSIF x =- 18379 THEN
            exp_f := 0;
        ELSIF x =- 18378 THEN
            exp_f := 0;
        ELSIF x =- 18377 THEN
            exp_f := 0;
        ELSIF x =- 18376 THEN
            exp_f := 0;
        ELSIF x =- 18375 THEN
            exp_f := 0;
        ELSIF x =- 18374 THEN
            exp_f := 0;
        ELSIF x =- 18373 THEN
            exp_f := 0;
        ELSIF x =- 18372 THEN
            exp_f := 0;
        ELSIF x =- 18371 THEN
            exp_f := 0;
        ELSIF x =- 18370 THEN
            exp_f := 0;
        ELSIF x =- 18369 THEN
            exp_f := 0;
        ELSIF x =- 18368 THEN
            exp_f := 0;
        ELSIF x =- 18367 THEN
            exp_f := 0;
        ELSIF x =- 18366 THEN
            exp_f := 0;
        ELSIF x =- 18365 THEN
            exp_f := 0;
        ELSIF x =- 18364 THEN
            exp_f := 0;
        ELSIF x =- 18363 THEN
            exp_f := 0;
        ELSIF x =- 18362 THEN
            exp_f := 0;
        ELSIF x =- 18361 THEN
            exp_f := 0;
        ELSIF x =- 18360 THEN
            exp_f := 0;
        ELSIF x =- 18359 THEN
            exp_f := 0;
        ELSIF x =- 18358 THEN
            exp_f := 0;
        ELSIF x =- 18357 THEN
            exp_f := 0;
        ELSIF x =- 18356 THEN
            exp_f := 0;
        ELSIF x =- 18355 THEN
            exp_f := 0;
        ELSIF x =- 18354 THEN
            exp_f := 0;
        ELSIF x =- 18353 THEN
            exp_f := 0;
        ELSIF x =- 18352 THEN
            exp_f := 0;
        ELSIF x =- 18351 THEN
            exp_f := 0;
        ELSIF x =- 18350 THEN
            exp_f := 0;
        ELSIF x =- 18349 THEN
            exp_f := 0;
        ELSIF x =- 18348 THEN
            exp_f := 0;
        ELSIF x =- 18347 THEN
            exp_f := 0;
        ELSIF x =- 18346 THEN
            exp_f := 0;
        ELSIF x =- 18345 THEN
            exp_f := 0;
        ELSIF x =- 18344 THEN
            exp_f := 0;
        ELSIF x =- 18343 THEN
            exp_f := 0;
        ELSIF x =- 18342 THEN
            exp_f := 0;
        ELSIF x =- 18341 THEN
            exp_f := 0;
        ELSIF x =- 18340 THEN
            exp_f := 0;
        ELSIF x =- 18339 THEN
            exp_f := 0;
        ELSIF x =- 18338 THEN
            exp_f := 0;
        ELSIF x =- 18337 THEN
            exp_f := 0;
        ELSIF x =- 18336 THEN
            exp_f := 0;
        ELSIF x =- 18335 THEN
            exp_f := 0;
        ELSIF x =- 18334 THEN
            exp_f := 0;
        ELSIF x =- 18333 THEN
            exp_f := 0;
        ELSIF x =- 18332 THEN
            exp_f := 0;
        ELSIF x =- 18331 THEN
            exp_f := 0;
        ELSIF x =- 18330 THEN
            exp_f := 0;
        ELSIF x =- 18329 THEN
            exp_f := 0;
        ELSIF x =- 18328 THEN
            exp_f := 0;
        ELSIF x =- 18327 THEN
            exp_f := 0;
        ELSIF x =- 18326 THEN
            exp_f := 0;
        ELSIF x =- 18325 THEN
            exp_f := 0;
        ELSIF x =- 18324 THEN
            exp_f := 0;
        ELSIF x =- 18323 THEN
            exp_f := 0;
        ELSIF x =- 18322 THEN
            exp_f := 0;
        ELSIF x =- 18321 THEN
            exp_f := 0;
        ELSIF x =- 18320 THEN
            exp_f := 0;
        ELSIF x =- 18319 THEN
            exp_f := 0;
        ELSIF x =- 18318 THEN
            exp_f := 0;
        ELSIF x =- 18317 THEN
            exp_f := 0;
        ELSIF x =- 18316 THEN
            exp_f := 0;
        ELSIF x =- 18315 THEN
            exp_f := 0;
        ELSIF x =- 18314 THEN
            exp_f := 0;
        ELSIF x =- 18313 THEN
            exp_f := 0;
        ELSIF x =- 18312 THEN
            exp_f := 0;
        ELSIF x =- 18311 THEN
            exp_f := 0;
        ELSIF x =- 18310 THEN
            exp_f := 0;
        ELSIF x =- 18309 THEN
            exp_f := 0;
        ELSIF x =- 18308 THEN
            exp_f := 0;
        ELSIF x =- 18307 THEN
            exp_f := 0;
        ELSIF x =- 18306 THEN
            exp_f := 0;
        ELSIF x =- 18305 THEN
            exp_f := 0;
        ELSIF x =- 18304 THEN
            exp_f := 0;
        ELSIF x =- 18303 THEN
            exp_f := 0;
        ELSIF x =- 18302 THEN
            exp_f := 0;
        ELSIF x =- 18301 THEN
            exp_f := 0;
        ELSIF x =- 18300 THEN
            exp_f := 0;
        ELSIF x =- 18299 THEN
            exp_f := 0;
        ELSIF x =- 18298 THEN
            exp_f := 0;
        ELSIF x =- 18297 THEN
            exp_f := 0;
        ELSIF x =- 18296 THEN
            exp_f := 0;
        ELSIF x =- 18295 THEN
            exp_f := 0;
        ELSIF x =- 18294 THEN
            exp_f := 0;
        ELSIF x =- 18293 THEN
            exp_f := 0;
        ELSIF x =- 18292 THEN
            exp_f := 0;
        ELSIF x =- 18291 THEN
            exp_f := 0;
        ELSIF x =- 18290 THEN
            exp_f := 0;
        ELSIF x =- 18289 THEN
            exp_f := 0;
        ELSIF x =- 18288 THEN
            exp_f := 0;
        ELSIF x =- 18287 THEN
            exp_f := 0;
        ELSIF x =- 18286 THEN
            exp_f := 0;
        ELSIF x =- 18285 THEN
            exp_f := 0;
        ELSIF x =- 18284 THEN
            exp_f := 0;
        ELSIF x =- 18283 THEN
            exp_f := 0;
        ELSIF x =- 18282 THEN
            exp_f := 0;
        ELSIF x =- 18281 THEN
            exp_f := 0;
        ELSIF x =- 18280 THEN
            exp_f := 0;
        ELSIF x =- 18279 THEN
            exp_f := 0;
        ELSIF x =- 18278 THEN
            exp_f := 0;
        ELSIF x =- 18277 THEN
            exp_f := 0;
        ELSIF x =- 18276 THEN
            exp_f := 0;
        ELSIF x =- 18275 THEN
            exp_f := 0;
        ELSIF x =- 18274 THEN
            exp_f := 0;
        ELSIF x =- 18273 THEN
            exp_f := 0;
        ELSIF x =- 18272 THEN
            exp_f := 0;
        ELSIF x =- 18271 THEN
            exp_f := 0;
        ELSIF x =- 18270 THEN
            exp_f := 0;
        ELSIF x =- 18269 THEN
            exp_f := 0;
        ELSIF x =- 18268 THEN
            exp_f := 0;
        ELSIF x =- 18267 THEN
            exp_f := 0;
        ELSIF x =- 18266 THEN
            exp_f := 0;
        ELSIF x =- 18265 THEN
            exp_f := 0;
        ELSIF x =- 18264 THEN
            exp_f := 0;
        ELSIF x =- 18263 THEN
            exp_f := 0;
        ELSIF x =- 18262 THEN
            exp_f := 0;
        ELSIF x =- 18261 THEN
            exp_f := 0;
        ELSIF x =- 18260 THEN
            exp_f := 0;
        ELSIF x =- 18259 THEN
            exp_f := 0;
        ELSIF x =- 18258 THEN
            exp_f := 0;
        ELSIF x =- 18257 THEN
            exp_f := 0;
        ELSIF x =- 18256 THEN
            exp_f := 0;
        ELSIF x =- 18255 THEN
            exp_f := 0;
        ELSIF x =- 18254 THEN
            exp_f := 0;
        ELSIF x =- 18253 THEN
            exp_f := 0;
        ELSIF x =- 18252 THEN
            exp_f := 0;
        ELSIF x =- 18251 THEN
            exp_f := 0;
        ELSIF x =- 18250 THEN
            exp_f := 0;
        ELSIF x =- 18249 THEN
            exp_f := 0;
        ELSIF x =- 18248 THEN
            exp_f := 0;
        ELSIF x =- 18247 THEN
            exp_f := 0;
        ELSIF x =- 18246 THEN
            exp_f := 0;
        ELSIF x =- 18245 THEN
            exp_f := 0;
        ELSIF x =- 18244 THEN
            exp_f := 0;
        ELSIF x =- 18243 THEN
            exp_f := 0;
        ELSIF x =- 18242 THEN
            exp_f := 0;
        ELSIF x =- 18241 THEN
            exp_f := 0;
        ELSIF x =- 18240 THEN
            exp_f := 0;
        ELSIF x =- 18239 THEN
            exp_f := 0;
        ELSIF x =- 18238 THEN
            exp_f := 0;
        ELSIF x =- 18237 THEN
            exp_f := 0;
        ELSIF x =- 18236 THEN
            exp_f := 0;
        ELSIF x =- 18235 THEN
            exp_f := 0;
        ELSIF x =- 18234 THEN
            exp_f := 0;
        ELSIF x =- 18233 THEN
            exp_f := 0;
        ELSIF x =- 18232 THEN
            exp_f := 0;
        ELSIF x =- 18231 THEN
            exp_f := 0;
        ELSIF x =- 18230 THEN
            exp_f := 0;
        ELSIF x =- 18229 THEN
            exp_f := 0;
        ELSIF x =- 18228 THEN
            exp_f := 0;
        ELSIF x =- 18227 THEN
            exp_f := 0;
        ELSIF x =- 18226 THEN
            exp_f := 0;
        ELSIF x =- 18225 THEN
            exp_f := 0;
        ELSIF x =- 18224 THEN
            exp_f := 0;
        ELSIF x =- 18223 THEN
            exp_f := 0;
        ELSIF x =- 18222 THEN
            exp_f := 0;
        ELSIF x =- 18221 THEN
            exp_f := 0;
        ELSIF x =- 18220 THEN
            exp_f := 0;
        ELSIF x =- 18219 THEN
            exp_f := 0;
        ELSIF x =- 18218 THEN
            exp_f := 0;
        ELSIF x =- 18217 THEN
            exp_f := 0;
        ELSIF x =- 18216 THEN
            exp_f := 0;
        ELSIF x =- 18215 THEN
            exp_f := 0;
        ELSIF x =- 18214 THEN
            exp_f := 0;
        ELSIF x =- 18213 THEN
            exp_f := 0;
        ELSIF x =- 18212 THEN
            exp_f := 0;
        ELSIF x =- 18211 THEN
            exp_f := 0;
        ELSIF x =- 18210 THEN
            exp_f := 0;
        ELSIF x =- 18209 THEN
            exp_f := 0;
        ELSIF x =- 18208 THEN
            exp_f := 0;
        ELSIF x =- 18207 THEN
            exp_f := 0;
        ELSIF x =- 18206 THEN
            exp_f := 0;
        ELSIF x =- 18205 THEN
            exp_f := 0;
        ELSIF x =- 18204 THEN
            exp_f := 0;
        ELSIF x =- 18203 THEN
            exp_f := 0;
        ELSIF x =- 18202 THEN
            exp_f := 0;
        ELSIF x =- 18201 THEN
            exp_f := 0;
        ELSIF x =- 18200 THEN
            exp_f := 0;
        ELSIF x =- 18199 THEN
            exp_f := 0;
        ELSIF x =- 18198 THEN
            exp_f := 0;
        ELSIF x =- 18197 THEN
            exp_f := 0;
        ELSIF x =- 18196 THEN
            exp_f := 0;
        ELSIF x =- 18195 THEN
            exp_f := 0;
        ELSIF x =- 18194 THEN
            exp_f := 0;
        ELSIF x =- 18193 THEN
            exp_f := 0;
        ELSIF x =- 18192 THEN
            exp_f := 0;
        ELSIF x =- 18191 THEN
            exp_f := 0;
        ELSIF x =- 18190 THEN
            exp_f := 0;
        ELSIF x =- 18189 THEN
            exp_f := 0;
        ELSIF x =- 18188 THEN
            exp_f := 0;
        ELSIF x =- 18187 THEN
            exp_f := 0;
        ELSIF x =- 18186 THEN
            exp_f := 0;
        ELSIF x =- 18185 THEN
            exp_f := 0;
        ELSIF x =- 18184 THEN
            exp_f := 0;
        ELSIF x =- 18183 THEN
            exp_f := 0;
        ELSIF x =- 18182 THEN
            exp_f := 0;
        ELSIF x =- 18181 THEN
            exp_f := 0;
        ELSIF x =- 18180 THEN
            exp_f := 0;
        ELSIF x =- 18179 THEN
            exp_f := 0;
        ELSIF x =- 18178 THEN
            exp_f := 0;
        ELSIF x =- 18177 THEN
            exp_f := 0;
        ELSIF x =- 18176 THEN
            exp_f := 0;
        ELSIF x =- 18175 THEN
            exp_f := 0;
        ELSIF x =- 18174 THEN
            exp_f := 0;
        ELSIF x =- 18173 THEN
            exp_f := 0;
        ELSIF x =- 18172 THEN
            exp_f := 0;
        ELSIF x =- 18171 THEN
            exp_f := 0;
        ELSIF x =- 18170 THEN
            exp_f := 0;
        ELSIF x =- 18169 THEN
            exp_f := 0;
        ELSIF x =- 18168 THEN
            exp_f := 0;
        ELSIF x =- 18167 THEN
            exp_f := 0;
        ELSIF x =- 18166 THEN
            exp_f := 0;
        ELSIF x =- 18165 THEN
            exp_f := 0;
        ELSIF x =- 18164 THEN
            exp_f := 0;
        ELSIF x =- 18163 THEN
            exp_f := 0;
        ELSIF x =- 18162 THEN
            exp_f := 0;
        ELSIF x =- 18161 THEN
            exp_f := 0;
        ELSIF x =- 18160 THEN
            exp_f := 0;
        ELSIF x =- 18159 THEN
            exp_f := 0;
        ELSIF x =- 18158 THEN
            exp_f := 0;
        ELSIF x =- 18157 THEN
            exp_f := 0;
        ELSIF x =- 18156 THEN
            exp_f := 0;
        ELSIF x =- 18155 THEN
            exp_f := 0;
        ELSIF x =- 18154 THEN
            exp_f := 0;
        ELSIF x =- 18153 THEN
            exp_f := 0;
        ELSIF x =- 18152 THEN
            exp_f := 0;
        ELSIF x =- 18151 THEN
            exp_f := 0;
        ELSIF x =- 18150 THEN
            exp_f := 0;
        ELSIF x =- 18149 THEN
            exp_f := 0;
        ELSIF x =- 18148 THEN
            exp_f := 0;
        ELSIF x =- 18147 THEN
            exp_f := 0;
        ELSIF x =- 18146 THEN
            exp_f := 0;
        ELSIF x =- 18145 THEN
            exp_f := 0;
        ELSIF x =- 18144 THEN
            exp_f := 0;
        ELSIF x =- 18143 THEN
            exp_f := 0;
        ELSIF x =- 18142 THEN
            exp_f := 0;
        ELSIF x =- 18141 THEN
            exp_f := 0;
        ELSIF x =- 18140 THEN
            exp_f := 0;
        ELSIF x =- 18139 THEN
            exp_f := 0;
        ELSIF x =- 18138 THEN
            exp_f := 0;
        ELSIF x =- 18137 THEN
            exp_f := 0;
        ELSIF x =- 18136 THEN
            exp_f := 0;
        ELSIF x =- 18135 THEN
            exp_f := 0;
        ELSIF x =- 18134 THEN
            exp_f := 0;
        ELSIF x =- 18133 THEN
            exp_f := 0;
        ELSIF x =- 18132 THEN
            exp_f := 0;
        ELSIF x =- 18131 THEN
            exp_f := 0;
        ELSIF x =- 18130 THEN
            exp_f := 0;
        ELSIF x =- 18129 THEN
            exp_f := 0;
        ELSIF x =- 18128 THEN
            exp_f := 0;
        ELSIF x =- 18127 THEN
            exp_f := 0;
        ELSIF x =- 18126 THEN
            exp_f := 0;
        ELSIF x =- 18125 THEN
            exp_f := 0;
        ELSIF x =- 18124 THEN
            exp_f := 0;
        ELSIF x =- 18123 THEN
            exp_f := 0;
        ELSIF x =- 18122 THEN
            exp_f := 0;
        ELSIF x =- 18121 THEN
            exp_f := 0;
        ELSIF x =- 18120 THEN
            exp_f := 0;
        ELSIF x =- 18119 THEN
            exp_f := 0;
        ELSIF x =- 18118 THEN
            exp_f := 0;
        ELSIF x =- 18117 THEN
            exp_f := 0;
        ELSIF x =- 18116 THEN
            exp_f := 0;
        ELSIF x =- 18115 THEN
            exp_f := 0;
        ELSIF x =- 18114 THEN
            exp_f := 0;
        ELSIF x =- 18113 THEN
            exp_f := 0;
        ELSIF x =- 18112 THEN
            exp_f := 0;
        ELSIF x =- 18111 THEN
            exp_f := 0;
        ELSIF x =- 18110 THEN
            exp_f := 0;
        ELSIF x =- 18109 THEN
            exp_f := 0;
        ELSIF x =- 18108 THEN
            exp_f := 0;
        ELSIF x =- 18107 THEN
            exp_f := 0;
        ELSIF x =- 18106 THEN
            exp_f := 0;
        ELSIF x =- 18105 THEN
            exp_f := 0;
        ELSIF x =- 18104 THEN
            exp_f := 0;
        ELSIF x =- 18103 THEN
            exp_f := 0;
        ELSIF x =- 18102 THEN
            exp_f := 0;
        ELSIF x =- 18101 THEN
            exp_f := 0;
        ELSIF x =- 18100 THEN
            exp_f := 0;
        ELSIF x =- 18099 THEN
            exp_f := 0;
        ELSIF x =- 18098 THEN
            exp_f := 0;
        ELSIF x =- 18097 THEN
            exp_f := 0;
        ELSIF x =- 18096 THEN
            exp_f := 0;
        ELSIF x =- 18095 THEN
            exp_f := 0;
        ELSIF x =- 18094 THEN
            exp_f := 0;
        ELSIF x =- 18093 THEN
            exp_f := 0;
        ELSIF x =- 18092 THEN
            exp_f := 0;
        ELSIF x =- 18091 THEN
            exp_f := 0;
        ELSIF x =- 18090 THEN
            exp_f := 0;
        ELSIF x =- 18089 THEN
            exp_f := 0;
        ELSIF x =- 18088 THEN
            exp_f := 0;
        ELSIF x =- 18087 THEN
            exp_f := 0;
        ELSIF x =- 18086 THEN
            exp_f := 0;
        ELSIF x =- 18085 THEN
            exp_f := 0;
        ELSIF x =- 18084 THEN
            exp_f := 0;
        ELSIF x =- 18083 THEN
            exp_f := 0;
        ELSIF x =- 18082 THEN
            exp_f := 0;
        ELSIF x =- 18081 THEN
            exp_f := 0;
        ELSIF x =- 18080 THEN
            exp_f := 0;
        ELSIF x =- 18079 THEN
            exp_f := 0;
        ELSIF x =- 18078 THEN
            exp_f := 0;
        ELSIF x =- 18077 THEN
            exp_f := 0;
        ELSIF x =- 18076 THEN
            exp_f := 0;
        ELSIF x =- 18075 THEN
            exp_f := 0;
        ELSIF x =- 18074 THEN
            exp_f := 0;
        ELSIF x =- 18073 THEN
            exp_f := 0;
        ELSIF x =- 18072 THEN
            exp_f := 0;
        ELSIF x =- 18071 THEN
            exp_f := 0;
        ELSIF x =- 18070 THEN
            exp_f := 0;
        ELSIF x =- 18069 THEN
            exp_f := 0;
        ELSIF x =- 18068 THEN
            exp_f := 0;
        ELSIF x =- 18067 THEN
            exp_f := 0;
        ELSIF x =- 18066 THEN
            exp_f := 0;
        ELSIF x =- 18065 THEN
            exp_f := 0;
        ELSIF x =- 18064 THEN
            exp_f := 0;
        ELSIF x =- 18063 THEN
            exp_f := 0;
        ELSIF x =- 18062 THEN
            exp_f := 0;
        ELSIF x =- 18061 THEN
            exp_f := 0;
        ELSIF x =- 18060 THEN
            exp_f := 0;
        ELSIF x =- 18059 THEN
            exp_f := 0;
        ELSIF x =- 18058 THEN
            exp_f := 0;
        ELSIF x =- 18057 THEN
            exp_f := 0;
        ELSIF x =- 18056 THEN
            exp_f := 0;
        ELSIF x =- 18055 THEN
            exp_f := 0;
        ELSIF x =- 18054 THEN
            exp_f := 0;
        ELSIF x =- 18053 THEN
            exp_f := 0;
        ELSIF x =- 18052 THEN
            exp_f := 0;
        ELSIF x =- 18051 THEN
            exp_f := 0;
        ELSIF x =- 18050 THEN
            exp_f := 0;
        ELSIF x =- 18049 THEN
            exp_f := 0;
        ELSIF x =- 18048 THEN
            exp_f := 0;
        ELSIF x =- 18047 THEN
            exp_f := 0;
        ELSIF x =- 18046 THEN
            exp_f := 0;
        ELSIF x =- 18045 THEN
            exp_f := 0;
        ELSIF x =- 18044 THEN
            exp_f := 0;
        ELSIF x =- 18043 THEN
            exp_f := 0;
        ELSIF x =- 18042 THEN
            exp_f := 0;
        ELSIF x =- 18041 THEN
            exp_f := 0;
        ELSIF x =- 18040 THEN
            exp_f := 0;
        ELSIF x =- 18039 THEN
            exp_f := 0;
        ELSIF x =- 18038 THEN
            exp_f := 0;
        ELSIF x =- 18037 THEN
            exp_f := 0;
        ELSIF x =- 18036 THEN
            exp_f := 0;
        ELSIF x =- 18035 THEN
            exp_f := 0;
        ELSIF x =- 18034 THEN
            exp_f := 0;
        ELSIF x =- 18033 THEN
            exp_f := 0;
        ELSIF x =- 18032 THEN
            exp_f := 0;
        ELSIF x =- 18031 THEN
            exp_f := 0;
        ELSIF x =- 18030 THEN
            exp_f := 0;
        ELSIF x =- 18029 THEN
            exp_f := 0;
        ELSIF x =- 18028 THEN
            exp_f := 0;
        ELSIF x =- 18027 THEN
            exp_f := 0;
        ELSIF x =- 18026 THEN
            exp_f := 0;
        ELSIF x =- 18025 THEN
            exp_f := 0;
        ELSIF x =- 18024 THEN
            exp_f := 0;
        ELSIF x =- 18023 THEN
            exp_f := 0;
        ELSIF x =- 18022 THEN
            exp_f := 0;
        ELSIF x =- 18021 THEN
            exp_f := 0;
        ELSIF x =- 18020 THEN
            exp_f := 0;
        ELSIF x =- 18019 THEN
            exp_f := 0;
        ELSIF x =- 18018 THEN
            exp_f := 0;
        ELSIF x =- 18017 THEN
            exp_f := 0;
        ELSIF x =- 18016 THEN
            exp_f := 0;
        ELSIF x =- 18015 THEN
            exp_f := 0;
        ELSIF x =- 18014 THEN
            exp_f := 0;
        ELSIF x =- 18013 THEN
            exp_f := 0;
        ELSIF x =- 18012 THEN
            exp_f := 0;
        ELSIF x =- 18011 THEN
            exp_f := 0;
        ELSIF x =- 18010 THEN
            exp_f := 0;
        ELSIF x =- 18009 THEN
            exp_f := 0;
        ELSIF x =- 18008 THEN
            exp_f := 0;
        ELSIF x =- 18007 THEN
            exp_f := 0;
        ELSIF x =- 18006 THEN
            exp_f := 0;
        ELSIF x =- 18005 THEN
            exp_f := 0;
        ELSIF x =- 18004 THEN
            exp_f := 0;
        ELSIF x =- 18003 THEN
            exp_f := 0;
        ELSIF x =- 18002 THEN
            exp_f := 0;
        ELSIF x =- 18001 THEN
            exp_f := 0;
        ELSIF x =- 18000 THEN
            exp_f := 0;
        ELSIF x =- 17999 THEN
            exp_f := 0;
        ELSIF x =- 17998 THEN
            exp_f := 0;
        ELSIF x =- 17997 THEN
            exp_f := 0;
        ELSIF x =- 17996 THEN
            exp_f := 0;
        ELSIF x =- 17995 THEN
            exp_f := 0;
        ELSIF x =- 17994 THEN
            exp_f := 0;
        ELSIF x =- 17993 THEN
            exp_f := 0;
        ELSIF x =- 17992 THEN
            exp_f := 0;
        ELSIF x =- 17991 THEN
            exp_f := 0;
        ELSIF x =- 17990 THEN
            exp_f := 0;
        ELSIF x =- 17989 THEN
            exp_f := 0;
        ELSIF x =- 17988 THEN
            exp_f := 0;
        ELSIF x =- 17987 THEN
            exp_f := 0;
        ELSIF x =- 17986 THEN
            exp_f := 0;
        ELSIF x =- 17985 THEN
            exp_f := 0;
        ELSIF x =- 17984 THEN
            exp_f := 0;
        ELSIF x =- 17983 THEN
            exp_f := 0;
        ELSIF x =- 17982 THEN
            exp_f := 0;
        ELSIF x =- 17981 THEN
            exp_f := 0;
        ELSIF x =- 17980 THEN
            exp_f := 0;
        ELSIF x =- 17979 THEN
            exp_f := 0;
        ELSIF x =- 17978 THEN
            exp_f := 0;
        ELSIF x =- 17977 THEN
            exp_f := 0;
        ELSIF x =- 17976 THEN
            exp_f := 0;
        ELSIF x =- 17975 THEN
            exp_f := 0;
        ELSIF x =- 17974 THEN
            exp_f := 0;
        ELSIF x =- 17973 THEN
            exp_f := 0;
        ELSIF x =- 17972 THEN
            exp_f := 0;
        ELSIF x =- 17971 THEN
            exp_f := 0;
        ELSIF x =- 17970 THEN
            exp_f := 0;
        ELSIF x =- 17969 THEN
            exp_f := 0;
        ELSIF x =- 17968 THEN
            exp_f := 0;
        ELSIF x =- 17967 THEN
            exp_f := 0;
        ELSIF x =- 17966 THEN
            exp_f := 0;
        ELSIF x =- 17965 THEN
            exp_f := 0;
        ELSIF x =- 17964 THEN
            exp_f := 0;
        ELSIF x =- 17963 THEN
            exp_f := 0;
        ELSIF x =- 17962 THEN
            exp_f := 0;
        ELSIF x =- 17961 THEN
            exp_f := 0;
        ELSIF x =- 17960 THEN
            exp_f := 0;
        ELSIF x =- 17959 THEN
            exp_f := 0;
        ELSIF x =- 17958 THEN
            exp_f := 0;
        ELSIF x =- 17957 THEN
            exp_f := 0;
        ELSIF x =- 17956 THEN
            exp_f := 0;
        ELSIF x =- 17955 THEN
            exp_f := 0;
        ELSIF x =- 17954 THEN
            exp_f := 0;
        ELSIF x =- 17953 THEN
            exp_f := 0;
        ELSIF x =- 17952 THEN
            exp_f := 0;
        ELSIF x =- 17951 THEN
            exp_f := 0;
        ELSIF x =- 17950 THEN
            exp_f := 0;
        ELSIF x =- 17949 THEN
            exp_f := 0;
        ELSIF x =- 17948 THEN
            exp_f := 0;
        ELSIF x =- 17947 THEN
            exp_f := 0;
        ELSIF x =- 17946 THEN
            exp_f := 0;
        ELSIF x =- 17945 THEN
            exp_f := 0;
        ELSIF x =- 17944 THEN
            exp_f := 0;
        ELSIF x =- 17943 THEN
            exp_f := 0;
        ELSIF x =- 17942 THEN
            exp_f := 0;
        ELSIF x =- 17941 THEN
            exp_f := 0;
        ELSIF x =- 17940 THEN
            exp_f := 0;
        ELSIF x =- 17939 THEN
            exp_f := 0;
        ELSIF x =- 17938 THEN
            exp_f := 0;
        ELSIF x =- 17937 THEN
            exp_f := 0;
        ELSIF x =- 17936 THEN
            exp_f := 0;
        ELSIF x =- 17935 THEN
            exp_f := 0;
        ELSIF x =- 17934 THEN
            exp_f := 0;
        ELSIF x =- 17933 THEN
            exp_f := 0;
        ELSIF x =- 17932 THEN
            exp_f := 0;
        ELSIF x =- 17931 THEN
            exp_f := 0;
        ELSIF x =- 17930 THEN
            exp_f := 0;
        ELSIF x =- 17929 THEN
            exp_f := 0;
        ELSIF x =- 17928 THEN
            exp_f := 0;
        ELSIF x =- 17927 THEN
            exp_f := 0;
        ELSIF x =- 17926 THEN
            exp_f := 0;
        ELSIF x =- 17925 THEN
            exp_f := 0;
        ELSIF x =- 17924 THEN
            exp_f := 0;
        ELSIF x =- 17923 THEN
            exp_f := 0;
        ELSIF x =- 17922 THEN
            exp_f := 0;
        ELSIF x =- 17921 THEN
            exp_f := 0;
        ELSIF x =- 17920 THEN
            exp_f := 0;
        ELSIF x =- 17919 THEN
            exp_f := 0;
        ELSIF x =- 17918 THEN
            exp_f := 0;
        ELSIF x =- 17917 THEN
            exp_f := 0;
        ELSIF x =- 17916 THEN
            exp_f := 0;
        ELSIF x =- 17915 THEN
            exp_f := 0;
        ELSIF x =- 17914 THEN
            exp_f := 0;
        ELSIF x =- 17913 THEN
            exp_f := 0;
        ELSIF x =- 17912 THEN
            exp_f := 0;
        ELSIF x =- 17911 THEN
            exp_f := 0;
        ELSIF x =- 17910 THEN
            exp_f := 0;
        ELSIF x =- 17909 THEN
            exp_f := 0;
        ELSIF x =- 17908 THEN
            exp_f := 0;
        ELSIF x =- 17907 THEN
            exp_f := 0;
        ELSIF x =- 17906 THEN
            exp_f := 0;
        ELSIF x =- 17905 THEN
            exp_f := 0;
        ELSIF x =- 17904 THEN
            exp_f := 0;
        ELSIF x =- 17903 THEN
            exp_f := 0;
        ELSIF x =- 17902 THEN
            exp_f := 0;
        ELSIF x =- 17901 THEN
            exp_f := 0;
        ELSIF x =- 17900 THEN
            exp_f := 0;
        ELSIF x =- 17899 THEN
            exp_f := 0;
        ELSIF x =- 17898 THEN
            exp_f := 0;
        ELSIF x =- 17897 THEN
            exp_f := 0;
        ELSIF x =- 17896 THEN
            exp_f := 0;
        ELSIF x =- 17895 THEN
            exp_f := 0;
        ELSIF x =- 17894 THEN
            exp_f := 0;
        ELSIF x =- 17893 THEN
            exp_f := 0;
        ELSIF x =- 17892 THEN
            exp_f := 0;
        ELSIF x =- 17891 THEN
            exp_f := 0;
        ELSIF x =- 17890 THEN
            exp_f := 0;
        ELSIF x =- 17889 THEN
            exp_f := 0;
        ELSIF x =- 17888 THEN
            exp_f := 0;
        ELSIF x =- 17887 THEN
            exp_f := 0;
        ELSIF x =- 17886 THEN
            exp_f := 0;
        ELSIF x =- 17885 THEN
            exp_f := 0;
        ELSIF x =- 17884 THEN
            exp_f := 0;
        ELSIF x =- 17883 THEN
            exp_f := 0;
        ELSIF x =- 17882 THEN
            exp_f := 0;
        ELSIF x =- 17881 THEN
            exp_f := 0;
        ELSIF x =- 17880 THEN
            exp_f := 0;
        ELSIF x =- 17879 THEN
            exp_f := 0;
        ELSIF x =- 17878 THEN
            exp_f := 0;
        ELSIF x =- 17877 THEN
            exp_f := 0;
        ELSIF x =- 17876 THEN
            exp_f := 0;
        ELSIF x =- 17875 THEN
            exp_f := 0;
        ELSIF x =- 17874 THEN
            exp_f := 0;
        ELSIF x =- 17873 THEN
            exp_f := 0;
        ELSIF x =- 17872 THEN
            exp_f := 0;
        ELSIF x =- 17871 THEN
            exp_f := 0;
        ELSIF x =- 17870 THEN
            exp_f := 0;
        ELSIF x =- 17869 THEN
            exp_f := 0;
        ELSIF x =- 17868 THEN
            exp_f := 0;
        ELSIF x =- 17867 THEN
            exp_f := 0;
        ELSIF x =- 17866 THEN
            exp_f := 0;
        ELSIF x =- 17865 THEN
            exp_f := 0;
        ELSIF x =- 17864 THEN
            exp_f := 0;
        ELSIF x =- 17863 THEN
            exp_f := 0;
        ELSIF x =- 17862 THEN
            exp_f := 0;
        ELSIF x =- 17861 THEN
            exp_f := 0;
        ELSIF x =- 17860 THEN
            exp_f := 0;
        ELSIF x =- 17859 THEN
            exp_f := 0;
        ELSIF x =- 17858 THEN
            exp_f := 0;
        ELSIF x =- 17857 THEN
            exp_f := 0;
        ELSIF x =- 17856 THEN
            exp_f := 0;
        ELSIF x =- 17855 THEN
            exp_f := 0;
        ELSIF x =- 17854 THEN
            exp_f := 0;
        ELSIF x =- 17853 THEN
            exp_f := 0;
        ELSIF x =- 17852 THEN
            exp_f := 0;
        ELSIF x =- 17851 THEN
            exp_f := 0;
        ELSIF x =- 17850 THEN
            exp_f := 0;
        ELSIF x =- 17849 THEN
            exp_f := 0;
        ELSIF x =- 17848 THEN
            exp_f := 0;
        ELSIF x =- 17847 THEN
            exp_f := 0;
        ELSIF x =- 17846 THEN
            exp_f := 0;
        ELSIF x =- 17845 THEN
            exp_f := 0;
        ELSIF x =- 17844 THEN
            exp_f := 0;
        ELSIF x =- 17843 THEN
            exp_f := 0;
        ELSIF x =- 17842 THEN
            exp_f := 0;
        ELSIF x =- 17841 THEN
            exp_f := 0;
        ELSIF x =- 17840 THEN
            exp_f := 0;
        ELSIF x =- 17839 THEN
            exp_f := 0;
        ELSIF x =- 17838 THEN
            exp_f := 0;
        ELSIF x =- 17837 THEN
            exp_f := 0;
        ELSIF x =- 17836 THEN
            exp_f := 0;
        ELSIF x =- 17835 THEN
            exp_f := 0;
        ELSIF x =- 17834 THEN
            exp_f := 0;
        ELSIF x =- 17833 THEN
            exp_f := 0;
        ELSIF x =- 17832 THEN
            exp_f := 0;
        ELSIF x =- 17831 THEN
            exp_f := 0;
        ELSIF x =- 17830 THEN
            exp_f := 0;
        ELSIF x =- 17829 THEN
            exp_f := 0;
        ELSIF x =- 17828 THEN
            exp_f := 0;
        ELSIF x =- 17827 THEN
            exp_f := 0;
        ELSIF x =- 17826 THEN
            exp_f := 0;
        ELSIF x =- 17825 THEN
            exp_f := 0;
        ELSIF x =- 17824 THEN
            exp_f := 0;
        ELSIF x =- 17823 THEN
            exp_f := 0;
        ELSIF x =- 17822 THEN
            exp_f := 0;
        ELSIF x =- 17821 THEN
            exp_f := 0;
        ELSIF x =- 17820 THEN
            exp_f := 0;
        ELSIF x =- 17819 THEN
            exp_f := 0;
        ELSIF x =- 17818 THEN
            exp_f := 0;
        ELSIF x =- 17817 THEN
            exp_f := 0;
        ELSIF x =- 17816 THEN
            exp_f := 0;
        ELSIF x =- 17815 THEN
            exp_f := 0;
        ELSIF x =- 17814 THEN
            exp_f := 0;
        ELSIF x =- 17813 THEN
            exp_f := 0;
        ELSIF x =- 17812 THEN
            exp_f := 0;
        ELSIF x =- 17811 THEN
            exp_f := 0;
        ELSIF x =- 17810 THEN
            exp_f := 0;
        ELSIF x =- 17809 THEN
            exp_f := 0;
        ELSIF x =- 17808 THEN
            exp_f := 0;
        ELSIF x =- 17807 THEN
            exp_f := 0;
        ELSIF x =- 17806 THEN
            exp_f := 0;
        ELSIF x =- 17805 THEN
            exp_f := 0;
        ELSIF x =- 17804 THEN
            exp_f := 0;
        ELSIF x =- 17803 THEN
            exp_f := 0;
        ELSIF x =- 17802 THEN
            exp_f := 0;
        ELSIF x =- 17801 THEN
            exp_f := 0;
        ELSIF x =- 17800 THEN
            exp_f := 0;
        ELSIF x =- 17799 THEN
            exp_f := 0;
        ELSIF x =- 17798 THEN
            exp_f := 0;
        ELSIF x =- 17797 THEN
            exp_f := 0;
        ELSIF x =- 17796 THEN
            exp_f := 0;
        ELSIF x =- 17795 THEN
            exp_f := 0;
        ELSIF x =- 17794 THEN
            exp_f := 0;
        ELSIF x =- 17793 THEN
            exp_f := 0;
        ELSIF x =- 17792 THEN
            exp_f := 0;
        ELSIF x =- 17791 THEN
            exp_f := 0;
        ELSIF x =- 17790 THEN
            exp_f := 0;
        ELSIF x =- 17789 THEN
            exp_f := 0;
        ELSIF x =- 17788 THEN
            exp_f := 0;
        ELSIF x =- 17787 THEN
            exp_f := 0;
        ELSIF x =- 17786 THEN
            exp_f := 0;
        ELSIF x =- 17785 THEN
            exp_f := 0;
        ELSIF x =- 17784 THEN
            exp_f := 0;
        ELSIF x =- 17783 THEN
            exp_f := 0;
        ELSIF x =- 17782 THEN
            exp_f := 0;
        ELSIF x =- 17781 THEN
            exp_f := 0;
        ELSIF x =- 17780 THEN
            exp_f := 0;
        ELSIF x =- 17779 THEN
            exp_f := 0;
        ELSIF x =- 17778 THEN
            exp_f := 0;
        ELSIF x =- 17777 THEN
            exp_f := 0;
        ELSIF x =- 17776 THEN
            exp_f := 0;
        ELSIF x =- 17775 THEN
            exp_f := 0;
        ELSIF x =- 17774 THEN
            exp_f := 0;
        ELSIF x =- 17773 THEN
            exp_f := 0;
        ELSIF x =- 17772 THEN
            exp_f := 0;
        ELSIF x =- 17771 THEN
            exp_f := 0;
        ELSIF x =- 17770 THEN
            exp_f := 0;
        ELSIF x =- 17769 THEN
            exp_f := 0;
        ELSIF x =- 17768 THEN
            exp_f := 0;
        ELSIF x =- 17767 THEN
            exp_f := 0;
        ELSIF x =- 17766 THEN
            exp_f := 0;
        ELSIF x =- 17765 THEN
            exp_f := 0;
        ELSIF x =- 17764 THEN
            exp_f := 0;
        ELSIF x =- 17763 THEN
            exp_f := 0;
        ELSIF x =- 17762 THEN
            exp_f := 0;
        ELSIF x =- 17761 THEN
            exp_f := 0;
        ELSIF x =- 17760 THEN
            exp_f := 0;
        ELSIF x =- 17759 THEN
            exp_f := 0;
        ELSIF x =- 17758 THEN
            exp_f := 0;
        ELSIF x =- 17757 THEN
            exp_f := 0;
        ELSIF x =- 17756 THEN
            exp_f := 0;
        ELSIF x =- 17755 THEN
            exp_f := 0;
        ELSIF x =- 17754 THEN
            exp_f := 0;
        ELSIF x =- 17753 THEN
            exp_f := 0;
        ELSIF x =- 17752 THEN
            exp_f := 0;
        ELSIF x =- 17751 THEN
            exp_f := 0;
        ELSIF x =- 17750 THEN
            exp_f := 0;
        ELSIF x =- 17749 THEN
            exp_f := 0;
        ELSIF x =- 17748 THEN
            exp_f := 0;
        ELSIF x =- 17747 THEN
            exp_f := 0;
        ELSIF x =- 17746 THEN
            exp_f := 0;
        ELSIF x =- 17745 THEN
            exp_f := 0;
        ELSIF x =- 17744 THEN
            exp_f := 0;
        ELSIF x =- 17743 THEN
            exp_f := 0;
        ELSIF x =- 17742 THEN
            exp_f := 0;
        ELSIF x =- 17741 THEN
            exp_f := 0;
        ELSIF x =- 17740 THEN
            exp_f := 0;
        ELSIF x =- 17739 THEN
            exp_f := 0;
        ELSIF x =- 17738 THEN
            exp_f := 0;
        ELSIF x =- 17737 THEN
            exp_f := 0;
        ELSIF x =- 17736 THEN
            exp_f := 0;
        ELSIF x =- 17735 THEN
            exp_f := 0;
        ELSIF x =- 17734 THEN
            exp_f := 0;
        ELSIF x =- 17733 THEN
            exp_f := 0;
        ELSIF x =- 17732 THEN
            exp_f := 0;
        ELSIF x =- 17731 THEN
            exp_f := 0;
        ELSIF x =- 17730 THEN
            exp_f := 0;
        ELSIF x =- 17729 THEN
            exp_f := 0;
        ELSIF x =- 17728 THEN
            exp_f := 0;
        ELSIF x =- 17727 THEN
            exp_f := 0;
        ELSIF x =- 17726 THEN
            exp_f := 0;
        ELSIF x =- 17725 THEN
            exp_f := 0;
        ELSIF x =- 17724 THEN
            exp_f := 0;
        ELSIF x =- 17723 THEN
            exp_f := 0;
        ELSIF x =- 17722 THEN
            exp_f := 0;
        ELSIF x =- 17721 THEN
            exp_f := 0;
        ELSIF x =- 17720 THEN
            exp_f := 0;
        ELSIF x =- 17719 THEN
            exp_f := 0;
        ELSIF x =- 17718 THEN
            exp_f := 0;
        ELSIF x =- 17717 THEN
            exp_f := 0;
        ELSIF x =- 17716 THEN
            exp_f := 0;
        ELSIF x =- 17715 THEN
            exp_f := 0;
        ELSIF x =- 17714 THEN
            exp_f := 0;
        ELSIF x =- 17713 THEN
            exp_f := 0;
        ELSIF x =- 17712 THEN
            exp_f := 0;
        ELSIF x =- 17711 THEN
            exp_f := 0;
        ELSIF x =- 17710 THEN
            exp_f := 0;
        ELSIF x =- 17709 THEN
            exp_f := 0;
        ELSIF x =- 17708 THEN
            exp_f := 0;
        ELSIF x =- 17707 THEN
            exp_f := 0;
        ELSIF x =- 17706 THEN
            exp_f := 0;
        ELSIF x =- 17705 THEN
            exp_f := 0;
        ELSIF x =- 17704 THEN
            exp_f := 0;
        ELSIF x =- 17703 THEN
            exp_f := 0;
        ELSIF x =- 17702 THEN
            exp_f := 0;
        ELSIF x =- 17701 THEN
            exp_f := 0;
        ELSIF x =- 17700 THEN
            exp_f := 0;
        ELSIF x =- 17699 THEN
            exp_f := 0;
        ELSIF x =- 17698 THEN
            exp_f := 0;
        ELSIF x =- 17697 THEN
            exp_f := 0;
        ELSIF x =- 17696 THEN
            exp_f := 0;
        ELSIF x =- 17695 THEN
            exp_f := 0;
        ELSIF x =- 17694 THEN
            exp_f := 0;
        ELSIF x =- 17693 THEN
            exp_f := 0;
        ELSIF x =- 17692 THEN
            exp_f := 0;
        ELSIF x =- 17691 THEN
            exp_f := 0;
        ELSIF x =- 17690 THEN
            exp_f := 0;
        ELSIF x =- 17689 THEN
            exp_f := 0;
        ELSIF x =- 17688 THEN
            exp_f := 0;
        ELSIF x =- 17687 THEN
            exp_f := 0;
        ELSIF x =- 17686 THEN
            exp_f := 0;
        ELSIF x =- 17685 THEN
            exp_f := 0;
        ELSIF x =- 17684 THEN
            exp_f := 0;
        ELSIF x =- 17683 THEN
            exp_f := 0;
        ELSIF x =- 17682 THEN
            exp_f := 0;
        ELSIF x =- 17681 THEN
            exp_f := 0;
        ELSIF x =- 17680 THEN
            exp_f := 0;
        ELSIF x =- 17679 THEN
            exp_f := 0;
        ELSIF x =- 17678 THEN
            exp_f := 0;
        ELSIF x =- 17677 THEN
            exp_f := 0;
        ELSIF x =- 17676 THEN
            exp_f := 0;
        ELSIF x =- 17675 THEN
            exp_f := 0;
        ELSIF x =- 17674 THEN
            exp_f := 0;
        ELSIF x =- 17673 THEN
            exp_f := 0;
        ELSIF x =- 17672 THEN
            exp_f := 0;
        ELSIF x =- 17671 THEN
            exp_f := 0;
        ELSIF x =- 17670 THEN
            exp_f := 0;
        ELSIF x =- 17669 THEN
            exp_f := 0;
        ELSIF x =- 17668 THEN
            exp_f := 0;
        ELSIF x =- 17667 THEN
            exp_f := 0;
        ELSIF x =- 17666 THEN
            exp_f := 0;
        ELSIF x =- 17665 THEN
            exp_f := 0;
        ELSIF x =- 17664 THEN
            exp_f := 0;
        ELSIF x =- 17663 THEN
            exp_f := 0;
        ELSIF x =- 17662 THEN
            exp_f := 0;
        ELSIF x =- 17661 THEN
            exp_f := 0;
        ELSIF x =- 17660 THEN
            exp_f := 0;
        ELSIF x =- 17659 THEN
            exp_f := 0;
        ELSIF x =- 17658 THEN
            exp_f := 0;
        ELSIF x =- 17657 THEN
            exp_f := 0;
        ELSIF x =- 17656 THEN
            exp_f := 0;
        ELSIF x =- 17655 THEN
            exp_f := 0;
        ELSIF x =- 17654 THEN
            exp_f := 0;
        ELSIF x =- 17653 THEN
            exp_f := 0;
        ELSIF x =- 17652 THEN
            exp_f := 0;
        ELSIF x =- 17651 THEN
            exp_f := 0;
        ELSIF x =- 17650 THEN
            exp_f := 0;
        ELSIF x =- 17649 THEN
            exp_f := 0;
        ELSIF x =- 17648 THEN
            exp_f := 0;
        ELSIF x =- 17647 THEN
            exp_f := 0;
        ELSIF x =- 17646 THEN
            exp_f := 0;
        ELSIF x =- 17645 THEN
            exp_f := 0;
        ELSIF x =- 17644 THEN
            exp_f := 0;
        ELSIF x =- 17643 THEN
            exp_f := 0;
        ELSIF x =- 17642 THEN
            exp_f := 0;
        ELSIF x =- 17641 THEN
            exp_f := 0;
        ELSIF x =- 17640 THEN
            exp_f := 0;
        ELSIF x =- 17639 THEN
            exp_f := 0;
        ELSIF x =- 17638 THEN
            exp_f := 0;
        ELSIF x =- 17637 THEN
            exp_f := 0;
        ELSIF x =- 17636 THEN
            exp_f := 0;
        ELSIF x =- 17635 THEN
            exp_f := 0;
        ELSIF x =- 17634 THEN
            exp_f := 0;
        ELSIF x =- 17633 THEN
            exp_f := 0;
        ELSIF x =- 17632 THEN
            exp_f := 0;
        ELSIF x =- 17631 THEN
            exp_f := 0;
        ELSIF x =- 17630 THEN
            exp_f := 0;
        ELSIF x =- 17629 THEN
            exp_f := 0;
        ELSIF x =- 17628 THEN
            exp_f := 0;
        ELSIF x =- 17627 THEN
            exp_f := 0;
        ELSIF x =- 17626 THEN
            exp_f := 0;
        ELSIF x =- 17625 THEN
            exp_f := 0;
        ELSIF x =- 17624 THEN
            exp_f := 0;
        ELSIF x =- 17623 THEN
            exp_f := 0;
        ELSIF x =- 17622 THEN
            exp_f := 0;
        ELSIF x =- 17621 THEN
            exp_f := 0;
        ELSIF x =- 17620 THEN
            exp_f := 0;
        ELSIF x =- 17619 THEN
            exp_f := 0;
        ELSIF x =- 17618 THEN
            exp_f := 0;
        ELSIF x =- 17617 THEN
            exp_f := 0;
        ELSIF x =- 17616 THEN
            exp_f := 0;
        ELSIF x =- 17615 THEN
            exp_f := 0;
        ELSIF x =- 17614 THEN
            exp_f := 0;
        ELSIF x =- 17613 THEN
            exp_f := 0;
        ELSIF x =- 17612 THEN
            exp_f := 0;
        ELSIF x =- 17611 THEN
            exp_f := 0;
        ELSIF x =- 17610 THEN
            exp_f := 0;
        ELSIF x =- 17609 THEN
            exp_f := 0;
        ELSIF x =- 17608 THEN
            exp_f := 0;
        ELSIF x =- 17607 THEN
            exp_f := 0;
        ELSIF x =- 17606 THEN
            exp_f := 0;
        ELSIF x =- 17605 THEN
            exp_f := 0;
        ELSIF x =- 17604 THEN
            exp_f := 0;
        ELSIF x =- 17603 THEN
            exp_f := 0;
        ELSIF x =- 17602 THEN
            exp_f := 0;
        ELSIF x =- 17601 THEN
            exp_f := 0;
        ELSIF x =- 17600 THEN
            exp_f := 0;
        ELSIF x =- 17599 THEN
            exp_f := 0;
        ELSIF x =- 17598 THEN
            exp_f := 0;
        ELSIF x =- 17597 THEN
            exp_f := 0;
        ELSIF x =- 17596 THEN
            exp_f := 0;
        ELSIF x =- 17595 THEN
            exp_f := 0;
        ELSIF x =- 17594 THEN
            exp_f := 0;
        ELSIF x =- 17593 THEN
            exp_f := 0;
        ELSIF x =- 17592 THEN
            exp_f := 0;
        ELSIF x =- 17591 THEN
            exp_f := 0;
        ELSIF x =- 17590 THEN
            exp_f := 0;
        ELSIF x =- 17589 THEN
            exp_f := 0;
        ELSIF x =- 17588 THEN
            exp_f := 0;
        ELSIF x =- 17587 THEN
            exp_f := 0;
        ELSIF x =- 17586 THEN
            exp_f := 0;
        ELSIF x =- 17585 THEN
            exp_f := 0;
        ELSIF x =- 17584 THEN
            exp_f := 0;
        ELSIF x =- 17583 THEN
            exp_f := 0;
        ELSIF x =- 17582 THEN
            exp_f := 0;
        ELSIF x =- 17581 THEN
            exp_f := 0;
        ELSIF x =- 17580 THEN
            exp_f := 0;
        ELSIF x =- 17579 THEN
            exp_f := 0;
        ELSIF x =- 17578 THEN
            exp_f := 0;
        ELSIF x =- 17577 THEN
            exp_f := 0;
        ELSIF x =- 17576 THEN
            exp_f := 0;
        ELSIF x =- 17575 THEN
            exp_f := 0;
        ELSIF x =- 17574 THEN
            exp_f := 0;
        ELSIF x =- 17573 THEN
            exp_f := 0;
        ELSIF x =- 17572 THEN
            exp_f := 0;
        ELSIF x =- 17571 THEN
            exp_f := 0;
        ELSIF x =- 17570 THEN
            exp_f := 0;
        ELSIF x =- 17569 THEN
            exp_f := 0;
        ELSIF x =- 17568 THEN
            exp_f := 0;
        ELSIF x =- 17567 THEN
            exp_f := 0;
        ELSIF x =- 17566 THEN
            exp_f := 0;
        ELSIF x =- 17565 THEN
            exp_f := 0;
        ELSIF x =- 17564 THEN
            exp_f := 0;
        ELSIF x =- 17563 THEN
            exp_f := 0;
        ELSIF x =- 17562 THEN
            exp_f := 0;
        ELSIF x =- 17561 THEN
            exp_f := 0;
        ELSIF x =- 17560 THEN
            exp_f := 0;
        ELSIF x =- 17559 THEN
            exp_f := 0;
        ELSIF x =- 17558 THEN
            exp_f := 0;
        ELSIF x =- 17557 THEN
            exp_f := 0;
        ELSIF x =- 17556 THEN
            exp_f := 0;
        ELSIF x =- 17555 THEN
            exp_f := 0;
        ELSIF x =- 17554 THEN
            exp_f := 0;
        ELSIF x =- 17553 THEN
            exp_f := 0;
        ELSIF x =- 17552 THEN
            exp_f := 0;
        ELSIF x =- 17551 THEN
            exp_f := 0;
        ELSIF x =- 17550 THEN
            exp_f := 0;
        ELSIF x =- 17549 THEN
            exp_f := 0;
        ELSIF x =- 17548 THEN
            exp_f := 0;
        ELSIF x =- 17547 THEN
            exp_f := 0;
        ELSIF x =- 17546 THEN
            exp_f := 0;
        ELSIF x =- 17545 THEN
            exp_f := 0;
        ELSIF x =- 17544 THEN
            exp_f := 0;
        ELSIF x =- 17543 THEN
            exp_f := 0;
        ELSIF x =- 17542 THEN
            exp_f := 0;
        ELSIF x =- 17541 THEN
            exp_f := 0;
        ELSIF x =- 17540 THEN
            exp_f := 0;
        ELSIF x =- 17539 THEN
            exp_f := 0;
        ELSIF x =- 17538 THEN
            exp_f := 0;
        ELSIF x =- 17537 THEN
            exp_f := 0;
        ELSIF x =- 17536 THEN
            exp_f := 0;
        ELSIF x =- 17535 THEN
            exp_f := 0;
        ELSIF x =- 17534 THEN
            exp_f := 0;
        ELSIF x =- 17533 THEN
            exp_f := 0;
        ELSIF x =- 17532 THEN
            exp_f := 0;
        ELSIF x =- 17531 THEN
            exp_f := 0;
        ELSIF x =- 17530 THEN
            exp_f := 0;
        ELSIF x =- 17529 THEN
            exp_f := 0;
        ELSIF x =- 17528 THEN
            exp_f := 0;
        ELSIF x =- 17527 THEN
            exp_f := 0;
        ELSIF x =- 17526 THEN
            exp_f := 0;
        ELSIF x =- 17525 THEN
            exp_f := 0;
        ELSIF x =- 17524 THEN
            exp_f := 0;
        ELSIF x =- 17523 THEN
            exp_f := 0;
        ELSIF x =- 17522 THEN
            exp_f := 0;
        ELSIF x =- 17521 THEN
            exp_f := 0;
        ELSIF x =- 17520 THEN
            exp_f := 0;
        ELSIF x =- 17519 THEN
            exp_f := 0;
        ELSIF x =- 17518 THEN
            exp_f := 0;
        ELSIF x =- 17517 THEN
            exp_f := 0;
        ELSIF x =- 17516 THEN
            exp_f := 0;
        ELSIF x =- 17515 THEN
            exp_f := 0;
        ELSIF x =- 17514 THEN
            exp_f := 0;
        ELSIF x =- 17513 THEN
            exp_f := 0;
        ELSIF x =- 17512 THEN
            exp_f := 0;
        ELSIF x =- 17511 THEN
            exp_f := 0;
        ELSIF x =- 17510 THEN
            exp_f := 0;
        ELSIF x =- 17509 THEN
            exp_f := 0;
        ELSIF x =- 17508 THEN
            exp_f := 0;
        ELSIF x =- 17507 THEN
            exp_f := 0;
        ELSIF x =- 17506 THEN
            exp_f := 0;
        ELSIF x =- 17505 THEN
            exp_f := 0;
        ELSIF x =- 17504 THEN
            exp_f := 0;
        ELSIF x =- 17503 THEN
            exp_f := 0;
        ELSIF x =- 17502 THEN
            exp_f := 0;
        ELSIF x =- 17501 THEN
            exp_f := 0;
        ELSIF x =- 17500 THEN
            exp_f := 0;
        ELSIF x =- 17499 THEN
            exp_f := 0;
        ELSIF x =- 17498 THEN
            exp_f := 0;
        ELSIF x =- 17497 THEN
            exp_f := 0;
        ELSIF x =- 17496 THEN
            exp_f := 0;
        ELSIF x =- 17495 THEN
            exp_f := 0;
        ELSIF x =- 17494 THEN
            exp_f := 0;
        ELSIF x =- 17493 THEN
            exp_f := 0;
        ELSIF x =- 17492 THEN
            exp_f := 0;
        ELSIF x =- 17491 THEN
            exp_f := 0;
        ELSIF x =- 17490 THEN
            exp_f := 0;
        ELSIF x =- 17489 THEN
            exp_f := 0;
        ELSIF x =- 17488 THEN
            exp_f := 0;
        ELSIF x =- 17487 THEN
            exp_f := 0;
        ELSIF x =- 17486 THEN
            exp_f := 0;
        ELSIF x =- 17485 THEN
            exp_f := 0;
        ELSIF x =- 17484 THEN
            exp_f := 0;
        ELSIF x =- 17483 THEN
            exp_f := 0;
        ELSIF x =- 17482 THEN
            exp_f := 0;
        ELSIF x =- 17481 THEN
            exp_f := 0;
        ELSIF x =- 17480 THEN
            exp_f := 0;
        ELSIF x =- 17479 THEN
            exp_f := 0;
        ELSIF x =- 17478 THEN
            exp_f := 0;
        ELSIF x =- 17477 THEN
            exp_f := 0;
        ELSIF x =- 17476 THEN
            exp_f := 0;
        ELSIF x =- 17475 THEN
            exp_f := 0;
        ELSIF x =- 17474 THEN
            exp_f := 0;
        ELSIF x =- 17473 THEN
            exp_f := 0;
        ELSIF x =- 17472 THEN
            exp_f := 0;
        ELSIF x =- 17471 THEN
            exp_f := 0;
        ELSIF x =- 17470 THEN
            exp_f := 0;
        ELSIF x =- 17469 THEN
            exp_f := 0;
        ELSIF x =- 17468 THEN
            exp_f := 0;
        ELSIF x =- 17467 THEN
            exp_f := 0;
        ELSIF x =- 17466 THEN
            exp_f := 0;
        ELSIF x =- 17465 THEN
            exp_f := 0;
        ELSIF x =- 17464 THEN
            exp_f := 0;
        ELSIF x =- 17463 THEN
            exp_f := 0;
        ELSIF x =- 17462 THEN
            exp_f := 0;
        ELSIF x =- 17461 THEN
            exp_f := 0;
        ELSIF x =- 17460 THEN
            exp_f := 0;
        ELSIF x =- 17459 THEN
            exp_f := 0;
        ELSIF x =- 17458 THEN
            exp_f := 0;
        ELSIF x =- 17457 THEN
            exp_f := 0;
        ELSIF x =- 17456 THEN
            exp_f := 0;
        ELSIF x =- 17455 THEN
            exp_f := 0;
        ELSIF x =- 17454 THEN
            exp_f := 0;
        ELSIF x =- 17453 THEN
            exp_f := 0;
        ELSIF x =- 17452 THEN
            exp_f := 0;
        ELSIF x =- 17451 THEN
            exp_f := 0;
        ELSIF x =- 17450 THEN
            exp_f := 0;
        ELSIF x =- 17449 THEN
            exp_f := 0;
        ELSIF x =- 17448 THEN
            exp_f := 0;
        ELSIF x =- 17447 THEN
            exp_f := 0;
        ELSIF x =- 17446 THEN
            exp_f := 0;
        ELSIF x =- 17445 THEN
            exp_f := 0;
        ELSIF x =- 17444 THEN
            exp_f := 0;
        ELSIF x =- 17443 THEN
            exp_f := 0;
        ELSIF x =- 17442 THEN
            exp_f := 0;
        ELSIF x =- 17441 THEN
            exp_f := 0;
        ELSIF x =- 17440 THEN
            exp_f := 0;
        ELSIF x =- 17439 THEN
            exp_f := 0;
        ELSIF x =- 17438 THEN
            exp_f := 0;
        ELSIF x =- 17437 THEN
            exp_f := 0;
        ELSIF x =- 17436 THEN
            exp_f := 0;
        ELSIF x =- 17435 THEN
            exp_f := 0;
        ELSIF x =- 17434 THEN
            exp_f := 0;
        ELSIF x =- 17433 THEN
            exp_f := 0;
        ELSIF x =- 17432 THEN
            exp_f := 0;
        ELSIF x =- 17431 THEN
            exp_f := 0;
        ELSIF x =- 17430 THEN
            exp_f := 0;
        ELSIF x =- 17429 THEN
            exp_f := 0;
        ELSIF x =- 17428 THEN
            exp_f := 0;
        ELSIF x =- 17427 THEN
            exp_f := 0;
        ELSIF x =- 17426 THEN
            exp_f := 0;
        ELSIF x =- 17425 THEN
            exp_f := 0;
        ELSIF x =- 17424 THEN
            exp_f := 0;
        ELSIF x =- 17423 THEN
            exp_f := 0;
        ELSIF x =- 17422 THEN
            exp_f := 0;
        ELSIF x =- 17421 THEN
            exp_f := 0;
        ELSIF x =- 17420 THEN
            exp_f := 0;
        ELSIF x =- 17419 THEN
            exp_f := 0;
        ELSIF x =- 17418 THEN
            exp_f := 0;
        ELSIF x =- 17417 THEN
            exp_f := 0;
        ELSIF x =- 17416 THEN
            exp_f := 0;
        ELSIF x =- 17415 THEN
            exp_f := 0;
        ELSIF x =- 17414 THEN
            exp_f := 0;
        ELSIF x =- 17413 THEN
            exp_f := 0;
        ELSIF x =- 17412 THEN
            exp_f := 0;
        ELSIF x =- 17411 THEN
            exp_f := 0;
        ELSIF x =- 17410 THEN
            exp_f := 0;
        ELSIF x =- 17409 THEN
            exp_f := 0;
        ELSIF x =- 17408 THEN
            exp_f := 0;
        ELSIF x =- 17407 THEN
            exp_f := 0;
        ELSIF x =- 17406 THEN
            exp_f := 0;
        ELSIF x =- 17405 THEN
            exp_f := 0;
        ELSIF x =- 17404 THEN
            exp_f := 0;
        ELSIF x =- 17403 THEN
            exp_f := 0;
        ELSIF x =- 17402 THEN
            exp_f := 0;
        ELSIF x =- 17401 THEN
            exp_f := 0;
        ELSIF x =- 17400 THEN
            exp_f := 0;
        ELSIF x =- 17399 THEN
            exp_f := 0;
        ELSIF x =- 17398 THEN
            exp_f := 0;
        ELSIF x =- 17397 THEN
            exp_f := 0;
        ELSIF x =- 17396 THEN
            exp_f := 0;
        ELSIF x =- 17395 THEN
            exp_f := 0;
        ELSIF x =- 17394 THEN
            exp_f := 0;
        ELSIF x =- 17393 THEN
            exp_f := 0;
        ELSIF x =- 17392 THEN
            exp_f := 0;
        ELSIF x =- 17391 THEN
            exp_f := 0;
        ELSIF x =- 17390 THEN
            exp_f := 0;
        ELSIF x =- 17389 THEN
            exp_f := 0;
        ELSIF x =- 17388 THEN
            exp_f := 0;
        ELSIF x =- 17387 THEN
            exp_f := 0;
        ELSIF x =- 17386 THEN
            exp_f := 0;
        ELSIF x =- 17385 THEN
            exp_f := 0;
        ELSIF x =- 17384 THEN
            exp_f := 0;
        ELSIF x =- 17383 THEN
            exp_f := 0;
        ELSIF x =- 17382 THEN
            exp_f := 0;
        ELSIF x =- 17381 THEN
            exp_f := 0;
        ELSIF x =- 17380 THEN
            exp_f := 0;
        ELSIF x =- 17379 THEN
            exp_f := 0;
        ELSIF x =- 17378 THEN
            exp_f := 0;
        ELSIF x =- 17377 THEN
            exp_f := 0;
        ELSIF x =- 17376 THEN
            exp_f := 0;
        ELSIF x =- 17375 THEN
            exp_f := 0;
        ELSIF x =- 17374 THEN
            exp_f := 0;
        ELSIF x =- 17373 THEN
            exp_f := 0;
        ELSIF x =- 17372 THEN
            exp_f := 0;
        ELSIF x =- 17371 THEN
            exp_f := 0;
        ELSIF x =- 17370 THEN
            exp_f := 0;
        ELSIF x =- 17369 THEN
            exp_f := 0;
        ELSIF x =- 17368 THEN
            exp_f := 0;
        ELSIF x =- 17367 THEN
            exp_f := 0;
        ELSIF x =- 17366 THEN
            exp_f := 0;
        ELSIF x =- 17365 THEN
            exp_f := 0;
        ELSIF x =- 17364 THEN
            exp_f := 0;
        ELSIF x =- 17363 THEN
            exp_f := 0;
        ELSIF x =- 17362 THEN
            exp_f := 0;
        ELSIF x =- 17361 THEN
            exp_f := 0;
        ELSIF x =- 17360 THEN
            exp_f := 0;
        ELSIF x =- 17359 THEN
            exp_f := 0;
        ELSIF x =- 17358 THEN
            exp_f := 0;
        ELSIF x =- 17357 THEN
            exp_f := 0;
        ELSIF x =- 17356 THEN
            exp_f := 0;
        ELSIF x =- 17355 THEN
            exp_f := 0;
        ELSIF x =- 17354 THEN
            exp_f := 0;
        ELSIF x =- 17353 THEN
            exp_f := 0;
        ELSIF x =- 17352 THEN
            exp_f := 0;
        ELSIF x =- 17351 THEN
            exp_f := 0;
        ELSIF x =- 17350 THEN
            exp_f := 0;
        ELSIF x =- 17349 THEN
            exp_f := 0;
        ELSIF x =- 17348 THEN
            exp_f := 0;
        ELSIF x =- 17347 THEN
            exp_f := 0;
        ELSIF x =- 17346 THEN
            exp_f := 0;
        ELSIF x =- 17345 THEN
            exp_f := 0;
        ELSIF x =- 17344 THEN
            exp_f := 0;
        ELSIF x =- 17343 THEN
            exp_f := 0;
        ELSIF x =- 17342 THEN
            exp_f := 0;
        ELSIF x =- 17341 THEN
            exp_f := 0;
        ELSIF x =- 17340 THEN
            exp_f := 0;
        ELSIF x =- 17339 THEN
            exp_f := 0;
        ELSIF x =- 17338 THEN
            exp_f := 0;
        ELSIF x =- 17337 THEN
            exp_f := 0;
        ELSIF x =- 17336 THEN
            exp_f := 0;
        ELSIF x =- 17335 THEN
            exp_f := 0;
        ELSIF x =- 17334 THEN
            exp_f := 0;
        ELSIF x =- 17333 THEN
            exp_f := 0;
        ELSIF x =- 17332 THEN
            exp_f := 0;
        ELSIF x =- 17331 THEN
            exp_f := 0;
        ELSIF x =- 17330 THEN
            exp_f := 0;
        ELSIF x =- 17329 THEN
            exp_f := 0;
        ELSIF x =- 17328 THEN
            exp_f := 0;
        ELSIF x =- 17327 THEN
            exp_f := 0;
        ELSIF x =- 17326 THEN
            exp_f := 0;
        ELSIF x =- 17325 THEN
            exp_f := 0;
        ELSIF x =- 17324 THEN
            exp_f := 0;
        ELSIF x =- 17323 THEN
            exp_f := 0;
        ELSIF x =- 17322 THEN
            exp_f := 0;
        ELSIF x =- 17321 THEN
            exp_f := 0;
        ELSIF x =- 17320 THEN
            exp_f := 0;
        ELSIF x =- 17319 THEN
            exp_f := 0;
        ELSIF x =- 17318 THEN
            exp_f := 0;
        ELSIF x =- 17317 THEN
            exp_f := 0;
        ELSIF x =- 17316 THEN
            exp_f := 0;
        ELSIF x =- 17315 THEN
            exp_f := 0;
        ELSIF x =- 17314 THEN
            exp_f := 0;
        ELSIF x =- 17313 THEN
            exp_f := 0;
        ELSIF x =- 17312 THEN
            exp_f := 0;
        ELSIF x =- 17311 THEN
            exp_f := 0;
        ELSIF x =- 17310 THEN
            exp_f := 0;
        ELSIF x =- 17309 THEN
            exp_f := 0;
        ELSIF x =- 17308 THEN
            exp_f := 0;
        ELSIF x =- 17307 THEN
            exp_f := 0;
        ELSIF x =- 17306 THEN
            exp_f := 0;
        ELSIF x =- 17305 THEN
            exp_f := 0;
        ELSIF x =- 17304 THEN
            exp_f := 0;
        ELSIF x =- 17303 THEN
            exp_f := 0;
        ELSIF x =- 17302 THEN
            exp_f := 0;
        ELSIF x =- 17301 THEN
            exp_f := 0;
        ELSIF x =- 17300 THEN
            exp_f := 0;
        ELSIF x =- 17299 THEN
            exp_f := 0;
        ELSIF x =- 17298 THEN
            exp_f := 0;
        ELSIF x =- 17297 THEN
            exp_f := 0;
        ELSIF x =- 17296 THEN
            exp_f := 0;
        ELSIF x =- 17295 THEN
            exp_f := 0;
        ELSIF x =- 17294 THEN
            exp_f := 0;
        ELSIF x =- 17293 THEN
            exp_f := 0;
        ELSIF x =- 17292 THEN
            exp_f := 0;
        ELSIF x =- 17291 THEN
            exp_f := 0;
        ELSIF x =- 17290 THEN
            exp_f := 0;
        ELSIF x =- 17289 THEN
            exp_f := 0;
        ELSIF x =- 17288 THEN
            exp_f := 0;
        ELSIF x =- 17287 THEN
            exp_f := 0;
        ELSIF x =- 17286 THEN
            exp_f := 0;
        ELSIF x =- 17285 THEN
            exp_f := 0;
        ELSIF x =- 17284 THEN
            exp_f := 0;
        ELSIF x =- 17283 THEN
            exp_f := 0;
        ELSIF x =- 17282 THEN
            exp_f := 0;
        ELSIF x =- 17281 THEN
            exp_f := 0;
        ELSIF x =- 17280 THEN
            exp_f := 0;
        ELSIF x =- 17279 THEN
            exp_f := 0;
        ELSIF x =- 17278 THEN
            exp_f := 0;
        ELSIF x =- 17277 THEN
            exp_f := 0;
        ELSIF x =- 17276 THEN
            exp_f := 0;
        ELSIF x =- 17275 THEN
            exp_f := 0;
        ELSIF x =- 17274 THEN
            exp_f := 0;
        ELSIF x =- 17273 THEN
            exp_f := 0;
        ELSIF x =- 17272 THEN
            exp_f := 0;
        ELSIF x =- 17271 THEN
            exp_f := 0;
        ELSIF x =- 17270 THEN
            exp_f := 0;
        ELSIF x =- 17269 THEN
            exp_f := 0;
        ELSIF x =- 17268 THEN
            exp_f := 0;
        ELSIF x =- 17267 THEN
            exp_f := 0;
        ELSIF x =- 17266 THEN
            exp_f := 0;
        ELSIF x =- 17265 THEN
            exp_f := 0;
        ELSIF x =- 17264 THEN
            exp_f := 0;
        ELSIF x =- 17263 THEN
            exp_f := 0;
        ELSIF x =- 17262 THEN
            exp_f := 0;
        ELSIF x =- 17261 THEN
            exp_f := 0;
        ELSIF x =- 17260 THEN
            exp_f := 0;
        ELSIF x =- 17259 THEN
            exp_f := 0;
        ELSIF x =- 17258 THEN
            exp_f := 0;
        ELSIF x =- 17257 THEN
            exp_f := 0;
        ELSIF x =- 17256 THEN
            exp_f := 0;
        ELSIF x =- 17255 THEN
            exp_f := 0;
        ELSIF x =- 17254 THEN
            exp_f := 0;
        ELSIF x =- 17253 THEN
            exp_f := 0;
        ELSIF x =- 17252 THEN
            exp_f := 0;
        ELSIF x =- 17251 THEN
            exp_f := 0;
        ELSIF x =- 17250 THEN
            exp_f := 0;
        ELSIF x =- 17249 THEN
            exp_f := 0;
        ELSIF x =- 17248 THEN
            exp_f := 0;
        ELSIF x =- 17247 THEN
            exp_f := 0;
        ELSIF x =- 17246 THEN
            exp_f := 0;
        ELSIF x =- 17245 THEN
            exp_f := 0;
        ELSIF x =- 17244 THEN
            exp_f := 0;
        ELSIF x =- 17243 THEN
            exp_f := 0;
        ELSIF x =- 17242 THEN
            exp_f := 0;
        ELSIF x =- 17241 THEN
            exp_f := 0;
        ELSIF x =- 17240 THEN
            exp_f := 0;
        ELSIF x =- 17239 THEN
            exp_f := 0;
        ELSIF x =- 17238 THEN
            exp_f := 0;
        ELSIF x =- 17237 THEN
            exp_f := 0;
        ELSIF x =- 17236 THEN
            exp_f := 0;
        ELSIF x =- 17235 THEN
            exp_f := 0;
        ELSIF x =- 17234 THEN
            exp_f := 0;
        ELSIF x =- 17233 THEN
            exp_f := 0;
        ELSIF x =- 17232 THEN
            exp_f := 0;
        ELSIF x =- 17231 THEN
            exp_f := 0;
        ELSIF x =- 17230 THEN
            exp_f := 0;
        ELSIF x =- 17229 THEN
            exp_f := 0;
        ELSIF x =- 17228 THEN
            exp_f := 0;
        ELSIF x =- 17227 THEN
            exp_f := 0;
        ELSIF x =- 17226 THEN
            exp_f := 0;
        ELSIF x =- 17225 THEN
            exp_f := 0;
        ELSIF x =- 17224 THEN
            exp_f := 0;
        ELSIF x =- 17223 THEN
            exp_f := 0;
        ELSIF x =- 17222 THEN
            exp_f := 0;
        ELSIF x =- 17221 THEN
            exp_f := 0;
        ELSIF x =- 17220 THEN
            exp_f := 0;
        ELSIF x =- 17219 THEN
            exp_f := 0;
        ELSIF x =- 17218 THEN
            exp_f := 0;
        ELSIF x =- 17217 THEN
            exp_f := 0;
        ELSIF x =- 17216 THEN
            exp_f := 0;
        ELSIF x =- 17215 THEN
            exp_f := 0;
        ELSIF x =- 17214 THEN
            exp_f := 0;
        ELSIF x =- 17213 THEN
            exp_f := 0;
        ELSIF x =- 17212 THEN
            exp_f := 0;
        ELSIF x =- 17211 THEN
            exp_f := 0;
        ELSIF x =- 17210 THEN
            exp_f := 0;
        ELSIF x =- 17209 THEN
            exp_f := 0;
        ELSIF x =- 17208 THEN
            exp_f := 0;
        ELSIF x =- 17207 THEN
            exp_f := 0;
        ELSIF x =- 17206 THEN
            exp_f := 0;
        ELSIF x =- 17205 THEN
            exp_f := 0;
        ELSIF x =- 17204 THEN
            exp_f := 0;
        ELSIF x =- 17203 THEN
            exp_f := 0;
        ELSIF x =- 17202 THEN
            exp_f := 0;
        ELSIF x =- 17201 THEN
            exp_f := 0;
        ELSIF x =- 17200 THEN
            exp_f := 0;
        ELSIF x =- 17199 THEN
            exp_f := 0;
        ELSIF x =- 17198 THEN
            exp_f := 0;
        ELSIF x =- 17197 THEN
            exp_f := 0;
        ELSIF x =- 17196 THEN
            exp_f := 0;
        ELSIF x =- 17195 THEN
            exp_f := 0;
        ELSIF x =- 17194 THEN
            exp_f := 0;
        ELSIF x =- 17193 THEN
            exp_f := 0;
        ELSIF x =- 17192 THEN
            exp_f := 0;
        ELSIF x =- 17191 THEN
            exp_f := 0;
        ELSIF x =- 17190 THEN
            exp_f := 0;
        ELSIF x =- 17189 THEN
            exp_f := 0;
        ELSIF x =- 17188 THEN
            exp_f := 0;
        ELSIF x =- 17187 THEN
            exp_f := 0;
        ELSIF x =- 17186 THEN
            exp_f := 0;
        ELSIF x =- 17185 THEN
            exp_f := 0;
        ELSIF x =- 17184 THEN
            exp_f := 0;
        ELSIF x =- 17183 THEN
            exp_f := 0;
        ELSIF x =- 17182 THEN
            exp_f := 0;
        ELSIF x =- 17181 THEN
            exp_f := 0;
        ELSIF x =- 17180 THEN
            exp_f := 0;
        ELSIF x =- 17179 THEN
            exp_f := 0;
        ELSIF x =- 17178 THEN
            exp_f := 0;
        ELSIF x =- 17177 THEN
            exp_f := 0;
        ELSIF x =- 17176 THEN
            exp_f := 0;
        ELSIF x =- 17175 THEN
            exp_f := 0;
        ELSIF x =- 17174 THEN
            exp_f := 0;
        ELSIF x =- 17173 THEN
            exp_f := 0;
        ELSIF x =- 17172 THEN
            exp_f := 0;
        ELSIF x =- 17171 THEN
            exp_f := 0;
        ELSIF x =- 17170 THEN
            exp_f := 0;
        ELSIF x =- 17169 THEN
            exp_f := 0;
        ELSIF x =- 17168 THEN
            exp_f := 0;
        ELSIF x =- 17167 THEN
            exp_f := 0;
        ELSIF x =- 17166 THEN
            exp_f := 0;
        ELSIF x =- 17165 THEN
            exp_f := 0;
        ELSIF x =- 17164 THEN
            exp_f := 0;
        ELSIF x =- 17163 THEN
            exp_f := 0;
        ELSIF x =- 17162 THEN
            exp_f := 0;
        ELSIF x =- 17161 THEN
            exp_f := 0;
        ELSIF x =- 17160 THEN
            exp_f := 0;
        ELSIF x =- 17159 THEN
            exp_f := 0;
        ELSIF x =- 17158 THEN
            exp_f := 0;
        ELSIF x =- 17157 THEN
            exp_f := 0;
        ELSIF x =- 17156 THEN
            exp_f := 0;
        ELSIF x =- 17155 THEN
            exp_f := 0;
        ELSIF x =- 17154 THEN
            exp_f := 0;
        ELSIF x =- 17153 THEN
            exp_f := 0;
        ELSIF x =- 17152 THEN
            exp_f := 0;
        ELSIF x =- 17151 THEN
            exp_f := 0;
        ELSIF x =- 17150 THEN
            exp_f := 0;
        ELSIF x =- 17149 THEN
            exp_f := 0;
        ELSIF x =- 17148 THEN
            exp_f := 0;
        ELSIF x =- 17147 THEN
            exp_f := 0;
        ELSIF x =- 17146 THEN
            exp_f := 0;
        ELSIF x =- 17145 THEN
            exp_f := 0;
        ELSIF x =- 17144 THEN
            exp_f := 0;
        ELSIF x =- 17143 THEN
            exp_f := 0;
        ELSIF x =- 17142 THEN
            exp_f := 0;
        ELSIF x =- 17141 THEN
            exp_f := 0;
        ELSIF x =- 17140 THEN
            exp_f := 0;
        ELSIF x =- 17139 THEN
            exp_f := 0;
        ELSIF x =- 17138 THEN
            exp_f := 0;
        ELSIF x =- 17137 THEN
            exp_f := 0;
        ELSIF x =- 17136 THEN
            exp_f := 0;
        ELSIF x =- 17135 THEN
            exp_f := 0;
        ELSIF x =- 17134 THEN
            exp_f := 0;
        ELSIF x =- 17133 THEN
            exp_f := 0;
        ELSIF x =- 17132 THEN
            exp_f := 0;
        ELSIF x =- 17131 THEN
            exp_f := 0;
        ELSIF x =- 17130 THEN
            exp_f := 0;
        ELSIF x =- 17129 THEN
            exp_f := 0;
        ELSIF x =- 17128 THEN
            exp_f := 0;
        ELSIF x =- 17127 THEN
            exp_f := 0;
        ELSIF x =- 17126 THEN
            exp_f := 0;
        ELSIF x =- 17125 THEN
            exp_f := 0;
        ELSIF x =- 17124 THEN
            exp_f := 0;
        ELSIF x =- 17123 THEN
            exp_f := 0;
        ELSIF x =- 17122 THEN
            exp_f := 0;
        ELSIF x =- 17121 THEN
            exp_f := 0;
        ELSIF x =- 17120 THEN
            exp_f := 0;
        ELSIF x =- 17119 THEN
            exp_f := 0;
        ELSIF x =- 17118 THEN
            exp_f := 0;
        ELSIF x =- 17117 THEN
            exp_f := 0;
        ELSIF x =- 17116 THEN
            exp_f := 0;
        ELSIF x =- 17115 THEN
            exp_f := 0;
        ELSIF x =- 17114 THEN
            exp_f := 0;
        ELSIF x =- 17113 THEN
            exp_f := 0;
        ELSIF x =- 17112 THEN
            exp_f := 0;
        ELSIF x =- 17111 THEN
            exp_f := 0;
        ELSIF x =- 17110 THEN
            exp_f := 0;
        ELSIF x =- 17109 THEN
            exp_f := 0;
        ELSIF x =- 17108 THEN
            exp_f := 0;
        ELSIF x =- 17107 THEN
            exp_f := 0;
        ELSIF x =- 17106 THEN
            exp_f := 0;
        ELSIF x =- 17105 THEN
            exp_f := 0;
        ELSIF x =- 17104 THEN
            exp_f := 0;
        ELSIF x =- 17103 THEN
            exp_f := 0;
        ELSIF x =- 17102 THEN
            exp_f := 0;
        ELSIF x =- 17101 THEN
            exp_f := 0;
        ELSIF x =- 17100 THEN
            exp_f := 0;
        ELSIF x =- 17099 THEN
            exp_f := 0;
        ELSIF x =- 17098 THEN
            exp_f := 0;
        ELSIF x =- 17097 THEN
            exp_f := 0;
        ELSIF x =- 17096 THEN
            exp_f := 0;
        ELSIF x =- 17095 THEN
            exp_f := 0;
        ELSIF x =- 17094 THEN
            exp_f := 0;
        ELSIF x =- 17093 THEN
            exp_f := 0;
        ELSIF x =- 17092 THEN
            exp_f := 0;
        ELSIF x =- 17091 THEN
            exp_f := 0;
        ELSIF x =- 17090 THEN
            exp_f := 0;
        ELSIF x =- 17089 THEN
            exp_f := 0;
        ELSIF x =- 17088 THEN
            exp_f := 0;
        ELSIF x =- 17087 THEN
            exp_f := 0;
        ELSIF x =- 17086 THEN
            exp_f := 0;
        ELSIF x =- 17085 THEN
            exp_f := 0;
        ELSIF x =- 17084 THEN
            exp_f := 0;
        ELSIF x =- 17083 THEN
            exp_f := 0;
        ELSIF x =- 17082 THEN
            exp_f := 0;
        ELSIF x =- 17081 THEN
            exp_f := 0;
        ELSIF x =- 17080 THEN
            exp_f := 0;
        ELSIF x =- 17079 THEN
            exp_f := 0;
        ELSIF x =- 17078 THEN
            exp_f := 0;
        ELSIF x =- 17077 THEN
            exp_f := 0;
        ELSIF x =- 17076 THEN
            exp_f := 0;
        ELSIF x =- 17075 THEN
            exp_f := 0;
        ELSIF x =- 17074 THEN
            exp_f := 0;
        ELSIF x =- 17073 THEN
            exp_f := 0;
        ELSIF x =- 17072 THEN
            exp_f := 0;
        ELSIF x =- 17071 THEN
            exp_f := 0;
        ELSIF x =- 17070 THEN
            exp_f := 0;
        ELSIF x =- 17069 THEN
            exp_f := 0;
        ELSIF x =- 17068 THEN
            exp_f := 0;
        ELSIF x =- 17067 THEN
            exp_f := 0;
        ELSIF x =- 17066 THEN
            exp_f := 0;
        ELSIF x =- 17065 THEN
            exp_f := 0;
        ELSIF x =- 17064 THEN
            exp_f := 0;
        ELSIF x =- 17063 THEN
            exp_f := 0;
        ELSIF x =- 17062 THEN
            exp_f := 0;
        ELSIF x =- 17061 THEN
            exp_f := 0;
        ELSIF x =- 17060 THEN
            exp_f := 0;
        ELSIF x =- 17059 THEN
            exp_f := 0;
        ELSIF x =- 17058 THEN
            exp_f := 0;
        ELSIF x =- 17057 THEN
            exp_f := 0;
        ELSIF x =- 17056 THEN
            exp_f := 0;
        ELSIF x =- 17055 THEN
            exp_f := 0;
        ELSIF x =- 17054 THEN
            exp_f := 0;
        ELSIF x =- 17053 THEN
            exp_f := 0;
        ELSIF x =- 17052 THEN
            exp_f := 0;
        ELSIF x =- 17051 THEN
            exp_f := 0;
        ELSIF x =- 17050 THEN
            exp_f := 0;
        ELSIF x =- 17049 THEN
            exp_f := 0;
        ELSIF x =- 17048 THEN
            exp_f := 0;
        ELSIF x =- 17047 THEN
            exp_f := 0;
        ELSIF x =- 17046 THEN
            exp_f := 0;
        ELSIF x =- 17045 THEN
            exp_f := 0;
        ELSIF x =- 17044 THEN
            exp_f := 0;
        ELSIF x =- 17043 THEN
            exp_f := 0;
        ELSIF x =- 17042 THEN
            exp_f := 0;
        ELSIF x =- 17041 THEN
            exp_f := 0;
        ELSIF x =- 17040 THEN
            exp_f := 0;
        ELSIF x =- 17039 THEN
            exp_f := 0;
        ELSIF x =- 17038 THEN
            exp_f := 0;
        ELSIF x =- 17037 THEN
            exp_f := 0;
        ELSIF x =- 17036 THEN
            exp_f := 0;
        ELSIF x =- 17035 THEN
            exp_f := 0;
        ELSIF x =- 17034 THEN
            exp_f := 0;
        ELSIF x =- 17033 THEN
            exp_f := 0;
        ELSIF x =- 17032 THEN
            exp_f := 0;
        ELSIF x =- 17031 THEN
            exp_f := 0;
        ELSIF x =- 17030 THEN
            exp_f := 0;
        ELSIF x =- 17029 THEN
            exp_f := 0;
        ELSIF x =- 17028 THEN
            exp_f := 0;
        ELSIF x =- 17027 THEN
            exp_f := 0;
        ELSIF x =- 17026 THEN
            exp_f := 0;
        ELSIF x =- 17025 THEN
            exp_f := 0;
        ELSIF x =- 17024 THEN
            exp_f := 0;
        ELSIF x =- 17023 THEN
            exp_f := 0;
        ELSIF x =- 17022 THEN
            exp_f := 0;
        ELSIF x =- 17021 THEN
            exp_f := 0;
        ELSIF x =- 17020 THEN
            exp_f := 0;
        ELSIF x =- 17019 THEN
            exp_f := 0;
        ELSIF x =- 17018 THEN
            exp_f := 0;
        ELSIF x =- 17017 THEN
            exp_f := 0;
        ELSIF x =- 17016 THEN
            exp_f := 0;
        ELSIF x =- 17015 THEN
            exp_f := 0;
        ELSIF x =- 17014 THEN
            exp_f := 0;
        ELSIF x =- 17013 THEN
            exp_f := 0;
        ELSIF x =- 17012 THEN
            exp_f := 0;
        ELSIF x =- 17011 THEN
            exp_f := 0;
        ELSIF x =- 17010 THEN
            exp_f := 0;
        ELSIF x =- 17009 THEN
            exp_f := 0;
        ELSIF x =- 17008 THEN
            exp_f := 0;
        ELSIF x =- 17007 THEN
            exp_f := 0;
        ELSIF x =- 17006 THEN
            exp_f := 0;
        ELSIF x =- 17005 THEN
            exp_f := 0;
        ELSIF x =- 17004 THEN
            exp_f := 0;
        ELSIF x =- 17003 THEN
            exp_f := 0;
        ELSIF x =- 17002 THEN
            exp_f := 0;
        ELSIF x =- 17001 THEN
            exp_f := 0;
        ELSIF x =- 17000 THEN
            exp_f := 0;
        ELSIF x =- 16999 THEN
            exp_f := 0;
        ELSIF x =- 16998 THEN
            exp_f := 0;
        ELSIF x =- 16997 THEN
            exp_f := 0;
        ELSIF x =- 16996 THEN
            exp_f := 0;
        ELSIF x =- 16995 THEN
            exp_f := 0;
        ELSIF x =- 16994 THEN
            exp_f := 0;
        ELSIF x =- 16993 THEN
            exp_f := 0;
        ELSIF x =- 16992 THEN
            exp_f := 0;
        ELSIF x =- 16991 THEN
            exp_f := 0;
        ELSIF x =- 16990 THEN
            exp_f := 0;
        ELSIF x =- 16989 THEN
            exp_f := 0;
        ELSIF x =- 16988 THEN
            exp_f := 0;
        ELSIF x =- 16987 THEN
            exp_f := 0;
        ELSIF x =- 16986 THEN
            exp_f := 0;
        ELSIF x =- 16985 THEN
            exp_f := 0;
        ELSIF x =- 16984 THEN
            exp_f := 0;
        ELSIF x =- 16983 THEN
            exp_f := 0;
        ELSIF x =- 16982 THEN
            exp_f := 0;
        ELSIF x =- 16981 THEN
            exp_f := 0;
        ELSIF x =- 16980 THEN
            exp_f := 0;
        ELSIF x =- 16979 THEN
            exp_f := 0;
        ELSIF x =- 16978 THEN
            exp_f := 0;
        ELSIF x =- 16977 THEN
            exp_f := 0;
        ELSIF x =- 16976 THEN
            exp_f := 0;
        ELSIF x =- 16975 THEN
            exp_f := 0;
        ELSIF x =- 16974 THEN
            exp_f := 0;
        ELSIF x =- 16973 THEN
            exp_f := 0;
        ELSIF x =- 16972 THEN
            exp_f := 0;
        ELSIF x =- 16971 THEN
            exp_f := 0;
        ELSIF x =- 16970 THEN
            exp_f := 0;
        ELSIF x =- 16969 THEN
            exp_f := 0;
        ELSIF x =- 16968 THEN
            exp_f := 0;
        ELSIF x =- 16967 THEN
            exp_f := 0;
        ELSIF x =- 16966 THEN
            exp_f := 0;
        ELSIF x =- 16965 THEN
            exp_f := 0;
        ELSIF x =- 16964 THEN
            exp_f := 0;
        ELSIF x =- 16963 THEN
            exp_f := 0;
        ELSIF x =- 16962 THEN
            exp_f := 0;
        ELSIF x =- 16961 THEN
            exp_f := 0;
        ELSIF x =- 16960 THEN
            exp_f := 0;
        ELSIF x =- 16959 THEN
            exp_f := 0;
        ELSIF x =- 16958 THEN
            exp_f := 0;
        ELSIF x =- 16957 THEN
            exp_f := 0;
        ELSIF x =- 16956 THEN
            exp_f := 0;
        ELSIF x =- 16955 THEN
            exp_f := 0;
        ELSIF x =- 16954 THEN
            exp_f := 0;
        ELSIF x =- 16953 THEN
            exp_f := 0;
        ELSIF x =- 16952 THEN
            exp_f := 0;
        ELSIF x =- 16951 THEN
            exp_f := 0;
        ELSIF x =- 16950 THEN
            exp_f := 0;
        ELSIF x =- 16949 THEN
            exp_f := 0;
        ELSIF x =- 16948 THEN
            exp_f := 0;
        ELSIF x =- 16947 THEN
            exp_f := 0;
        ELSIF x =- 16946 THEN
            exp_f := 0;
        ELSIF x =- 16945 THEN
            exp_f := 0;
        ELSIF x =- 16944 THEN
            exp_f := 0;
        ELSIF x =- 16943 THEN
            exp_f := 0;
        ELSIF x =- 16942 THEN
            exp_f := 0;
        ELSIF x =- 16941 THEN
            exp_f := 0;
        ELSIF x =- 16940 THEN
            exp_f := 0;
        ELSIF x =- 16939 THEN
            exp_f := 0;
        ELSIF x =- 16938 THEN
            exp_f := 0;
        ELSIF x =- 16937 THEN
            exp_f := 0;
        ELSIF x =- 16936 THEN
            exp_f := 0;
        ELSIF x =- 16935 THEN
            exp_f := 0;
        ELSIF x =- 16934 THEN
            exp_f := 0;
        ELSIF x =- 16933 THEN
            exp_f := 0;
        ELSIF x =- 16932 THEN
            exp_f := 0;
        ELSIF x =- 16931 THEN
            exp_f := 0;
        ELSIF x =- 16930 THEN
            exp_f := 0;
        ELSIF x =- 16929 THEN
            exp_f := 0;
        ELSIF x =- 16928 THEN
            exp_f := 0;
        ELSIF x =- 16927 THEN
            exp_f := 0;
        ELSIF x =- 16926 THEN
            exp_f := 0;
        ELSIF x =- 16925 THEN
            exp_f := 0;
        ELSIF x =- 16924 THEN
            exp_f := 0;
        ELSIF x =- 16923 THEN
            exp_f := 0;
        ELSIF x =- 16922 THEN
            exp_f := 0;
        ELSIF x =- 16921 THEN
            exp_f := 0;
        ELSIF x =- 16920 THEN
            exp_f := 0;
        ELSIF x =- 16919 THEN
            exp_f := 0;
        ELSIF x =- 16918 THEN
            exp_f := 0;
        ELSIF x =- 16917 THEN
            exp_f := 0;
        ELSIF x =- 16916 THEN
            exp_f := 0;
        ELSIF x =- 16915 THEN
            exp_f := 0;
        ELSIF x =- 16914 THEN
            exp_f := 0;
        ELSIF x =- 16913 THEN
            exp_f := 0;
        ELSIF x =- 16912 THEN
            exp_f := 0;
        ELSIF x =- 16911 THEN
            exp_f := 0;
        ELSIF x =- 16910 THEN
            exp_f := 0;
        ELSIF x =- 16909 THEN
            exp_f := 0;
        ELSIF x =- 16908 THEN
            exp_f := 0;
        ELSIF x =- 16907 THEN
            exp_f := 0;
        ELSIF x =- 16906 THEN
            exp_f := 0;
        ELSIF x =- 16905 THEN
            exp_f := 0;
        ELSIF x =- 16904 THEN
            exp_f := 0;
        ELSIF x =- 16903 THEN
            exp_f := 0;
        ELSIF x =- 16902 THEN
            exp_f := 0;
        ELSIF x =- 16901 THEN
            exp_f := 0;
        ELSIF x =- 16900 THEN
            exp_f := 0;
        ELSIF x =- 16899 THEN
            exp_f := 0;
        ELSIF x =- 16898 THEN
            exp_f := 0;
        ELSIF x =- 16897 THEN
            exp_f := 0;
        ELSIF x =- 16896 THEN
            exp_f := 0;
        ELSIF x =- 16895 THEN
            exp_f := 1;
        ELSIF x =- 16894 THEN
            exp_f := 1;
        ELSIF x =- 16893 THEN
            exp_f := 1;
        ELSIF x =- 16892 THEN
            exp_f := 1;
        ELSIF x =- 16891 THEN
            exp_f := 1;
        ELSIF x =- 16890 THEN
            exp_f := 1;
        ELSIF x =- 16889 THEN
            exp_f := 1;
        ELSIF x =- 16888 THEN
            exp_f := 1;
        ELSIF x =- 16887 THEN
            exp_f := 1;
        ELSIF x =- 16886 THEN
            exp_f := 1;
        ELSIF x =- 16885 THEN
            exp_f := 1;
        ELSIF x =- 16884 THEN
            exp_f := 1;
        ELSIF x =- 16883 THEN
            exp_f := 1;
        ELSIF x =- 16882 THEN
            exp_f := 1;
        ELSIF x =- 16881 THEN
            exp_f := 1;
        ELSIF x =- 16880 THEN
            exp_f := 1;
        ELSIF x =- 16879 THEN
            exp_f := 1;
        ELSIF x =- 16878 THEN
            exp_f := 1;
        ELSIF x =- 16877 THEN
            exp_f := 1;
        ELSIF x =- 16876 THEN
            exp_f := 1;
        ELSIF x =- 16875 THEN
            exp_f := 1;
        ELSIF x =- 16874 THEN
            exp_f := 1;
        ELSIF x =- 16873 THEN
            exp_f := 1;
        ELSIF x =- 16872 THEN
            exp_f := 1;
        ELSIF x =- 16871 THEN
            exp_f := 1;
        ELSIF x =- 16870 THEN
            exp_f := 1;
        ELSIF x =- 16869 THEN
            exp_f := 1;
        ELSIF x =- 16868 THEN
            exp_f := 1;
        ELSIF x =- 16867 THEN
            exp_f := 1;
        ELSIF x =- 16866 THEN
            exp_f := 1;
        ELSIF x =- 16865 THEN
            exp_f := 1;
        ELSIF x =- 16864 THEN
            exp_f := 1;
        ELSIF x =- 16863 THEN
            exp_f := 1;
        ELSIF x =- 16862 THEN
            exp_f := 1;
        ELSIF x =- 16861 THEN
            exp_f := 1;
        ELSIF x =- 16860 THEN
            exp_f := 1;
        ELSIF x =- 16859 THEN
            exp_f := 1;
        ELSIF x =- 16858 THEN
            exp_f := 1;
        ELSIF x =- 16857 THEN
            exp_f := 1;
        ELSIF x =- 16856 THEN
            exp_f := 1;
        ELSIF x =- 16855 THEN
            exp_f := 1;
        ELSIF x =- 16854 THEN
            exp_f := 1;
        ELSIF x =- 16853 THEN
            exp_f := 1;
        ELSIF x =- 16852 THEN
            exp_f := 1;
        ELSIF x =- 16851 THEN
            exp_f := 1;
        ELSIF x =- 16850 THEN
            exp_f := 1;
        ELSIF x =- 16849 THEN
            exp_f := 1;
        ELSIF x =- 16848 THEN
            exp_f := 1;
        ELSIF x =- 16847 THEN
            exp_f := 1;
        ELSIF x =- 16846 THEN
            exp_f := 1;
        ELSIF x =- 16845 THEN
            exp_f := 1;
        ELSIF x =- 16844 THEN
            exp_f := 1;
        ELSIF x =- 16843 THEN
            exp_f := 1;
        ELSIF x =- 16842 THEN
            exp_f := 1;
        ELSIF x =- 16841 THEN
            exp_f := 1;
        ELSIF x =- 16840 THEN
            exp_f := 1;
        ELSIF x =- 16839 THEN
            exp_f := 1;
        ELSIF x =- 16838 THEN
            exp_f := 1;
        ELSIF x =- 16837 THEN
            exp_f := 1;
        ELSIF x =- 16836 THEN
            exp_f := 1;
        ELSIF x =- 16835 THEN
            exp_f := 1;
        ELSIF x =- 16834 THEN
            exp_f := 1;
        ELSIF x =- 16833 THEN
            exp_f := 1;
        ELSIF x =- 16832 THEN
            exp_f := 1;
        ELSIF x =- 16831 THEN
            exp_f := 1;
        ELSIF x =- 16830 THEN
            exp_f := 1;
        ELSIF x =- 16829 THEN
            exp_f := 1;
        ELSIF x =- 16828 THEN
            exp_f := 1;
        ELSIF x =- 16827 THEN
            exp_f := 1;
        ELSIF x =- 16826 THEN
            exp_f := 1;
        ELSIF x =- 16825 THEN
            exp_f := 1;
        ELSIF x =- 16824 THEN
            exp_f := 1;
        ELSIF x =- 16823 THEN
            exp_f := 1;
        ELSIF x =- 16822 THEN
            exp_f := 1;
        ELSIF x =- 16821 THEN
            exp_f := 1;
        ELSIF x =- 16820 THEN
            exp_f := 1;
        ELSIF x =- 16819 THEN
            exp_f := 1;
        ELSIF x =- 16818 THEN
            exp_f := 1;
        ELSIF x =- 16817 THEN
            exp_f := 1;
        ELSIF x =- 16816 THEN
            exp_f := 1;
        ELSIF x =- 16815 THEN
            exp_f := 1;
        ELSIF x =- 16814 THEN
            exp_f := 1;
        ELSIF x =- 16813 THEN
            exp_f := 1;
        ELSIF x =- 16812 THEN
            exp_f := 1;
        ELSIF x =- 16811 THEN
            exp_f := 1;
        ELSIF x =- 16810 THEN
            exp_f := 1;
        ELSIF x =- 16809 THEN
            exp_f := 1;
        ELSIF x =- 16808 THEN
            exp_f := 1;
        ELSIF x =- 16807 THEN
            exp_f := 1;
        ELSIF x =- 16806 THEN
            exp_f := 1;
        ELSIF x =- 16805 THEN
            exp_f := 1;
        ELSIF x =- 16804 THEN
            exp_f := 1;
        ELSIF x =- 16803 THEN
            exp_f := 1;
        ELSIF x =- 16802 THEN
            exp_f := 1;
        ELSIF x =- 16801 THEN
            exp_f := 1;
        ELSIF x =- 16800 THEN
            exp_f := 1;
        ELSIF x =- 16799 THEN
            exp_f := 1;
        ELSIF x =- 16798 THEN
            exp_f := 1;
        ELSIF x =- 16797 THEN
            exp_f := 1;
        ELSIF x =- 16796 THEN
            exp_f := 1;
        ELSIF x =- 16795 THEN
            exp_f := 1;
        ELSIF x =- 16794 THEN
            exp_f := 1;
        ELSIF x =- 16793 THEN
            exp_f := 1;
        ELSIF x =- 16792 THEN
            exp_f := 1;
        ELSIF x =- 16791 THEN
            exp_f := 1;
        ELSIF x =- 16790 THEN
            exp_f := 1;
        ELSIF x =- 16789 THEN
            exp_f := 1;
        ELSIF x =- 16788 THEN
            exp_f := 1;
        ELSIF x =- 16787 THEN
            exp_f := 1;
        ELSIF x =- 16786 THEN
            exp_f := 1;
        ELSIF x =- 16785 THEN
            exp_f := 1;
        ELSIF x =- 16784 THEN
            exp_f := 1;
        ELSIF x =- 16783 THEN
            exp_f := 1;
        ELSIF x =- 16782 THEN
            exp_f := 1;
        ELSIF x =- 16781 THEN
            exp_f := 1;
        ELSIF x =- 16780 THEN
            exp_f := 1;
        ELSIF x =- 16779 THEN
            exp_f := 1;
        ELSIF x =- 16778 THEN
            exp_f := 1;
        ELSIF x =- 16777 THEN
            exp_f := 1;
        ELSIF x =- 16776 THEN
            exp_f := 1;
        ELSIF x =- 16775 THEN
            exp_f := 1;
        ELSIF x =- 16774 THEN
            exp_f := 1;
        ELSIF x =- 16773 THEN
            exp_f := 1;
        ELSIF x =- 16772 THEN
            exp_f := 1;
        ELSIF x =- 16771 THEN
            exp_f := 1;
        ELSIF x =- 16770 THEN
            exp_f := 1;
        ELSIF x =- 16769 THEN
            exp_f := 1;
        ELSIF x =- 16768 THEN
            exp_f := 1;
        ELSIF x =- 16767 THEN
            exp_f := 1;
        ELSIF x =- 16766 THEN
            exp_f := 1;
        ELSIF x =- 16765 THEN
            exp_f := 1;
        ELSIF x =- 16764 THEN
            exp_f := 1;
        ELSIF x =- 16763 THEN
            exp_f := 1;
        ELSIF x =- 16762 THEN
            exp_f := 1;
        ELSIF x =- 16761 THEN
            exp_f := 1;
        ELSIF x =- 16760 THEN
            exp_f := 1;
        ELSIF x =- 16759 THEN
            exp_f := 1;
        ELSIF x =- 16758 THEN
            exp_f := 1;
        ELSIF x =- 16757 THEN
            exp_f := 1;
        ELSIF x =- 16756 THEN
            exp_f := 1;
        ELSIF x =- 16755 THEN
            exp_f := 1;
        ELSIF x =- 16754 THEN
            exp_f := 1;
        ELSIF x =- 16753 THEN
            exp_f := 1;
        ELSIF x =- 16752 THEN
            exp_f := 1;
        ELSIF x =- 16751 THEN
            exp_f := 1;
        ELSIF x =- 16750 THEN
            exp_f := 1;
        ELSIF x =- 16749 THEN
            exp_f := 1;
        ELSIF x =- 16748 THEN
            exp_f := 1;
        ELSIF x =- 16747 THEN
            exp_f := 1;
        ELSIF x =- 16746 THEN
            exp_f := 1;
        ELSIF x =- 16745 THEN
            exp_f := 1;
        ELSIF x =- 16744 THEN
            exp_f := 1;
        ELSIF x =- 16743 THEN
            exp_f := 1;
        ELSIF x =- 16742 THEN
            exp_f := 1;
        ELSIF x =- 16741 THEN
            exp_f := 1;
        ELSIF x =- 16740 THEN
            exp_f := 1;
        ELSIF x =- 16739 THEN
            exp_f := 1;
        ELSIF x =- 16738 THEN
            exp_f := 1;
        ELSIF x =- 16737 THEN
            exp_f := 1;
        ELSIF x =- 16736 THEN
            exp_f := 1;
        ELSIF x =- 16735 THEN
            exp_f := 1;
        ELSIF x =- 16734 THEN
            exp_f := 1;
        ELSIF x =- 16733 THEN
            exp_f := 1;
        ELSIF x =- 16732 THEN
            exp_f := 1;
        ELSIF x =- 16731 THEN
            exp_f := 1;
        ELSIF x =- 16730 THEN
            exp_f := 1;
        ELSIF x =- 16729 THEN
            exp_f := 1;
        ELSIF x =- 16728 THEN
            exp_f := 1;
        ELSIF x =- 16727 THEN
            exp_f := 1;
        ELSIF x =- 16726 THEN
            exp_f := 1;
        ELSIF x =- 16725 THEN
            exp_f := 1;
        ELSIF x =- 16724 THEN
            exp_f := 1;
        ELSIF x =- 16723 THEN
            exp_f := 1;
        ELSIF x =- 16722 THEN
            exp_f := 1;
        ELSIF x =- 16721 THEN
            exp_f := 1;
        ELSIF x =- 16720 THEN
            exp_f := 1;
        ELSIF x =- 16719 THEN
            exp_f := 1;
        ELSIF x =- 16718 THEN
            exp_f := 1;
        ELSIF x =- 16717 THEN
            exp_f := 1;
        ELSIF x =- 16716 THEN
            exp_f := 1;
        ELSIF x =- 16715 THEN
            exp_f := 1;
        ELSIF x =- 16714 THEN
            exp_f := 1;
        ELSIF x =- 16713 THEN
            exp_f := 1;
        ELSIF x =- 16712 THEN
            exp_f := 1;
        ELSIF x =- 16711 THEN
            exp_f := 1;
        ELSIF x =- 16710 THEN
            exp_f := 1;
        ELSIF x =- 16709 THEN
            exp_f := 1;
        ELSIF x =- 16708 THEN
            exp_f := 1;
        ELSIF x =- 16707 THEN
            exp_f := 1;
        ELSIF x =- 16706 THEN
            exp_f := 1;
        ELSIF x =- 16705 THEN
            exp_f := 1;
        ELSIF x =- 16704 THEN
            exp_f := 1;
        ELSIF x =- 16703 THEN
            exp_f := 1;
        ELSIF x =- 16702 THEN
            exp_f := 1;
        ELSIF x =- 16701 THEN
            exp_f := 1;
        ELSIF x =- 16700 THEN
            exp_f := 1;
        ELSIF x =- 16699 THEN
            exp_f := 1;
        ELSIF x =- 16698 THEN
            exp_f := 1;
        ELSIF x =- 16697 THEN
            exp_f := 1;
        ELSIF x =- 16696 THEN
            exp_f := 1;
        ELSIF x =- 16695 THEN
            exp_f := 1;
        ELSIF x =- 16694 THEN
            exp_f := 1;
        ELSIF x =- 16693 THEN
            exp_f := 1;
        ELSIF x =- 16692 THEN
            exp_f := 1;
        ELSIF x =- 16691 THEN
            exp_f := 1;
        ELSIF x =- 16690 THEN
            exp_f := 1;
        ELSIF x =- 16689 THEN
            exp_f := 1;
        ELSIF x =- 16688 THEN
            exp_f := 1;
        ELSIF x =- 16687 THEN
            exp_f := 1;
        ELSIF x =- 16686 THEN
            exp_f := 1;
        ELSIF x =- 16685 THEN
            exp_f := 1;
        ELSIF x =- 16684 THEN
            exp_f := 1;
        ELSIF x =- 16683 THEN
            exp_f := 1;
        ELSIF x =- 16682 THEN
            exp_f := 1;
        ELSIF x =- 16681 THEN
            exp_f := 1;
        ELSIF x =- 16680 THEN
            exp_f := 1;
        ELSIF x =- 16679 THEN
            exp_f := 1;
        ELSIF x =- 16678 THEN
            exp_f := 1;
        ELSIF x =- 16677 THEN
            exp_f := 1;
        ELSIF x =- 16676 THEN
            exp_f := 1;
        ELSIF x =- 16675 THEN
            exp_f := 1;
        ELSIF x =- 16674 THEN
            exp_f := 1;
        ELSIF x =- 16673 THEN
            exp_f := 1;
        ELSIF x =- 16672 THEN
            exp_f := 1;
        ELSIF x =- 16671 THEN
            exp_f := 1;
        ELSIF x =- 16670 THEN
            exp_f := 1;
        ELSIF x =- 16669 THEN
            exp_f := 1;
        ELSIF x =- 16668 THEN
            exp_f := 1;
        ELSIF x =- 16667 THEN
            exp_f := 1;
        ELSIF x =- 16666 THEN
            exp_f := 1;
        ELSIF x =- 16665 THEN
            exp_f := 1;
        ELSIF x =- 16664 THEN
            exp_f := 1;
        ELSIF x =- 16663 THEN
            exp_f := 1;
        ELSIF x =- 16662 THEN
            exp_f := 1;
        ELSIF x =- 16661 THEN
            exp_f := 1;
        ELSIF x =- 16660 THEN
            exp_f := 1;
        ELSIF x =- 16659 THEN
            exp_f := 1;
        ELSIF x =- 16658 THEN
            exp_f := 1;
        ELSIF x =- 16657 THEN
            exp_f := 1;
        ELSIF x =- 16656 THEN
            exp_f := 1;
        ELSIF x =- 16655 THEN
            exp_f := 1;
        ELSIF x =- 16654 THEN
            exp_f := 1;
        ELSIF x =- 16653 THEN
            exp_f := 1;
        ELSIF x =- 16652 THEN
            exp_f := 1;
        ELSIF x =- 16651 THEN
            exp_f := 1;
        ELSIF x =- 16650 THEN
            exp_f := 1;
        ELSIF x =- 16649 THEN
            exp_f := 1;
        ELSIF x =- 16648 THEN
            exp_f := 1;
        ELSIF x =- 16647 THEN
            exp_f := 1;
        ELSIF x =- 16646 THEN
            exp_f := 1;
        ELSIF x =- 16645 THEN
            exp_f := 1;
        ELSIF x =- 16644 THEN
            exp_f := 1;
        ELSIF x =- 16643 THEN
            exp_f := 1;
        ELSIF x =- 16642 THEN
            exp_f := 1;
        ELSIF x =- 16641 THEN
            exp_f := 1;
        ELSIF x =- 16640 THEN
            exp_f := 1;
        ELSIF x =- 16639 THEN
            exp_f := 1;
        ELSIF x =- 16638 THEN
            exp_f := 1;
        ELSIF x =- 16637 THEN
            exp_f := 1;
        ELSIF x =- 16636 THEN
            exp_f := 1;
        ELSIF x =- 16635 THEN
            exp_f := 1;
        ELSIF x =- 16634 THEN
            exp_f := 1;
        ELSIF x =- 16633 THEN
            exp_f := 1;
        ELSIF x =- 16632 THEN
            exp_f := 1;
        ELSIF x =- 16631 THEN
            exp_f := 1;
        ELSIF x =- 16630 THEN
            exp_f := 1;
        ELSIF x =- 16629 THEN
            exp_f := 1;
        ELSIF x =- 16628 THEN
            exp_f := 1;
        ELSIF x =- 16627 THEN
            exp_f := 1;
        ELSIF x =- 16626 THEN
            exp_f := 1;
        ELSIF x =- 16625 THEN
            exp_f := 1;
        ELSIF x =- 16624 THEN
            exp_f := 1;
        ELSIF x =- 16623 THEN
            exp_f := 1;
        ELSIF x =- 16622 THEN
            exp_f := 1;
        ELSIF x =- 16621 THEN
            exp_f := 1;
        ELSIF x =- 16620 THEN
            exp_f := 1;
        ELSIF x =- 16619 THEN
            exp_f := 1;
        ELSIF x =- 16618 THEN
            exp_f := 1;
        ELSIF x =- 16617 THEN
            exp_f := 1;
        ELSIF x =- 16616 THEN
            exp_f := 1;
        ELSIF x =- 16615 THEN
            exp_f := 1;
        ELSIF x =- 16614 THEN
            exp_f := 1;
        ELSIF x =- 16613 THEN
            exp_f := 1;
        ELSIF x =- 16612 THEN
            exp_f := 1;
        ELSIF x =- 16611 THEN
            exp_f := 1;
        ELSIF x =- 16610 THEN
            exp_f := 1;
        ELSIF x =- 16609 THEN
            exp_f := 1;
        ELSIF x =- 16608 THEN
            exp_f := 1;
        ELSIF x =- 16607 THEN
            exp_f := 1;
        ELSIF x =- 16606 THEN
            exp_f := 1;
        ELSIF x =- 16605 THEN
            exp_f := 1;
        ELSIF x =- 16604 THEN
            exp_f := 1;
        ELSIF x =- 16603 THEN
            exp_f := 1;
        ELSIF x =- 16602 THEN
            exp_f := 1;
        ELSIF x =- 16601 THEN
            exp_f := 1;
        ELSIF x =- 16600 THEN
            exp_f := 1;
        ELSIF x =- 16599 THEN
            exp_f := 1;
        ELSIF x =- 16598 THEN
            exp_f := 1;
        ELSIF x =- 16597 THEN
            exp_f := 1;
        ELSIF x =- 16596 THEN
            exp_f := 1;
        ELSIF x =- 16595 THEN
            exp_f := 1;
        ELSIF x =- 16594 THEN
            exp_f := 1;
        ELSIF x =- 16593 THEN
            exp_f := 1;
        ELSIF x =- 16592 THEN
            exp_f := 1;
        ELSIF x =- 16591 THEN
            exp_f := 1;
        ELSIF x =- 16590 THEN
            exp_f := 1;
        ELSIF x =- 16589 THEN
            exp_f := 1;
        ELSIF x =- 16588 THEN
            exp_f := 1;
        ELSIF x =- 16587 THEN
            exp_f := 1;
        ELSIF x =- 16586 THEN
            exp_f := 1;
        ELSIF x =- 16585 THEN
            exp_f := 1;
        ELSIF x =- 16584 THEN
            exp_f := 1;
        ELSIF x =- 16583 THEN
            exp_f := 1;
        ELSIF x =- 16582 THEN
            exp_f := 1;
        ELSIF x =- 16581 THEN
            exp_f := 1;
        ELSIF x =- 16580 THEN
            exp_f := 1;
        ELSIF x =- 16579 THEN
            exp_f := 1;
        ELSIF x =- 16578 THEN
            exp_f := 1;
        ELSIF x =- 16577 THEN
            exp_f := 1;
        ELSIF x =- 16576 THEN
            exp_f := 1;
        ELSIF x =- 16575 THEN
            exp_f := 1;
        ELSIF x =- 16574 THEN
            exp_f := 1;
        ELSIF x =- 16573 THEN
            exp_f := 1;
        ELSIF x =- 16572 THEN
            exp_f := 1;
        ELSIF x =- 16571 THEN
            exp_f := 1;
        ELSIF x =- 16570 THEN
            exp_f := 1;
        ELSIF x =- 16569 THEN
            exp_f := 1;
        ELSIF x =- 16568 THEN
            exp_f := 1;
        ELSIF x =- 16567 THEN
            exp_f := 1;
        ELSIF x =- 16566 THEN
            exp_f := 1;
        ELSIF x =- 16565 THEN
            exp_f := 1;
        ELSIF x =- 16564 THEN
            exp_f := 1;
        ELSIF x =- 16563 THEN
            exp_f := 1;
        ELSIF x =- 16562 THEN
            exp_f := 1;
        ELSIF x =- 16561 THEN
            exp_f := 1;
        ELSIF x =- 16560 THEN
            exp_f := 1;
        ELSIF x =- 16559 THEN
            exp_f := 1;
        ELSIF x =- 16558 THEN
            exp_f := 1;
        ELSIF x =- 16557 THEN
            exp_f := 1;
        ELSIF x =- 16556 THEN
            exp_f := 1;
        ELSIF x =- 16555 THEN
            exp_f := 1;
        ELSIF x =- 16554 THEN
            exp_f := 1;
        ELSIF x =- 16553 THEN
            exp_f := 1;
        ELSIF x =- 16552 THEN
            exp_f := 1;
        ELSIF x =- 16551 THEN
            exp_f := 1;
        ELSIF x =- 16550 THEN
            exp_f := 1;
        ELSIF x =- 16549 THEN
            exp_f := 1;
        ELSIF x =- 16548 THEN
            exp_f := 1;
        ELSIF x =- 16547 THEN
            exp_f := 1;
        ELSIF x =- 16546 THEN
            exp_f := 1;
        ELSIF x =- 16545 THEN
            exp_f := 1;
        ELSIF x =- 16544 THEN
            exp_f := 1;
        ELSIF x =- 16543 THEN
            exp_f := 1;
        ELSIF x =- 16542 THEN
            exp_f := 1;
        ELSIF x =- 16541 THEN
            exp_f := 1;
        ELSIF x =- 16540 THEN
            exp_f := 1;
        ELSIF x =- 16539 THEN
            exp_f := 1;
        ELSIF x =- 16538 THEN
            exp_f := 1;
        ELSIF x =- 16537 THEN
            exp_f := 1;
        ELSIF x =- 16536 THEN
            exp_f := 1;
        ELSIF x =- 16535 THEN
            exp_f := 1;
        ELSIF x =- 16534 THEN
            exp_f := 1;
        ELSIF x =- 16533 THEN
            exp_f := 1;
        ELSIF x =- 16532 THEN
            exp_f := 1;
        ELSIF x =- 16531 THEN
            exp_f := 1;
        ELSIF x =- 16530 THEN
            exp_f := 1;
        ELSIF x =- 16529 THEN
            exp_f := 1;
        ELSIF x =- 16528 THEN
            exp_f := 1;
        ELSIF x =- 16527 THEN
            exp_f := 1;
        ELSIF x =- 16526 THEN
            exp_f := 1;
        ELSIF x =- 16525 THEN
            exp_f := 1;
        ELSIF x =- 16524 THEN
            exp_f := 1;
        ELSIF x =- 16523 THEN
            exp_f := 1;
        ELSIF x =- 16522 THEN
            exp_f := 1;
        ELSIF x =- 16521 THEN
            exp_f := 1;
        ELSIF x =- 16520 THEN
            exp_f := 1;
        ELSIF x =- 16519 THEN
            exp_f := 1;
        ELSIF x =- 16518 THEN
            exp_f := 1;
        ELSIF x =- 16517 THEN
            exp_f := 1;
        ELSIF x =- 16516 THEN
            exp_f := 1;
        ELSIF x =- 16515 THEN
            exp_f := 1;
        ELSIF x =- 16514 THEN
            exp_f := 1;
        ELSIF x =- 16513 THEN
            exp_f := 1;
        ELSIF x =- 16512 THEN
            exp_f := 1;
        ELSIF x =- 16511 THEN
            exp_f := 1;
        ELSIF x =- 16510 THEN
            exp_f := 1;
        ELSIF x =- 16509 THEN
            exp_f := 1;
        ELSIF x =- 16508 THEN
            exp_f := 1;
        ELSIF x =- 16507 THEN
            exp_f := 1;
        ELSIF x =- 16506 THEN
            exp_f := 1;
        ELSIF x =- 16505 THEN
            exp_f := 1;
        ELSIF x =- 16504 THEN
            exp_f := 1;
        ELSIF x =- 16503 THEN
            exp_f := 1;
        ELSIF x =- 16502 THEN
            exp_f := 1;
        ELSIF x =- 16501 THEN
            exp_f := 1;
        ELSIF x =- 16500 THEN
            exp_f := 1;
        ELSIF x =- 16499 THEN
            exp_f := 1;
        ELSIF x =- 16498 THEN
            exp_f := 1;
        ELSIF x =- 16497 THEN
            exp_f := 1;
        ELSIF x =- 16496 THEN
            exp_f := 1;
        ELSIF x =- 16495 THEN
            exp_f := 1;
        ELSIF x =- 16494 THEN
            exp_f := 1;
        ELSIF x =- 16493 THEN
            exp_f := 1;
        ELSIF x =- 16492 THEN
            exp_f := 1;
        ELSIF x =- 16491 THEN
            exp_f := 1;
        ELSIF x =- 16490 THEN
            exp_f := 1;
        ELSIF x =- 16489 THEN
            exp_f := 1;
        ELSIF x =- 16488 THEN
            exp_f := 1;
        ELSIF x =- 16487 THEN
            exp_f := 1;
        ELSIF x =- 16486 THEN
            exp_f := 1;
        ELSIF x =- 16485 THEN
            exp_f := 1;
        ELSIF x =- 16484 THEN
            exp_f := 1;
        ELSIF x =- 16483 THEN
            exp_f := 1;
        ELSIF x =- 16482 THEN
            exp_f := 1;
        ELSIF x =- 16481 THEN
            exp_f := 1;
        ELSIF x =- 16480 THEN
            exp_f := 1;
        ELSIF x =- 16479 THEN
            exp_f := 1;
        ELSIF x =- 16478 THEN
            exp_f := 1;
        ELSIF x =- 16477 THEN
            exp_f := 1;
        ELSIF x =- 16476 THEN
            exp_f := 1;
        ELSIF x =- 16475 THEN
            exp_f := 1;
        ELSIF x =- 16474 THEN
            exp_f := 1;
        ELSIF x =- 16473 THEN
            exp_f := 1;
        ELSIF x =- 16472 THEN
            exp_f := 1;
        ELSIF x =- 16471 THEN
            exp_f := 1;
        ELSIF x =- 16470 THEN
            exp_f := 1;
        ELSIF x =- 16469 THEN
            exp_f := 1;
        ELSIF x =- 16468 THEN
            exp_f := 1;
        ELSIF x =- 16467 THEN
            exp_f := 1;
        ELSIF x =- 16466 THEN
            exp_f := 1;
        ELSIF x =- 16465 THEN
            exp_f := 1;
        ELSIF x =- 16464 THEN
            exp_f := 1;
        ELSIF x =- 16463 THEN
            exp_f := 1;
        ELSIF x =- 16462 THEN
            exp_f := 1;
        ELSIF x =- 16461 THEN
            exp_f := 1;
        ELSIF x =- 16460 THEN
            exp_f := 1;
        ELSIF x =- 16459 THEN
            exp_f := 1;
        ELSIF x =- 16458 THEN
            exp_f := 1;
        ELSIF x =- 16457 THEN
            exp_f := 1;
        ELSIF x =- 16456 THEN
            exp_f := 1;
        ELSIF x =- 16455 THEN
            exp_f := 1;
        ELSIF x =- 16454 THEN
            exp_f := 1;
        ELSIF x =- 16453 THEN
            exp_f := 1;
        ELSIF x =- 16452 THEN
            exp_f := 1;
        ELSIF x =- 16451 THEN
            exp_f := 1;
        ELSIF x =- 16450 THEN
            exp_f := 1;
        ELSIF x =- 16449 THEN
            exp_f := 1;
        ELSIF x =- 16448 THEN
            exp_f := 1;
        ELSIF x =- 16447 THEN
            exp_f := 1;
        ELSIF x =- 16446 THEN
            exp_f := 1;
        ELSIF x =- 16445 THEN
            exp_f := 1;
        ELSIF x =- 16444 THEN
            exp_f := 1;
        ELSIF x =- 16443 THEN
            exp_f := 1;
        ELSIF x =- 16442 THEN
            exp_f := 1;
        ELSIF x =- 16441 THEN
            exp_f := 1;
        ELSIF x =- 16440 THEN
            exp_f := 1;
        ELSIF x =- 16439 THEN
            exp_f := 1;
        ELSIF x =- 16438 THEN
            exp_f := 1;
        ELSIF x =- 16437 THEN
            exp_f := 1;
        ELSIF x =- 16436 THEN
            exp_f := 1;
        ELSIF x =- 16435 THEN
            exp_f := 1;
        ELSIF x =- 16434 THEN
            exp_f := 1;
        ELSIF x =- 16433 THEN
            exp_f := 1;
        ELSIF x =- 16432 THEN
            exp_f := 1;
        ELSIF x =- 16431 THEN
            exp_f := 1;
        ELSIF x =- 16430 THEN
            exp_f := 1;
        ELSIF x =- 16429 THEN
            exp_f := 1;
        ELSIF x =- 16428 THEN
            exp_f := 1;
        ELSIF x =- 16427 THEN
            exp_f := 1;
        ELSIF x =- 16426 THEN
            exp_f := 1;
        ELSIF x =- 16425 THEN
            exp_f := 1;
        ELSIF x =- 16424 THEN
            exp_f := 1;
        ELSIF x =- 16423 THEN
            exp_f := 1;
        ELSIF x =- 16422 THEN
            exp_f := 1;
        ELSIF x =- 16421 THEN
            exp_f := 1;
        ELSIF x =- 16420 THEN
            exp_f := 1;
        ELSIF x =- 16419 THEN
            exp_f := 1;
        ELSIF x =- 16418 THEN
            exp_f := 1;
        ELSIF x =- 16417 THEN
            exp_f := 1;
        ELSIF x =- 16416 THEN
            exp_f := 1;
        ELSIF x =- 16415 THEN
            exp_f := 1;
        ELSIF x =- 16414 THEN
            exp_f := 1;
        ELSIF x =- 16413 THEN
            exp_f := 1;
        ELSIF x =- 16412 THEN
            exp_f := 1;
        ELSIF x =- 16411 THEN
            exp_f := 1;
        ELSIF x =- 16410 THEN
            exp_f := 1;
        ELSIF x =- 16409 THEN
            exp_f := 1;
        ELSIF x =- 16408 THEN
            exp_f := 1;
        ELSIF x =- 16407 THEN
            exp_f := 1;
        ELSIF x =- 16406 THEN
            exp_f := 1;
        ELSIF x =- 16405 THEN
            exp_f := 1;
        ELSIF x =- 16404 THEN
            exp_f := 1;
        ELSIF x =- 16403 THEN
            exp_f := 1;
        ELSIF x =- 16402 THEN
            exp_f := 1;
        ELSIF x =- 16401 THEN
            exp_f := 1;
        ELSIF x =- 16400 THEN
            exp_f := 1;
        ELSIF x =- 16399 THEN
            exp_f := 1;
        ELSIF x =- 16398 THEN
            exp_f := 1;
        ELSIF x =- 16397 THEN
            exp_f := 1;
        ELSIF x =- 16396 THEN
            exp_f := 1;
        ELSIF x =- 16395 THEN
            exp_f := 1;
        ELSIF x =- 16394 THEN
            exp_f := 1;
        ELSIF x =- 16393 THEN
            exp_f := 1;
        ELSIF x =- 16392 THEN
            exp_f := 1;
        ELSIF x =- 16391 THEN
            exp_f := 1;
        ELSIF x =- 16390 THEN
            exp_f := 1;
        ELSIF x =- 16389 THEN
            exp_f := 1;
        ELSIF x =- 16388 THEN
            exp_f := 1;
        ELSIF x =- 16387 THEN
            exp_f := 1;
        ELSIF x =- 16386 THEN
            exp_f := 1;
        ELSIF x =- 16385 THEN
            exp_f := 1;
        ELSIF x =- 16384 THEN
            exp_f := 1;
        ELSIF x =- 16383 THEN
            exp_f := 1;
        ELSIF x =- 16382 THEN
            exp_f := 1;
        ELSIF x =- 16381 THEN
            exp_f := 1;
        ELSIF x =- 16380 THEN
            exp_f := 1;
        ELSIF x =- 16379 THEN
            exp_f := 1;
        ELSIF x =- 16378 THEN
            exp_f := 1;
        ELSIF x =- 16377 THEN
            exp_f := 1;
        ELSIF x =- 16376 THEN
            exp_f := 1;
        ELSIF x =- 16375 THEN
            exp_f := 1;
        ELSIF x =- 16374 THEN
            exp_f := 1;
        ELSIF x =- 16373 THEN
            exp_f := 1;
        ELSIF x =- 16372 THEN
            exp_f := 1;
        ELSIF x =- 16371 THEN
            exp_f := 1;
        ELSIF x =- 16370 THEN
            exp_f := 1;
        ELSIF x =- 16369 THEN
            exp_f := 1;
        ELSIF x =- 16368 THEN
            exp_f := 1;
        ELSIF x =- 16367 THEN
            exp_f := 1;
        ELSIF x =- 16366 THEN
            exp_f := 1;
        ELSIF x =- 16365 THEN
            exp_f := 1;
        ELSIF x =- 16364 THEN
            exp_f := 1;
        ELSIF x =- 16363 THEN
            exp_f := 1;
        ELSIF x =- 16362 THEN
            exp_f := 1;
        ELSIF x =- 16361 THEN
            exp_f := 1;
        ELSIF x =- 16360 THEN
            exp_f := 1;
        ELSIF x =- 16359 THEN
            exp_f := 1;
        ELSIF x =- 16358 THEN
            exp_f := 1;
        ELSIF x =- 16357 THEN
            exp_f := 1;
        ELSIF x =- 16356 THEN
            exp_f := 1;
        ELSIF x =- 16355 THEN
            exp_f := 1;
        ELSIF x =- 16354 THEN
            exp_f := 1;
        ELSIF x =- 16353 THEN
            exp_f := 1;
        ELSIF x =- 16352 THEN
            exp_f := 1;
        ELSIF x =- 16351 THEN
            exp_f := 1;
        ELSIF x =- 16350 THEN
            exp_f := 1;
        ELSIF x =- 16349 THEN
            exp_f := 1;
        ELSIF x =- 16348 THEN
            exp_f := 1;
        ELSIF x =- 16347 THEN
            exp_f := 1;
        ELSIF x =- 16346 THEN
            exp_f := 1;
        ELSIF x =- 16345 THEN
            exp_f := 1;
        ELSIF x =- 16344 THEN
            exp_f := 1;
        ELSIF x =- 16343 THEN
            exp_f := 1;
        ELSIF x =- 16342 THEN
            exp_f := 1;
        ELSIF x =- 16341 THEN
            exp_f := 1;
        ELSIF x =- 16340 THEN
            exp_f := 1;
        ELSIF x =- 16339 THEN
            exp_f := 1;
        ELSIF x =- 16338 THEN
            exp_f := 1;
        ELSIF x =- 16337 THEN
            exp_f := 1;
        ELSIF x =- 16336 THEN
            exp_f := 1;
        ELSIF x =- 16335 THEN
            exp_f := 1;
        ELSIF x =- 16334 THEN
            exp_f := 1;
        ELSIF x =- 16333 THEN
            exp_f := 1;
        ELSIF x =- 16332 THEN
            exp_f := 1;
        ELSIF x =- 16331 THEN
            exp_f := 1;
        ELSIF x =- 16330 THEN
            exp_f := 1;
        ELSIF x =- 16329 THEN
            exp_f := 1;
        ELSIF x =- 16328 THEN
            exp_f := 1;
        ELSIF x =- 16327 THEN
            exp_f := 1;
        ELSIF x =- 16326 THEN
            exp_f := 1;
        ELSIF x =- 16325 THEN
            exp_f := 1;
        ELSIF x =- 16324 THEN
            exp_f := 1;
        ELSIF x =- 16323 THEN
            exp_f := 1;
        ELSIF x =- 16322 THEN
            exp_f := 1;
        ELSIF x =- 16321 THEN
            exp_f := 1;
        ELSIF x =- 16320 THEN
            exp_f := 1;
        ELSIF x =- 16319 THEN
            exp_f := 1;
        ELSIF x =- 16318 THEN
            exp_f := 1;
        ELSIF x =- 16317 THEN
            exp_f := 1;
        ELSIF x =- 16316 THEN
            exp_f := 1;
        ELSIF x =- 16315 THEN
            exp_f := 1;
        ELSIF x =- 16314 THEN
            exp_f := 1;
        ELSIF x =- 16313 THEN
            exp_f := 1;
        ELSIF x =- 16312 THEN
            exp_f := 1;
        ELSIF x =- 16311 THEN
            exp_f := 1;
        ELSIF x =- 16310 THEN
            exp_f := 1;
        ELSIF x =- 16309 THEN
            exp_f := 1;
        ELSIF x =- 16308 THEN
            exp_f := 1;
        ELSIF x =- 16307 THEN
            exp_f := 1;
        ELSIF x =- 16306 THEN
            exp_f := 1;
        ELSIF x =- 16305 THEN
            exp_f := 1;
        ELSIF x =- 16304 THEN
            exp_f := 1;
        ELSIF x =- 16303 THEN
            exp_f := 1;
        ELSIF x =- 16302 THEN
            exp_f := 1;
        ELSIF x =- 16301 THEN
            exp_f := 1;
        ELSIF x =- 16300 THEN
            exp_f := 1;
        ELSIF x =- 16299 THEN
            exp_f := 1;
        ELSIF x =- 16298 THEN
            exp_f := 1;
        ELSIF x =- 16297 THEN
            exp_f := 1;
        ELSIF x =- 16296 THEN
            exp_f := 1;
        ELSIF x =- 16295 THEN
            exp_f := 1;
        ELSIF x =- 16294 THEN
            exp_f := 1;
        ELSIF x =- 16293 THEN
            exp_f := 1;
        ELSIF x =- 16292 THEN
            exp_f := 1;
        ELSIF x =- 16291 THEN
            exp_f := 1;
        ELSIF x =- 16290 THEN
            exp_f := 1;
        ELSIF x =- 16289 THEN
            exp_f := 1;
        ELSIF x =- 16288 THEN
            exp_f := 1;
        ELSIF x =- 16287 THEN
            exp_f := 1;
        ELSIF x =- 16286 THEN
            exp_f := 1;
        ELSIF x =- 16285 THEN
            exp_f := 1;
        ELSIF x =- 16284 THEN
            exp_f := 1;
        ELSIF x =- 16283 THEN
            exp_f := 1;
        ELSIF x =- 16282 THEN
            exp_f := 1;
        ELSIF x =- 16281 THEN
            exp_f := 1;
        ELSIF x =- 16280 THEN
            exp_f := 1;
        ELSIF x =- 16279 THEN
            exp_f := 1;
        ELSIF x =- 16278 THEN
            exp_f := 1;
        ELSIF x =- 16277 THEN
            exp_f := 1;
        ELSIF x =- 16276 THEN
            exp_f := 1;
        ELSIF x =- 16275 THEN
            exp_f := 1;
        ELSIF x =- 16274 THEN
            exp_f := 1;
        ELSIF x =- 16273 THEN
            exp_f := 1;
        ELSIF x =- 16272 THEN
            exp_f := 1;
        ELSIF x =- 16271 THEN
            exp_f := 1;
        ELSIF x =- 16270 THEN
            exp_f := 1;
        ELSIF x =- 16269 THEN
            exp_f := 1;
        ELSIF x =- 16268 THEN
            exp_f := 1;
        ELSIF x =- 16267 THEN
            exp_f := 1;
        ELSIF x =- 16266 THEN
            exp_f := 1;
        ELSIF x =- 16265 THEN
            exp_f := 1;
        ELSIF x =- 16264 THEN
            exp_f := 1;
        ELSIF x =- 16263 THEN
            exp_f := 1;
        ELSIF x =- 16262 THEN
            exp_f := 1;
        ELSIF x =- 16261 THEN
            exp_f := 1;
        ELSIF x =- 16260 THEN
            exp_f := 1;
        ELSIF x =- 16259 THEN
            exp_f := 1;
        ELSIF x =- 16258 THEN
            exp_f := 1;
        ELSIF x =- 16257 THEN
            exp_f := 1;
        ELSIF x =- 16256 THEN
            exp_f := 1;
        ELSIF x =- 16255 THEN
            exp_f := 1;
        ELSIF x =- 16254 THEN
            exp_f := 1;
        ELSIF x =- 16253 THEN
            exp_f := 1;
        ELSIF x =- 16252 THEN
            exp_f := 1;
        ELSIF x =- 16251 THEN
            exp_f := 1;
        ELSIF x =- 16250 THEN
            exp_f := 1;
        ELSIF x =- 16249 THEN
            exp_f := 1;
        ELSIF x =- 16248 THEN
            exp_f := 1;
        ELSIF x =- 16247 THEN
            exp_f := 1;
        ELSIF x =- 16246 THEN
            exp_f := 1;
        ELSIF x =- 16245 THEN
            exp_f := 1;
        ELSIF x =- 16244 THEN
            exp_f := 1;
        ELSIF x =- 16243 THEN
            exp_f := 1;
        ELSIF x =- 16242 THEN
            exp_f := 1;
        ELSIF x =- 16241 THEN
            exp_f := 1;
        ELSIF x =- 16240 THEN
            exp_f := 1;
        ELSIF x =- 16239 THEN
            exp_f := 1;
        ELSIF x =- 16238 THEN
            exp_f := 1;
        ELSIF x =- 16237 THEN
            exp_f := 1;
        ELSIF x =- 16236 THEN
            exp_f := 1;
        ELSIF x =- 16235 THEN
            exp_f := 1;
        ELSIF x =- 16234 THEN
            exp_f := 1;
        ELSIF x =- 16233 THEN
            exp_f := 1;
        ELSIF x =- 16232 THEN
            exp_f := 1;
        ELSIF x =- 16231 THEN
            exp_f := 1;
        ELSIF x =- 16230 THEN
            exp_f := 1;
        ELSIF x =- 16229 THEN
            exp_f := 1;
        ELSIF x =- 16228 THEN
            exp_f := 1;
        ELSIF x =- 16227 THEN
            exp_f := 1;
        ELSIF x =- 16226 THEN
            exp_f := 1;
        ELSIF x =- 16225 THEN
            exp_f := 1;
        ELSIF x =- 16224 THEN
            exp_f := 1;
        ELSIF x =- 16223 THEN
            exp_f := 1;
        ELSIF x =- 16222 THEN
            exp_f := 1;
        ELSIF x =- 16221 THEN
            exp_f := 1;
        ELSIF x =- 16220 THEN
            exp_f := 1;
        ELSIF x =- 16219 THEN
            exp_f := 1;
        ELSIF x =- 16218 THEN
            exp_f := 1;
        ELSIF x =- 16217 THEN
            exp_f := 1;
        ELSIF x =- 16216 THEN
            exp_f := 1;
        ELSIF x =- 16215 THEN
            exp_f := 1;
        ELSIF x =- 16214 THEN
            exp_f := 1;
        ELSIF x =- 16213 THEN
            exp_f := 1;
        ELSIF x =- 16212 THEN
            exp_f := 1;
        ELSIF x =- 16211 THEN
            exp_f := 1;
        ELSIF x =- 16210 THEN
            exp_f := 1;
        ELSIF x =- 16209 THEN
            exp_f := 1;
        ELSIF x =- 16208 THEN
            exp_f := 1;
        ELSIF x =- 16207 THEN
            exp_f := 1;
        ELSIF x =- 16206 THEN
            exp_f := 1;
        ELSIF x =- 16205 THEN
            exp_f := 1;
        ELSIF x =- 16204 THEN
            exp_f := 1;
        ELSIF x =- 16203 THEN
            exp_f := 1;
        ELSIF x =- 16202 THEN
            exp_f := 1;
        ELSIF x =- 16201 THEN
            exp_f := 1;
        ELSIF x =- 16200 THEN
            exp_f := 1;
        ELSIF x =- 16199 THEN
            exp_f := 1;
        ELSIF x =- 16198 THEN
            exp_f := 1;
        ELSIF x =- 16197 THEN
            exp_f := 1;
        ELSIF x =- 16196 THEN
            exp_f := 1;
        ELSIF x =- 16195 THEN
            exp_f := 1;
        ELSIF x =- 16194 THEN
            exp_f := 1;
        ELSIF x =- 16193 THEN
            exp_f := 1;
        ELSIF x =- 16192 THEN
            exp_f := 1;
        ELSIF x =- 16191 THEN
            exp_f := 1;
        ELSIF x =- 16190 THEN
            exp_f := 1;
        ELSIF x =- 16189 THEN
            exp_f := 1;
        ELSIF x =- 16188 THEN
            exp_f := 1;
        ELSIF x =- 16187 THEN
            exp_f := 1;
        ELSIF x =- 16186 THEN
            exp_f := 1;
        ELSIF x =- 16185 THEN
            exp_f := 1;
        ELSIF x =- 16184 THEN
            exp_f := 1;
        ELSIF x =- 16183 THEN
            exp_f := 1;
        ELSIF x =- 16182 THEN
            exp_f := 1;
        ELSIF x =- 16181 THEN
            exp_f := 1;
        ELSIF x =- 16180 THEN
            exp_f := 1;
        ELSIF x =- 16179 THEN
            exp_f := 1;
        ELSIF x =- 16178 THEN
            exp_f := 1;
        ELSIF x =- 16177 THEN
            exp_f := 1;
        ELSIF x =- 16176 THEN
            exp_f := 1;
        ELSIF x =- 16175 THEN
            exp_f := 1;
        ELSIF x =- 16174 THEN
            exp_f := 1;
        ELSIF x =- 16173 THEN
            exp_f := 1;
        ELSIF x =- 16172 THEN
            exp_f := 1;
        ELSIF x =- 16171 THEN
            exp_f := 1;
        ELSIF x =- 16170 THEN
            exp_f := 1;
        ELSIF x =- 16169 THEN
            exp_f := 1;
        ELSIF x =- 16168 THEN
            exp_f := 1;
        ELSIF x =- 16167 THEN
            exp_f := 1;
        ELSIF x =- 16166 THEN
            exp_f := 1;
        ELSIF x =- 16165 THEN
            exp_f := 1;
        ELSIF x =- 16164 THEN
            exp_f := 1;
        ELSIF x =- 16163 THEN
            exp_f := 1;
        ELSIF x =- 16162 THEN
            exp_f := 1;
        ELSIF x =- 16161 THEN
            exp_f := 1;
        ELSIF x =- 16160 THEN
            exp_f := 1;
        ELSIF x =- 16159 THEN
            exp_f := 1;
        ELSIF x =- 16158 THEN
            exp_f := 1;
        ELSIF x =- 16157 THEN
            exp_f := 1;
        ELSIF x =- 16156 THEN
            exp_f := 1;
        ELSIF x =- 16155 THEN
            exp_f := 1;
        ELSIF x =- 16154 THEN
            exp_f := 1;
        ELSIF x =- 16153 THEN
            exp_f := 1;
        ELSIF x =- 16152 THEN
            exp_f := 1;
        ELSIF x =- 16151 THEN
            exp_f := 1;
        ELSIF x =- 16150 THEN
            exp_f := 1;
        ELSIF x =- 16149 THEN
            exp_f := 1;
        ELSIF x =- 16148 THEN
            exp_f := 1;
        ELSIF x =- 16147 THEN
            exp_f := 1;
        ELSIF x =- 16146 THEN
            exp_f := 1;
        ELSIF x =- 16145 THEN
            exp_f := 1;
        ELSIF x =- 16144 THEN
            exp_f := 1;
        ELSIF x =- 16143 THEN
            exp_f := 1;
        ELSIF x =- 16142 THEN
            exp_f := 1;
        ELSIF x =- 16141 THEN
            exp_f := 1;
        ELSIF x =- 16140 THEN
            exp_f := 1;
        ELSIF x =- 16139 THEN
            exp_f := 1;
        ELSIF x =- 16138 THEN
            exp_f := 1;
        ELSIF x =- 16137 THEN
            exp_f := 1;
        ELSIF x =- 16136 THEN
            exp_f := 1;
        ELSIF x =- 16135 THEN
            exp_f := 1;
        ELSIF x =- 16134 THEN
            exp_f := 1;
        ELSIF x =- 16133 THEN
            exp_f := 1;
        ELSIF x =- 16132 THEN
            exp_f := 1;
        ELSIF x =- 16131 THEN
            exp_f := 1;
        ELSIF x =- 16130 THEN
            exp_f := 1;
        ELSIF x =- 16129 THEN
            exp_f := 1;
        ELSIF x =- 16128 THEN
            exp_f := 1;
        ELSIF x =- 16127 THEN
            exp_f := 1;
        ELSIF x =- 16126 THEN
            exp_f := 1;
        ELSIF x =- 16125 THEN
            exp_f := 1;
        ELSIF x =- 16124 THEN
            exp_f := 1;
        ELSIF x =- 16123 THEN
            exp_f := 1;
        ELSIF x =- 16122 THEN
            exp_f := 1;
        ELSIF x =- 16121 THEN
            exp_f := 1;
        ELSIF x =- 16120 THEN
            exp_f := 1;
        ELSIF x =- 16119 THEN
            exp_f := 1;
        ELSIF x =- 16118 THEN
            exp_f := 1;
        ELSIF x =- 16117 THEN
            exp_f := 1;
        ELSIF x =- 16116 THEN
            exp_f := 1;
        ELSIF x =- 16115 THEN
            exp_f := 1;
        ELSIF x =- 16114 THEN
            exp_f := 1;
        ELSIF x =- 16113 THEN
            exp_f := 1;
        ELSIF x =- 16112 THEN
            exp_f := 1;
        ELSIF x =- 16111 THEN
            exp_f := 1;
        ELSIF x =- 16110 THEN
            exp_f := 1;
        ELSIF x =- 16109 THEN
            exp_f := 1;
        ELSIF x =- 16108 THEN
            exp_f := 1;
        ELSIF x =- 16107 THEN
            exp_f := 1;
        ELSIF x =- 16106 THEN
            exp_f := 1;
        ELSIF x =- 16105 THEN
            exp_f := 1;
        ELSIF x =- 16104 THEN
            exp_f := 1;
        ELSIF x =- 16103 THEN
            exp_f := 1;
        ELSIF x =- 16102 THEN
            exp_f := 1;
        ELSIF x =- 16101 THEN
            exp_f := 1;
        ELSIF x =- 16100 THEN
            exp_f := 1;
        ELSIF x =- 16099 THEN
            exp_f := 1;
        ELSIF x =- 16098 THEN
            exp_f := 1;
        ELSIF x =- 16097 THEN
            exp_f := 1;
        ELSIF x =- 16096 THEN
            exp_f := 1;
        ELSIF x =- 16095 THEN
            exp_f := 1;
        ELSIF x =- 16094 THEN
            exp_f := 1;
        ELSIF x =- 16093 THEN
            exp_f := 1;
        ELSIF x =- 16092 THEN
            exp_f := 1;
        ELSIF x =- 16091 THEN
            exp_f := 1;
        ELSIF x =- 16090 THEN
            exp_f := 1;
        ELSIF x =- 16089 THEN
            exp_f := 1;
        ELSIF x =- 16088 THEN
            exp_f := 1;
        ELSIF x =- 16087 THEN
            exp_f := 1;
        ELSIF x =- 16086 THEN
            exp_f := 1;
        ELSIF x =- 16085 THEN
            exp_f := 1;
        ELSIF x =- 16084 THEN
            exp_f := 1;
        ELSIF x =- 16083 THEN
            exp_f := 1;
        ELSIF x =- 16082 THEN
            exp_f := 1;
        ELSIF x =- 16081 THEN
            exp_f := 1;
        ELSIF x =- 16080 THEN
            exp_f := 1;
        ELSIF x =- 16079 THEN
            exp_f := 1;
        ELSIF x =- 16078 THEN
            exp_f := 1;
        ELSIF x =- 16077 THEN
            exp_f := 1;
        ELSIF x =- 16076 THEN
            exp_f := 1;
        ELSIF x =- 16075 THEN
            exp_f := 1;
        ELSIF x =- 16074 THEN
            exp_f := 1;
        ELSIF x =- 16073 THEN
            exp_f := 1;
        ELSIF x =- 16072 THEN
            exp_f := 1;
        ELSIF x =- 16071 THEN
            exp_f := 1;
        ELSIF x =- 16070 THEN
            exp_f := 1;
        ELSIF x =- 16069 THEN
            exp_f := 1;
        ELSIF x =- 16068 THEN
            exp_f := 1;
        ELSIF x =- 16067 THEN
            exp_f := 1;
        ELSIF x =- 16066 THEN
            exp_f := 1;
        ELSIF x =- 16065 THEN
            exp_f := 1;
        ELSIF x =- 16064 THEN
            exp_f := 1;
        ELSIF x =- 16063 THEN
            exp_f := 1;
        ELSIF x =- 16062 THEN
            exp_f := 1;
        ELSIF x =- 16061 THEN
            exp_f := 1;
        ELSIF x =- 16060 THEN
            exp_f := 1;
        ELSIF x =- 16059 THEN
            exp_f := 1;
        ELSIF x =- 16058 THEN
            exp_f := 1;
        ELSIF x =- 16057 THEN
            exp_f := 1;
        ELSIF x =- 16056 THEN
            exp_f := 1;
        ELSIF x =- 16055 THEN
            exp_f := 1;
        ELSIF x =- 16054 THEN
            exp_f := 1;
        ELSIF x =- 16053 THEN
            exp_f := 1;
        ELSIF x =- 16052 THEN
            exp_f := 1;
        ELSIF x =- 16051 THEN
            exp_f := 1;
        ELSIF x =- 16050 THEN
            exp_f := 1;
        ELSIF x =- 16049 THEN
            exp_f := 1;
        ELSIF x =- 16048 THEN
            exp_f := 1;
        ELSIF x =- 16047 THEN
            exp_f := 1;
        ELSIF x =- 16046 THEN
            exp_f := 1;
        ELSIF x =- 16045 THEN
            exp_f := 1;
        ELSIF x =- 16044 THEN
            exp_f := 1;
        ELSIF x =- 16043 THEN
            exp_f := 1;
        ELSIF x =- 16042 THEN
            exp_f := 1;
        ELSIF x =- 16041 THEN
            exp_f := 1;
        ELSIF x =- 16040 THEN
            exp_f := 1;
        ELSIF x =- 16039 THEN
            exp_f := 1;
        ELSIF x =- 16038 THEN
            exp_f := 1;
        ELSIF x =- 16037 THEN
            exp_f := 1;
        ELSIF x =- 16036 THEN
            exp_f := 1;
        ELSIF x =- 16035 THEN
            exp_f := 1;
        ELSIF x =- 16034 THEN
            exp_f := 1;
        ELSIF x =- 16033 THEN
            exp_f := 1;
        ELSIF x =- 16032 THEN
            exp_f := 1;
        ELSIF x =- 16031 THEN
            exp_f := 1;
        ELSIF x =- 16030 THEN
            exp_f := 1;
        ELSIF x =- 16029 THEN
            exp_f := 1;
        ELSIF x =- 16028 THEN
            exp_f := 1;
        ELSIF x =- 16027 THEN
            exp_f := 1;
        ELSIF x =- 16026 THEN
            exp_f := 1;
        ELSIF x =- 16025 THEN
            exp_f := 1;
        ELSIF x =- 16024 THEN
            exp_f := 1;
        ELSIF x =- 16023 THEN
            exp_f := 1;
        ELSIF x =- 16022 THEN
            exp_f := 1;
        ELSIF x =- 16021 THEN
            exp_f := 1;
        ELSIF x =- 16020 THEN
            exp_f := 1;
        ELSIF x =- 16019 THEN
            exp_f := 1;
        ELSIF x =- 16018 THEN
            exp_f := 1;
        ELSIF x =- 16017 THEN
            exp_f := 1;
        ELSIF x =- 16016 THEN
            exp_f := 1;
        ELSIF x =- 16015 THEN
            exp_f := 1;
        ELSIF x =- 16014 THEN
            exp_f := 1;
        ELSIF x =- 16013 THEN
            exp_f := 1;
        ELSIF x =- 16012 THEN
            exp_f := 1;
        ELSIF x =- 16011 THEN
            exp_f := 1;
        ELSIF x =- 16010 THEN
            exp_f := 1;
        ELSIF x =- 16009 THEN
            exp_f := 1;
        ELSIF x =- 16008 THEN
            exp_f := 1;
        ELSIF x =- 16007 THEN
            exp_f := 1;
        ELSIF x =- 16006 THEN
            exp_f := 1;
        ELSIF x =- 16005 THEN
            exp_f := 1;
        ELSIF x =- 16004 THEN
            exp_f := 1;
        ELSIF x =- 16003 THEN
            exp_f := 1;
        ELSIF x =- 16002 THEN
            exp_f := 1;
        ELSIF x =- 16001 THEN
            exp_f := 1;
        ELSIF x =- 16000 THEN
            exp_f := 1;
        ELSIF x =- 15999 THEN
            exp_f := 1;
        ELSIF x =- 15998 THEN
            exp_f := 1;
        ELSIF x =- 15997 THEN
            exp_f := 1;
        ELSIF x =- 15996 THEN
            exp_f := 1;
        ELSIF x =- 15995 THEN
            exp_f := 1;
        ELSIF x =- 15994 THEN
            exp_f := 1;
        ELSIF x =- 15993 THEN
            exp_f := 1;
        ELSIF x =- 15992 THEN
            exp_f := 1;
        ELSIF x =- 15991 THEN
            exp_f := 1;
        ELSIF x =- 15990 THEN
            exp_f := 1;
        ELSIF x =- 15989 THEN
            exp_f := 1;
        ELSIF x =- 15988 THEN
            exp_f := 1;
        ELSIF x =- 15987 THEN
            exp_f := 1;
        ELSIF x =- 15986 THEN
            exp_f := 1;
        ELSIF x =- 15985 THEN
            exp_f := 1;
        ELSIF x =- 15984 THEN
            exp_f := 1;
        ELSIF x =- 15983 THEN
            exp_f := 1;
        ELSIF x =- 15982 THEN
            exp_f := 1;
        ELSIF x =- 15981 THEN
            exp_f := 1;
        ELSIF x =- 15980 THEN
            exp_f := 1;
        ELSIF x =- 15979 THEN
            exp_f := 1;
        ELSIF x =- 15978 THEN
            exp_f := 1;
        ELSIF x =- 15977 THEN
            exp_f := 1;
        ELSIF x =- 15976 THEN
            exp_f := 1;
        ELSIF x =- 15975 THEN
            exp_f := 1;
        ELSIF x =- 15974 THEN
            exp_f := 1;
        ELSIF x =- 15973 THEN
            exp_f := 1;
        ELSIF x =- 15972 THEN
            exp_f := 1;
        ELSIF x =- 15971 THEN
            exp_f := 1;
        ELSIF x =- 15970 THEN
            exp_f := 1;
        ELSIF x =- 15969 THEN
            exp_f := 1;
        ELSIF x =- 15968 THEN
            exp_f := 1;
        ELSIF x =- 15967 THEN
            exp_f := 1;
        ELSIF x =- 15966 THEN
            exp_f := 1;
        ELSIF x =- 15965 THEN
            exp_f := 1;
        ELSIF x =- 15964 THEN
            exp_f := 1;
        ELSIF x =- 15963 THEN
            exp_f := 1;
        ELSIF x =- 15962 THEN
            exp_f := 1;
        ELSIF x =- 15961 THEN
            exp_f := 1;
        ELSIF x =- 15960 THEN
            exp_f := 1;
        ELSIF x =- 15959 THEN
            exp_f := 1;
        ELSIF x =- 15958 THEN
            exp_f := 1;
        ELSIF x =- 15957 THEN
            exp_f := 1;
        ELSIF x =- 15956 THEN
            exp_f := 1;
        ELSIF x =- 15955 THEN
            exp_f := 1;
        ELSIF x =- 15954 THEN
            exp_f := 1;
        ELSIF x =- 15953 THEN
            exp_f := 1;
        ELSIF x =- 15952 THEN
            exp_f := 1;
        ELSIF x =- 15951 THEN
            exp_f := 1;
        ELSIF x =- 15950 THEN
            exp_f := 1;
        ELSIF x =- 15949 THEN
            exp_f := 1;
        ELSIF x =- 15948 THEN
            exp_f := 1;
        ELSIF x =- 15947 THEN
            exp_f := 1;
        ELSIF x =- 15946 THEN
            exp_f := 1;
        ELSIF x =- 15945 THEN
            exp_f := 1;
        ELSIF x =- 15944 THEN
            exp_f := 1;
        ELSIF x =- 15943 THEN
            exp_f := 1;
        ELSIF x =- 15942 THEN
            exp_f := 1;
        ELSIF x =- 15941 THEN
            exp_f := 1;
        ELSIF x =- 15940 THEN
            exp_f := 1;
        ELSIF x =- 15939 THEN
            exp_f := 1;
        ELSIF x =- 15938 THEN
            exp_f := 1;
        ELSIF x =- 15937 THEN
            exp_f := 1;
        ELSIF x =- 15936 THEN
            exp_f := 1;
        ELSIF x =- 15935 THEN
            exp_f := 1;
        ELSIF x =- 15934 THEN
            exp_f := 1;
        ELSIF x =- 15933 THEN
            exp_f := 1;
        ELSIF x =- 15932 THEN
            exp_f := 1;
        ELSIF x =- 15931 THEN
            exp_f := 1;
        ELSIF x =- 15930 THEN
            exp_f := 1;
        ELSIF x =- 15929 THEN
            exp_f := 1;
        ELSIF x =- 15928 THEN
            exp_f := 1;
        ELSIF x =- 15927 THEN
            exp_f := 1;
        ELSIF x =- 15926 THEN
            exp_f := 1;
        ELSIF x =- 15925 THEN
            exp_f := 1;
        ELSIF x =- 15924 THEN
            exp_f := 1;
        ELSIF x =- 15923 THEN
            exp_f := 1;
        ELSIF x =- 15922 THEN
            exp_f := 1;
        ELSIF x =- 15921 THEN
            exp_f := 1;
        ELSIF x =- 15920 THEN
            exp_f := 1;
        ELSIF x =- 15919 THEN
            exp_f := 1;
        ELSIF x =- 15918 THEN
            exp_f := 1;
        ELSIF x =- 15917 THEN
            exp_f := 1;
        ELSIF x =- 15916 THEN
            exp_f := 1;
        ELSIF x =- 15915 THEN
            exp_f := 1;
        ELSIF x =- 15914 THEN
            exp_f := 1;
        ELSIF x =- 15913 THEN
            exp_f := 1;
        ELSIF x =- 15912 THEN
            exp_f := 1;
        ELSIF x =- 15911 THEN
            exp_f := 1;
        ELSIF x =- 15910 THEN
            exp_f := 1;
        ELSIF x =- 15909 THEN
            exp_f := 1;
        ELSIF x =- 15908 THEN
            exp_f := 1;
        ELSIF x =- 15907 THEN
            exp_f := 1;
        ELSIF x =- 15906 THEN
            exp_f := 1;
        ELSIF x =- 15905 THEN
            exp_f := 1;
        ELSIF x =- 15904 THEN
            exp_f := 1;
        ELSIF x =- 15903 THEN
            exp_f := 1;
        ELSIF x =- 15902 THEN
            exp_f := 1;
        ELSIF x =- 15901 THEN
            exp_f := 1;
        ELSIF x =- 15900 THEN
            exp_f := 1;
        ELSIF x =- 15899 THEN
            exp_f := 1;
        ELSIF x =- 15898 THEN
            exp_f := 1;
        ELSIF x =- 15897 THEN
            exp_f := 1;
        ELSIF x =- 15896 THEN
            exp_f := 1;
        ELSIF x =- 15895 THEN
            exp_f := 1;
        ELSIF x =- 15894 THEN
            exp_f := 1;
        ELSIF x =- 15893 THEN
            exp_f := 1;
        ELSIF x =- 15892 THEN
            exp_f := 1;
        ELSIF x =- 15891 THEN
            exp_f := 1;
        ELSIF x =- 15890 THEN
            exp_f := 1;
        ELSIF x =- 15889 THEN
            exp_f := 1;
        ELSIF x =- 15888 THEN
            exp_f := 1;
        ELSIF x =- 15887 THEN
            exp_f := 1;
        ELSIF x =- 15886 THEN
            exp_f := 1;
        ELSIF x =- 15885 THEN
            exp_f := 1;
        ELSIF x =- 15884 THEN
            exp_f := 1;
        ELSIF x =- 15883 THEN
            exp_f := 1;
        ELSIF x =- 15882 THEN
            exp_f := 1;
        ELSIF x =- 15881 THEN
            exp_f := 1;
        ELSIF x =- 15880 THEN
            exp_f := 1;
        ELSIF x =- 15879 THEN
            exp_f := 1;
        ELSIF x =- 15878 THEN
            exp_f := 1;
        ELSIF x =- 15877 THEN
            exp_f := 1;
        ELSIF x =- 15876 THEN
            exp_f := 1;
        ELSIF x =- 15875 THEN
            exp_f := 1;
        ELSIF x =- 15874 THEN
            exp_f := 1;
        ELSIF x =- 15873 THEN
            exp_f := 1;
        ELSIF x =- 15872 THEN
            exp_f := 1;
        ELSIF x =- 15871 THEN
            exp_f := 1;
        ELSIF x =- 15870 THEN
            exp_f := 1;
        ELSIF x =- 15869 THEN
            exp_f := 1;
        ELSIF x =- 15868 THEN
            exp_f := 1;
        ELSIF x =- 15867 THEN
            exp_f := 1;
        ELSIF x =- 15866 THEN
            exp_f := 1;
        ELSIF x =- 15865 THEN
            exp_f := 1;
        ELSIF x =- 15864 THEN
            exp_f := 1;
        ELSIF x =- 15863 THEN
            exp_f := 1;
        ELSIF x =- 15862 THEN
            exp_f := 1;
        ELSIF x =- 15861 THEN
            exp_f := 1;
        ELSIF x =- 15860 THEN
            exp_f := 1;
        ELSIF x =- 15859 THEN
            exp_f := 1;
        ELSIF x =- 15858 THEN
            exp_f := 1;
        ELSIF x =- 15857 THEN
            exp_f := 1;
        ELSIF x =- 15856 THEN
            exp_f := 1;
        ELSIF x =- 15855 THEN
            exp_f := 1;
        ELSIF x =- 15854 THEN
            exp_f := 1;
        ELSIF x =- 15853 THEN
            exp_f := 1;
        ELSIF x =- 15852 THEN
            exp_f := 1;
        ELSIF x =- 15851 THEN
            exp_f := 1;
        ELSIF x =- 15850 THEN
            exp_f := 1;
        ELSIF x =- 15849 THEN
            exp_f := 1;
        ELSIF x =- 15848 THEN
            exp_f := 1;
        ELSIF x =- 15847 THEN
            exp_f := 1;
        ELSIF x =- 15846 THEN
            exp_f := 1;
        ELSIF x =- 15845 THEN
            exp_f := 1;
        ELSIF x =- 15844 THEN
            exp_f := 1;
        ELSIF x =- 15843 THEN
            exp_f := 1;
        ELSIF x =- 15842 THEN
            exp_f := 1;
        ELSIF x =- 15841 THEN
            exp_f := 1;
        ELSIF x =- 15840 THEN
            exp_f := 1;
        ELSIF x =- 15839 THEN
            exp_f := 1;
        ELSIF x =- 15838 THEN
            exp_f := 1;
        ELSIF x =- 15837 THEN
            exp_f := 1;
        ELSIF x =- 15836 THEN
            exp_f := 1;
        ELSIF x =- 15835 THEN
            exp_f := 1;
        ELSIF x =- 15834 THEN
            exp_f := 1;
        ELSIF x =- 15833 THEN
            exp_f := 1;
        ELSIF x =- 15832 THEN
            exp_f := 1;
        ELSIF x =- 15831 THEN
            exp_f := 1;
        ELSIF x =- 15830 THEN
            exp_f := 1;
        ELSIF x =- 15829 THEN
            exp_f := 1;
        ELSIF x =- 15828 THEN
            exp_f := 1;
        ELSIF x =- 15827 THEN
            exp_f := 1;
        ELSIF x =- 15826 THEN
            exp_f := 1;
        ELSIF x =- 15825 THEN
            exp_f := 1;
        ELSIF x =- 15824 THEN
            exp_f := 1;
        ELSIF x =- 15823 THEN
            exp_f := 1;
        ELSIF x =- 15822 THEN
            exp_f := 1;
        ELSIF x =- 15821 THEN
            exp_f := 1;
        ELSIF x =- 15820 THEN
            exp_f := 1;
        ELSIF x =- 15819 THEN
            exp_f := 1;
        ELSIF x =- 15818 THEN
            exp_f := 1;
        ELSIF x =- 15817 THEN
            exp_f := 1;
        ELSIF x =- 15816 THEN
            exp_f := 1;
        ELSIF x =- 15815 THEN
            exp_f := 1;
        ELSIF x =- 15814 THEN
            exp_f := 1;
        ELSIF x =- 15813 THEN
            exp_f := 1;
        ELSIF x =- 15812 THEN
            exp_f := 1;
        ELSIF x =- 15811 THEN
            exp_f := 1;
        ELSIF x =- 15810 THEN
            exp_f := 1;
        ELSIF x =- 15809 THEN
            exp_f := 1;
        ELSIF x =- 15808 THEN
            exp_f := 1;
        ELSIF x =- 15807 THEN
            exp_f := 1;
        ELSIF x =- 15806 THEN
            exp_f := 1;
        ELSIF x =- 15805 THEN
            exp_f := 1;
        ELSIF x =- 15804 THEN
            exp_f := 1;
        ELSIF x =- 15803 THEN
            exp_f := 1;
        ELSIF x =- 15802 THEN
            exp_f := 1;
        ELSIF x =- 15801 THEN
            exp_f := 1;
        ELSIF x =- 15800 THEN
            exp_f := 1;
        ELSIF x =- 15799 THEN
            exp_f := 1;
        ELSIF x =- 15798 THEN
            exp_f := 1;
        ELSIF x =- 15797 THEN
            exp_f := 1;
        ELSIF x =- 15796 THEN
            exp_f := 1;
        ELSIF x =- 15795 THEN
            exp_f := 1;
        ELSIF x =- 15794 THEN
            exp_f := 1;
        ELSIF x =- 15793 THEN
            exp_f := 1;
        ELSIF x =- 15792 THEN
            exp_f := 1;
        ELSIF x =- 15791 THEN
            exp_f := 1;
        ELSIF x =- 15790 THEN
            exp_f := 1;
        ELSIF x =- 15789 THEN
            exp_f := 1;
        ELSIF x =- 15788 THEN
            exp_f := 1;
        ELSIF x =- 15787 THEN
            exp_f := 1;
        ELSIF x =- 15786 THEN
            exp_f := 1;
        ELSIF x =- 15785 THEN
            exp_f := 1;
        ELSIF x =- 15784 THEN
            exp_f := 1;
        ELSIF x =- 15783 THEN
            exp_f := 1;
        ELSIF x =- 15782 THEN
            exp_f := 1;
        ELSIF x =- 15781 THEN
            exp_f := 1;
        ELSIF x =- 15780 THEN
            exp_f := 1;
        ELSIF x =- 15779 THEN
            exp_f := 1;
        ELSIF x =- 15778 THEN
            exp_f := 1;
        ELSIF x =- 15777 THEN
            exp_f := 1;
        ELSIF x =- 15776 THEN
            exp_f := 1;
        ELSIF x =- 15775 THEN
            exp_f := 1;
        ELSIF x =- 15774 THEN
            exp_f := 1;
        ELSIF x =- 15773 THEN
            exp_f := 1;
        ELSIF x =- 15772 THEN
            exp_f := 1;
        ELSIF x =- 15771 THEN
            exp_f := 1;
        ELSIF x =- 15770 THEN
            exp_f := 1;
        ELSIF x =- 15769 THEN
            exp_f := 1;
        ELSIF x =- 15768 THEN
            exp_f := 1;
        ELSIF x =- 15767 THEN
            exp_f := 1;
        ELSIF x =- 15766 THEN
            exp_f := 1;
        ELSIF x =- 15765 THEN
            exp_f := 1;
        ELSIF x =- 15764 THEN
            exp_f := 1;
        ELSIF x =- 15763 THEN
            exp_f := 1;
        ELSIF x =- 15762 THEN
            exp_f := 1;
        ELSIF x =- 15761 THEN
            exp_f := 1;
        ELSIF x =- 15760 THEN
            exp_f := 1;
        ELSIF x =- 15759 THEN
            exp_f := 1;
        ELSIF x =- 15758 THEN
            exp_f := 1;
        ELSIF x =- 15757 THEN
            exp_f := 1;
        ELSIF x =- 15756 THEN
            exp_f := 1;
        ELSIF x =- 15755 THEN
            exp_f := 1;
        ELSIF x =- 15754 THEN
            exp_f := 1;
        ELSIF x =- 15753 THEN
            exp_f := 1;
        ELSIF x =- 15752 THEN
            exp_f := 1;
        ELSIF x =- 15751 THEN
            exp_f := 1;
        ELSIF x =- 15750 THEN
            exp_f := 1;
        ELSIF x =- 15749 THEN
            exp_f := 1;
        ELSIF x =- 15748 THEN
            exp_f := 1;
        ELSIF x =- 15747 THEN
            exp_f := 1;
        ELSIF x =- 15746 THEN
            exp_f := 1;
        ELSIF x =- 15745 THEN
            exp_f := 1;
        ELSIF x =- 15744 THEN
            exp_f := 1;
        ELSIF x =- 15743 THEN
            exp_f := 1;
        ELSIF x =- 15742 THEN
            exp_f := 1;
        ELSIF x =- 15741 THEN
            exp_f := 1;
        ELSIF x =- 15740 THEN
            exp_f := 1;
        ELSIF x =- 15739 THEN
            exp_f := 1;
        ELSIF x =- 15738 THEN
            exp_f := 1;
        ELSIF x =- 15737 THEN
            exp_f := 1;
        ELSIF x =- 15736 THEN
            exp_f := 1;
        ELSIF x =- 15735 THEN
            exp_f := 1;
        ELSIF x =- 15734 THEN
            exp_f := 1;
        ELSIF x =- 15733 THEN
            exp_f := 1;
        ELSIF x =- 15732 THEN
            exp_f := 1;
        ELSIF x =- 15731 THEN
            exp_f := 1;
        ELSIF x =- 15730 THEN
            exp_f := 1;
        ELSIF x =- 15729 THEN
            exp_f := 1;
        ELSIF x =- 15728 THEN
            exp_f := 1;
        ELSIF x =- 15727 THEN
            exp_f := 1;
        ELSIF x =- 15726 THEN
            exp_f := 1;
        ELSIF x =- 15725 THEN
            exp_f := 1;
        ELSIF x =- 15724 THEN
            exp_f := 1;
        ELSIF x =- 15723 THEN
            exp_f := 1;
        ELSIF x =- 15722 THEN
            exp_f := 1;
        ELSIF x =- 15721 THEN
            exp_f := 1;
        ELSIF x =- 15720 THEN
            exp_f := 1;
        ELSIF x =- 15719 THEN
            exp_f := 1;
        ELSIF x =- 15718 THEN
            exp_f := 1;
        ELSIF x =- 15717 THEN
            exp_f := 1;
        ELSIF x =- 15716 THEN
            exp_f := 1;
        ELSIF x =- 15715 THEN
            exp_f := 1;
        ELSIF x =- 15714 THEN
            exp_f := 1;
        ELSIF x =- 15713 THEN
            exp_f := 1;
        ELSIF x =- 15712 THEN
            exp_f := 1;
        ELSIF x =- 15711 THEN
            exp_f := 1;
        ELSIF x =- 15710 THEN
            exp_f := 1;
        ELSIF x =- 15709 THEN
            exp_f := 1;
        ELSIF x =- 15708 THEN
            exp_f := 1;
        ELSIF x =- 15707 THEN
            exp_f := 1;
        ELSIF x =- 15706 THEN
            exp_f := 1;
        ELSIF x =- 15705 THEN
            exp_f := 1;
        ELSIF x =- 15704 THEN
            exp_f := 1;
        ELSIF x =- 15703 THEN
            exp_f := 1;
        ELSIF x =- 15702 THEN
            exp_f := 1;
        ELSIF x =- 15701 THEN
            exp_f := 1;
        ELSIF x =- 15700 THEN
            exp_f := 1;
        ELSIF x =- 15699 THEN
            exp_f := 1;
        ELSIF x =- 15698 THEN
            exp_f := 1;
        ELSIF x =- 15697 THEN
            exp_f := 1;
        ELSIF x =- 15696 THEN
            exp_f := 1;
        ELSIF x =- 15695 THEN
            exp_f := 1;
        ELSIF x =- 15694 THEN
            exp_f := 1;
        ELSIF x =- 15693 THEN
            exp_f := 1;
        ELSIF x =- 15692 THEN
            exp_f := 1;
        ELSIF x =- 15691 THEN
            exp_f := 1;
        ELSIF x =- 15690 THEN
            exp_f := 1;
        ELSIF x =- 15689 THEN
            exp_f := 1;
        ELSIF x =- 15688 THEN
            exp_f := 1;
        ELSIF x =- 15687 THEN
            exp_f := 1;
        ELSIF x =- 15686 THEN
            exp_f := 1;
        ELSIF x =- 15685 THEN
            exp_f := 1;
        ELSIF x =- 15684 THEN
            exp_f := 1;
        ELSIF x =- 15683 THEN
            exp_f := 1;
        ELSIF x =- 15682 THEN
            exp_f := 1;
        ELSIF x =- 15681 THEN
            exp_f := 1;
        ELSIF x =- 15680 THEN
            exp_f := 1;
        ELSIF x =- 15679 THEN
            exp_f := 1;
        ELSIF x =- 15678 THEN
            exp_f := 1;
        ELSIF x =- 15677 THEN
            exp_f := 1;
        ELSIF x =- 15676 THEN
            exp_f := 1;
        ELSIF x =- 15675 THEN
            exp_f := 1;
        ELSIF x =- 15674 THEN
            exp_f := 1;
        ELSIF x =- 15673 THEN
            exp_f := 1;
        ELSIF x =- 15672 THEN
            exp_f := 1;
        ELSIF x =- 15671 THEN
            exp_f := 1;
        ELSIF x =- 15670 THEN
            exp_f := 1;
        ELSIF x =- 15669 THEN
            exp_f := 1;
        ELSIF x =- 15668 THEN
            exp_f := 1;
        ELSIF x =- 15667 THEN
            exp_f := 1;
        ELSIF x =- 15666 THEN
            exp_f := 1;
        ELSIF x =- 15665 THEN
            exp_f := 1;
        ELSIF x =- 15664 THEN
            exp_f := 1;
        ELSIF x =- 15663 THEN
            exp_f := 1;
        ELSIF x =- 15662 THEN
            exp_f := 1;
        ELSIF x =- 15661 THEN
            exp_f := 1;
        ELSIF x =- 15660 THEN
            exp_f := 1;
        ELSIF x =- 15659 THEN
            exp_f := 1;
        ELSIF x =- 15658 THEN
            exp_f := 1;
        ELSIF x =- 15657 THEN
            exp_f := 1;
        ELSIF x =- 15656 THEN
            exp_f := 1;
        ELSIF x =- 15655 THEN
            exp_f := 1;
        ELSIF x =- 15654 THEN
            exp_f := 1;
        ELSIF x =- 15653 THEN
            exp_f := 1;
        ELSIF x =- 15652 THEN
            exp_f := 1;
        ELSIF x =- 15651 THEN
            exp_f := 1;
        ELSIF x =- 15650 THEN
            exp_f := 1;
        ELSIF x =- 15649 THEN
            exp_f := 1;
        ELSIF x =- 15648 THEN
            exp_f := 1;
        ELSIF x =- 15647 THEN
            exp_f := 1;
        ELSIF x =- 15646 THEN
            exp_f := 1;
        ELSIF x =- 15645 THEN
            exp_f := 1;
        ELSIF x =- 15644 THEN
            exp_f := 1;
        ELSIF x =- 15643 THEN
            exp_f := 1;
        ELSIF x =- 15642 THEN
            exp_f := 1;
        ELSIF x =- 15641 THEN
            exp_f := 1;
        ELSIF x =- 15640 THEN
            exp_f := 1;
        ELSIF x =- 15639 THEN
            exp_f := 1;
        ELSIF x =- 15638 THEN
            exp_f := 1;
        ELSIF x =- 15637 THEN
            exp_f := 1;
        ELSIF x =- 15636 THEN
            exp_f := 1;
        ELSIF x =- 15635 THEN
            exp_f := 1;
        ELSIF x =- 15634 THEN
            exp_f := 1;
        ELSIF x =- 15633 THEN
            exp_f := 1;
        ELSIF x =- 15632 THEN
            exp_f := 1;
        ELSIF x =- 15631 THEN
            exp_f := 1;
        ELSIF x =- 15630 THEN
            exp_f := 1;
        ELSIF x =- 15629 THEN
            exp_f := 1;
        ELSIF x =- 15628 THEN
            exp_f := 1;
        ELSIF x =- 15627 THEN
            exp_f := 1;
        ELSIF x =- 15626 THEN
            exp_f := 1;
        ELSIF x =- 15625 THEN
            exp_f := 1;
        ELSIF x =- 15624 THEN
            exp_f := 1;
        ELSIF x =- 15623 THEN
            exp_f := 1;
        ELSIF x =- 15622 THEN
            exp_f := 1;
        ELSIF x =- 15621 THEN
            exp_f := 1;
        ELSIF x =- 15620 THEN
            exp_f := 1;
        ELSIF x =- 15619 THEN
            exp_f := 1;
        ELSIF x =- 15618 THEN
            exp_f := 1;
        ELSIF x =- 15617 THEN
            exp_f := 1;
        ELSIF x =- 15616 THEN
            exp_f := 1;
        ELSIF x =- 15615 THEN
            exp_f := 1;
        ELSIF x =- 15614 THEN
            exp_f := 1;
        ELSIF x =- 15613 THEN
            exp_f := 1;
        ELSIF x =- 15612 THEN
            exp_f := 1;
        ELSIF x =- 15611 THEN
            exp_f := 1;
        ELSIF x =- 15610 THEN
            exp_f := 1;
        ELSIF x =- 15609 THEN
            exp_f := 1;
        ELSIF x =- 15608 THEN
            exp_f := 1;
        ELSIF x =- 15607 THEN
            exp_f := 1;
        ELSIF x =- 15606 THEN
            exp_f := 1;
        ELSIF x =- 15605 THEN
            exp_f := 1;
        ELSIF x =- 15604 THEN
            exp_f := 1;
        ELSIF x =- 15603 THEN
            exp_f := 1;
        ELSIF x =- 15602 THEN
            exp_f := 1;
        ELSIF x =- 15601 THEN
            exp_f := 1;
        ELSIF x =- 15600 THEN
            exp_f := 1;
        ELSIF x =- 15599 THEN
            exp_f := 1;
        ELSIF x =- 15598 THEN
            exp_f := 1;
        ELSIF x =- 15597 THEN
            exp_f := 1;
        ELSIF x =- 15596 THEN
            exp_f := 1;
        ELSIF x =- 15595 THEN
            exp_f := 1;
        ELSIF x =- 15594 THEN
            exp_f := 1;
        ELSIF x =- 15593 THEN
            exp_f := 1;
        ELSIF x =- 15592 THEN
            exp_f := 1;
        ELSIF x =- 15591 THEN
            exp_f := 1;
        ELSIF x =- 15590 THEN
            exp_f := 1;
        ELSIF x =- 15589 THEN
            exp_f := 1;
        ELSIF x =- 15588 THEN
            exp_f := 1;
        ELSIF x =- 15587 THEN
            exp_f := 1;
        ELSIF x =- 15586 THEN
            exp_f := 1;
        ELSIF x =- 15585 THEN
            exp_f := 1;
        ELSIF x =- 15584 THEN
            exp_f := 1;
        ELSIF x =- 15583 THEN
            exp_f := 1;
        ELSIF x =- 15582 THEN
            exp_f := 1;
        ELSIF x =- 15581 THEN
            exp_f := 1;
        ELSIF x =- 15580 THEN
            exp_f := 1;
        ELSIF x =- 15579 THEN
            exp_f := 1;
        ELSIF x =- 15578 THEN
            exp_f := 1;
        ELSIF x =- 15577 THEN
            exp_f := 1;
        ELSIF x =- 15576 THEN
            exp_f := 1;
        ELSIF x =- 15575 THEN
            exp_f := 1;
        ELSIF x =- 15574 THEN
            exp_f := 1;
        ELSIF x =- 15573 THEN
            exp_f := 1;
        ELSIF x =- 15572 THEN
            exp_f := 1;
        ELSIF x =- 15571 THEN
            exp_f := 1;
        ELSIF x =- 15570 THEN
            exp_f := 1;
        ELSIF x =- 15569 THEN
            exp_f := 1;
        ELSIF x =- 15568 THEN
            exp_f := 1;
        ELSIF x =- 15567 THEN
            exp_f := 1;
        ELSIF x =- 15566 THEN
            exp_f := 1;
        ELSIF x =- 15565 THEN
            exp_f := 1;
        ELSIF x =- 15564 THEN
            exp_f := 1;
        ELSIF x =- 15563 THEN
            exp_f := 1;
        ELSIF x =- 15562 THEN
            exp_f := 1;
        ELSIF x =- 15561 THEN
            exp_f := 1;
        ELSIF x =- 15560 THEN
            exp_f := 1;
        ELSIF x =- 15559 THEN
            exp_f := 1;
        ELSIF x =- 15558 THEN
            exp_f := 1;
        ELSIF x =- 15557 THEN
            exp_f := 1;
        ELSIF x =- 15556 THEN
            exp_f := 1;
        ELSIF x =- 15555 THEN
            exp_f := 1;
        ELSIF x =- 15554 THEN
            exp_f := 1;
        ELSIF x =- 15553 THEN
            exp_f := 1;
        ELSIF x =- 15552 THEN
            exp_f := 1;
        ELSIF x =- 15551 THEN
            exp_f := 1;
        ELSIF x =- 15550 THEN
            exp_f := 1;
        ELSIF x =- 15549 THEN
            exp_f := 1;
        ELSIF x =- 15548 THEN
            exp_f := 1;
        ELSIF x =- 15547 THEN
            exp_f := 1;
        ELSIF x =- 15546 THEN
            exp_f := 1;
        ELSIF x =- 15545 THEN
            exp_f := 1;
        ELSIF x =- 15544 THEN
            exp_f := 1;
        ELSIF x =- 15543 THEN
            exp_f := 1;
        ELSIF x =- 15542 THEN
            exp_f := 1;
        ELSIF x =- 15541 THEN
            exp_f := 1;
        ELSIF x =- 15540 THEN
            exp_f := 1;
        ELSIF x =- 15539 THEN
            exp_f := 1;
        ELSIF x =- 15538 THEN
            exp_f := 1;
        ELSIF x =- 15537 THEN
            exp_f := 1;
        ELSIF x =- 15536 THEN
            exp_f := 1;
        ELSIF x =- 15535 THEN
            exp_f := 1;
        ELSIF x =- 15534 THEN
            exp_f := 1;
        ELSIF x =- 15533 THEN
            exp_f := 1;
        ELSIF x =- 15532 THEN
            exp_f := 1;
        ELSIF x =- 15531 THEN
            exp_f := 1;
        ELSIF x =- 15530 THEN
            exp_f := 1;
        ELSIF x =- 15529 THEN
            exp_f := 1;
        ELSIF x =- 15528 THEN
            exp_f := 1;
        ELSIF x =- 15527 THEN
            exp_f := 1;
        ELSIF x =- 15526 THEN
            exp_f := 1;
        ELSIF x =- 15525 THEN
            exp_f := 1;
        ELSIF x =- 15524 THEN
            exp_f := 1;
        ELSIF x =- 15523 THEN
            exp_f := 1;
        ELSIF x =- 15522 THEN
            exp_f := 1;
        ELSIF x =- 15521 THEN
            exp_f := 1;
        ELSIF x =- 15520 THEN
            exp_f := 1;
        ELSIF x =- 15519 THEN
            exp_f := 1;
        ELSIF x =- 15518 THEN
            exp_f := 1;
        ELSIF x =- 15517 THEN
            exp_f := 1;
        ELSIF x =- 15516 THEN
            exp_f := 1;
        ELSIF x =- 15515 THEN
            exp_f := 1;
        ELSIF x =- 15514 THEN
            exp_f := 1;
        ELSIF x =- 15513 THEN
            exp_f := 1;
        ELSIF x =- 15512 THEN
            exp_f := 1;
        ELSIF x =- 15511 THEN
            exp_f := 1;
        ELSIF x =- 15510 THEN
            exp_f := 1;
        ELSIF x =- 15509 THEN
            exp_f := 1;
        ELSIF x =- 15508 THEN
            exp_f := 1;
        ELSIF x =- 15507 THEN
            exp_f := 1;
        ELSIF x =- 15506 THEN
            exp_f := 1;
        ELSIF x =- 15505 THEN
            exp_f := 1;
        ELSIF x =- 15504 THEN
            exp_f := 1;
        ELSIF x =- 15503 THEN
            exp_f := 1;
        ELSIF x =- 15502 THEN
            exp_f := 1;
        ELSIF x =- 15501 THEN
            exp_f := 1;
        ELSIF x =- 15500 THEN
            exp_f := 1;
        ELSIF x =- 15499 THEN
            exp_f := 1;
        ELSIF x =- 15498 THEN
            exp_f := 1;
        ELSIF x =- 15497 THEN
            exp_f := 1;
        ELSIF x =- 15496 THEN
            exp_f := 1;
        ELSIF x =- 15495 THEN
            exp_f := 1;
        ELSIF x =- 15494 THEN
            exp_f := 1;
        ELSIF x =- 15493 THEN
            exp_f := 1;
        ELSIF x =- 15492 THEN
            exp_f := 1;
        ELSIF x =- 15491 THEN
            exp_f := 1;
        ELSIF x =- 15490 THEN
            exp_f := 1;
        ELSIF x =- 15489 THEN
            exp_f := 1;
        ELSIF x =- 15488 THEN
            exp_f := 1;
        ELSIF x =- 15487 THEN
            exp_f := 1;
        ELSIF x =- 15486 THEN
            exp_f := 1;
        ELSIF x =- 15485 THEN
            exp_f := 1;
        ELSIF x =- 15484 THEN
            exp_f := 1;
        ELSIF x =- 15483 THEN
            exp_f := 1;
        ELSIF x =- 15482 THEN
            exp_f := 1;
        ELSIF x =- 15481 THEN
            exp_f := 1;
        ELSIF x =- 15480 THEN
            exp_f := 1;
        ELSIF x =- 15479 THEN
            exp_f := 1;
        ELSIF x =- 15478 THEN
            exp_f := 1;
        ELSIF x =- 15477 THEN
            exp_f := 1;
        ELSIF x =- 15476 THEN
            exp_f := 1;
        ELSIF x =- 15475 THEN
            exp_f := 1;
        ELSIF x =- 15474 THEN
            exp_f := 1;
        ELSIF x =- 15473 THEN
            exp_f := 1;
        ELSIF x =- 15472 THEN
            exp_f := 1;
        ELSIF x =- 15471 THEN
            exp_f := 1;
        ELSIF x =- 15470 THEN
            exp_f := 1;
        ELSIF x =- 15469 THEN
            exp_f := 1;
        ELSIF x =- 15468 THEN
            exp_f := 1;
        ELSIF x =- 15467 THEN
            exp_f := 1;
        ELSIF x =- 15466 THEN
            exp_f := 1;
        ELSIF x =- 15465 THEN
            exp_f := 1;
        ELSIF x =- 15464 THEN
            exp_f := 1;
        ELSIF x =- 15463 THEN
            exp_f := 1;
        ELSIF x =- 15462 THEN
            exp_f := 1;
        ELSIF x =- 15461 THEN
            exp_f := 1;
        ELSIF x =- 15460 THEN
            exp_f := 1;
        ELSIF x =- 15459 THEN
            exp_f := 1;
        ELSIF x =- 15458 THEN
            exp_f := 1;
        ELSIF x =- 15457 THEN
            exp_f := 1;
        ELSIF x =- 15456 THEN
            exp_f := 1;
        ELSIF x =- 15455 THEN
            exp_f := 1;
        ELSIF x =- 15454 THEN
            exp_f := 1;
        ELSIF x =- 15453 THEN
            exp_f := 1;
        ELSIF x =- 15452 THEN
            exp_f := 1;
        ELSIF x =- 15451 THEN
            exp_f := 1;
        ELSIF x =- 15450 THEN
            exp_f := 1;
        ELSIF x =- 15449 THEN
            exp_f := 1;
        ELSIF x =- 15448 THEN
            exp_f := 1;
        ELSIF x =- 15447 THEN
            exp_f := 1;
        ELSIF x =- 15446 THEN
            exp_f := 1;
        ELSIF x =- 15445 THEN
            exp_f := 1;
        ELSIF x =- 15444 THEN
            exp_f := 1;
        ELSIF x =- 15443 THEN
            exp_f := 1;
        ELSIF x =- 15442 THEN
            exp_f := 1;
        ELSIF x =- 15441 THEN
            exp_f := 1;
        ELSIF x =- 15440 THEN
            exp_f := 1;
        ELSIF x =- 15439 THEN
            exp_f := 1;
        ELSIF x =- 15438 THEN
            exp_f := 1;
        ELSIF x =- 15437 THEN
            exp_f := 1;
        ELSIF x =- 15436 THEN
            exp_f := 1;
        ELSIF x =- 15435 THEN
            exp_f := 1;
        ELSIF x =- 15434 THEN
            exp_f := 1;
        ELSIF x =- 15433 THEN
            exp_f := 1;
        ELSIF x =- 15432 THEN
            exp_f := 1;
        ELSIF x =- 15431 THEN
            exp_f := 1;
        ELSIF x =- 15430 THEN
            exp_f := 1;
        ELSIF x =- 15429 THEN
            exp_f := 1;
        ELSIF x =- 15428 THEN
            exp_f := 1;
        ELSIF x =- 15427 THEN
            exp_f := 1;
        ELSIF x =- 15426 THEN
            exp_f := 1;
        ELSIF x =- 15425 THEN
            exp_f := 1;
        ELSIF x =- 15424 THEN
            exp_f := 1;
        ELSIF x =- 15423 THEN
            exp_f := 1;
        ELSIF x =- 15422 THEN
            exp_f := 1;
        ELSIF x =- 15421 THEN
            exp_f := 1;
        ELSIF x =- 15420 THEN
            exp_f := 1;
        ELSIF x =- 15419 THEN
            exp_f := 1;
        ELSIF x =- 15418 THEN
            exp_f := 1;
        ELSIF x =- 15417 THEN
            exp_f := 1;
        ELSIF x =- 15416 THEN
            exp_f := 1;
        ELSIF x =- 15415 THEN
            exp_f := 1;
        ELSIF x =- 15414 THEN
            exp_f := 1;
        ELSIF x =- 15413 THEN
            exp_f := 1;
        ELSIF x =- 15412 THEN
            exp_f := 1;
        ELSIF x =- 15411 THEN
            exp_f := 1;
        ELSIF x =- 15410 THEN
            exp_f := 1;
        ELSIF x =- 15409 THEN
            exp_f := 1;
        ELSIF x =- 15408 THEN
            exp_f := 1;
        ELSIF x =- 15407 THEN
            exp_f := 1;
        ELSIF x =- 15406 THEN
            exp_f := 1;
        ELSIF x =- 15405 THEN
            exp_f := 1;
        ELSIF x =- 15404 THEN
            exp_f := 1;
        ELSIF x =- 15403 THEN
            exp_f := 1;
        ELSIF x =- 15402 THEN
            exp_f := 1;
        ELSIF x =- 15401 THEN
            exp_f := 1;
        ELSIF x =- 15400 THEN
            exp_f := 1;
        ELSIF x =- 15399 THEN
            exp_f := 1;
        ELSIF x =- 15398 THEN
            exp_f := 1;
        ELSIF x =- 15397 THEN
            exp_f := 1;
        ELSIF x =- 15396 THEN
            exp_f := 1;
        ELSIF x =- 15395 THEN
            exp_f := 1;
        ELSIF x =- 15394 THEN
            exp_f := 1;
        ELSIF x =- 15393 THEN
            exp_f := 1;
        ELSIF x =- 15392 THEN
            exp_f := 1;
        ELSIF x =- 15391 THEN
            exp_f := 1;
        ELSIF x =- 15390 THEN
            exp_f := 1;
        ELSIF x =- 15389 THEN
            exp_f := 1;
        ELSIF x =- 15388 THEN
            exp_f := 1;
        ELSIF x =- 15387 THEN
            exp_f := 1;
        ELSIF x =- 15386 THEN
            exp_f := 1;
        ELSIF x =- 15385 THEN
            exp_f := 1;
        ELSIF x =- 15384 THEN
            exp_f := 1;
        ELSIF x =- 15383 THEN
            exp_f := 1;
        ELSIF x =- 15382 THEN
            exp_f := 1;
        ELSIF x =- 15381 THEN
            exp_f := 1;
        ELSIF x =- 15380 THEN
            exp_f := 1;
        ELSIF x =- 15379 THEN
            exp_f := 1;
        ELSIF x =- 15378 THEN
            exp_f := 1;
        ELSIF x =- 15377 THEN
            exp_f := 1;
        ELSIF x =- 15376 THEN
            exp_f := 1;
        ELSIF x =- 15375 THEN
            exp_f := 1;
        ELSIF x =- 15374 THEN
            exp_f := 1;
        ELSIF x =- 15373 THEN
            exp_f := 1;
        ELSIF x =- 15372 THEN
            exp_f := 1;
        ELSIF x =- 15371 THEN
            exp_f := 1;
        ELSIF x =- 15370 THEN
            exp_f := 1;
        ELSIF x =- 15369 THEN
            exp_f := 1;
        ELSIF x =- 15368 THEN
            exp_f := 1;
        ELSIF x =- 15367 THEN
            exp_f := 1;
        ELSIF x =- 15366 THEN
            exp_f := 1;
        ELSIF x =- 15365 THEN
            exp_f := 1;
        ELSIF x =- 15364 THEN
            exp_f := 1;
        ELSIF x =- 15363 THEN
            exp_f := 1;
        ELSIF x =- 15362 THEN
            exp_f := 1;
        ELSIF x =- 15361 THEN
            exp_f := 1;
        ELSIF x =- 15360 THEN
            exp_f := 1;
        ELSIF x =- 15359 THEN
            exp_f := 1;
        ELSIF x =- 15358 THEN
            exp_f := 1;
        ELSIF x =- 15357 THEN
            exp_f := 1;
        ELSIF x =- 15356 THEN
            exp_f := 1;
        ELSIF x =- 15355 THEN
            exp_f := 1;
        ELSIF x =- 15354 THEN
            exp_f := 1;
        ELSIF x =- 15353 THEN
            exp_f := 1;
        ELSIF x =- 15352 THEN
            exp_f := 1;
        ELSIF x =- 15351 THEN
            exp_f := 1;
        ELSIF x =- 15350 THEN
            exp_f := 1;
        ELSIF x =- 15349 THEN
            exp_f := 1;
        ELSIF x =- 15348 THEN
            exp_f := 1;
        ELSIF x =- 15347 THEN
            exp_f := 1;
        ELSIF x =- 15346 THEN
            exp_f := 1;
        ELSIF x =- 15345 THEN
            exp_f := 1;
        ELSIF x =- 15344 THEN
            exp_f := 1;
        ELSIF x =- 15343 THEN
            exp_f := 1;
        ELSIF x =- 15342 THEN
            exp_f := 1;
        ELSIF x =- 15341 THEN
            exp_f := 1;
        ELSIF x =- 15340 THEN
            exp_f := 1;
        ELSIF x =- 15339 THEN
            exp_f := 1;
        ELSIF x =- 15338 THEN
            exp_f := 1;
        ELSIF x =- 15337 THEN
            exp_f := 1;
        ELSIF x =- 15336 THEN
            exp_f := 1;
        ELSIF x =- 15335 THEN
            exp_f := 1;
        ELSIF x =- 15334 THEN
            exp_f := 1;
        ELSIF x =- 15333 THEN
            exp_f := 1;
        ELSIF x =- 15332 THEN
            exp_f := 1;
        ELSIF x =- 15331 THEN
            exp_f := 1;
        ELSIF x =- 15330 THEN
            exp_f := 1;
        ELSIF x =- 15329 THEN
            exp_f := 1;
        ELSIF x =- 15328 THEN
            exp_f := 1;
        ELSIF x =- 15327 THEN
            exp_f := 1;
        ELSIF x =- 15326 THEN
            exp_f := 1;
        ELSIF x =- 15325 THEN
            exp_f := 1;
        ELSIF x =- 15324 THEN
            exp_f := 1;
        ELSIF x =- 15323 THEN
            exp_f := 1;
        ELSIF x =- 15322 THEN
            exp_f := 1;
        ELSIF x =- 15321 THEN
            exp_f := 1;
        ELSIF x =- 15320 THEN
            exp_f := 1;
        ELSIF x =- 15319 THEN
            exp_f := 1;
        ELSIF x =- 15318 THEN
            exp_f := 1;
        ELSIF x =- 15317 THEN
            exp_f := 1;
        ELSIF x =- 15316 THEN
            exp_f := 1;
        ELSIF x =- 15315 THEN
            exp_f := 1;
        ELSIF x =- 15314 THEN
            exp_f := 1;
        ELSIF x =- 15313 THEN
            exp_f := 1;
        ELSIF x =- 15312 THEN
            exp_f := 1;
        ELSIF x =- 15311 THEN
            exp_f := 1;
        ELSIF x =- 15310 THEN
            exp_f := 1;
        ELSIF x =- 15309 THEN
            exp_f := 1;
        ELSIF x =- 15308 THEN
            exp_f := 1;
        ELSIF x =- 15307 THEN
            exp_f := 1;
        ELSIF x =- 15306 THEN
            exp_f := 1;
        ELSIF x =- 15305 THEN
            exp_f := 1;
        ELSIF x =- 15304 THEN
            exp_f := 1;
        ELSIF x =- 15303 THEN
            exp_f := 1;
        ELSIF x =- 15302 THEN
            exp_f := 1;
        ELSIF x =- 15301 THEN
            exp_f := 1;
        ELSIF x =- 15300 THEN
            exp_f := 1;
        ELSIF x =- 15299 THEN
            exp_f := 1;
        ELSIF x =- 15298 THEN
            exp_f := 1;
        ELSIF x =- 15297 THEN
            exp_f := 1;
        ELSIF x =- 15296 THEN
            exp_f := 1;
        ELSIF x =- 15295 THEN
            exp_f := 1;
        ELSIF x =- 15294 THEN
            exp_f := 1;
        ELSIF x =- 15293 THEN
            exp_f := 1;
        ELSIF x =- 15292 THEN
            exp_f := 1;
        ELSIF x =- 15291 THEN
            exp_f := 1;
        ELSIF x =- 15290 THEN
            exp_f := 1;
        ELSIF x =- 15289 THEN
            exp_f := 1;
        ELSIF x =- 15288 THEN
            exp_f := 1;
        ELSIF x =- 15287 THEN
            exp_f := 1;
        ELSIF x =- 15286 THEN
            exp_f := 1;
        ELSIF x =- 15285 THEN
            exp_f := 1;
        ELSIF x =- 15284 THEN
            exp_f := 1;
        ELSIF x =- 15283 THEN
            exp_f := 1;
        ELSIF x =- 15282 THEN
            exp_f := 1;
        ELSIF x =- 15281 THEN
            exp_f := 1;
        ELSIF x =- 15280 THEN
            exp_f := 1;
        ELSIF x =- 15279 THEN
            exp_f := 1;
        ELSIF x =- 15278 THEN
            exp_f := 1;
        ELSIF x =- 15277 THEN
            exp_f := 1;
        ELSIF x =- 15276 THEN
            exp_f := 1;
        ELSIF x =- 15275 THEN
            exp_f := 1;
        ELSIF x =- 15274 THEN
            exp_f := 1;
        ELSIF x =- 15273 THEN
            exp_f := 1;
        ELSIF x =- 15272 THEN
            exp_f := 1;
        ELSIF x =- 15271 THEN
            exp_f := 1;
        ELSIF x =- 15270 THEN
            exp_f := 1;
        ELSIF x =- 15269 THEN
            exp_f := 1;
        ELSIF x =- 15268 THEN
            exp_f := 1;
        ELSIF x =- 15267 THEN
            exp_f := 1;
        ELSIF x =- 15266 THEN
            exp_f := 1;
        ELSIF x =- 15265 THEN
            exp_f := 1;
        ELSIF x =- 15264 THEN
            exp_f := 1;
        ELSIF x =- 15263 THEN
            exp_f := 1;
        ELSIF x =- 15262 THEN
            exp_f := 1;
        ELSIF x =- 15261 THEN
            exp_f := 1;
        ELSIF x =- 15260 THEN
            exp_f := 1;
        ELSIF x =- 15259 THEN
            exp_f := 1;
        ELSIF x =- 15258 THEN
            exp_f := 1;
        ELSIF x =- 15257 THEN
            exp_f := 1;
        ELSIF x =- 15256 THEN
            exp_f := 1;
        ELSIF x =- 15255 THEN
            exp_f := 1;
        ELSIF x =- 15254 THEN
            exp_f := 1;
        ELSIF x =- 15253 THEN
            exp_f := 1;
        ELSIF x =- 15252 THEN
            exp_f := 1;
        ELSIF x =- 15251 THEN
            exp_f := 1;
        ELSIF x =- 15250 THEN
            exp_f := 1;
        ELSIF x =- 15249 THEN
            exp_f := 1;
        ELSIF x =- 15248 THEN
            exp_f := 1;
        ELSIF x =- 15247 THEN
            exp_f := 1;
        ELSIF x =- 15246 THEN
            exp_f := 1;
        ELSIF x =- 15245 THEN
            exp_f := 1;
        ELSIF x =- 15244 THEN
            exp_f := 1;
        ELSIF x =- 15243 THEN
            exp_f := 1;
        ELSIF x =- 15242 THEN
            exp_f := 1;
        ELSIF x =- 15241 THEN
            exp_f := 1;
        ELSIF x =- 15240 THEN
            exp_f := 1;
        ELSIF x =- 15239 THEN
            exp_f := 1;
        ELSIF x =- 15238 THEN
            exp_f := 1;
        ELSIF x =- 15237 THEN
            exp_f := 1;
        ELSIF x =- 15236 THEN
            exp_f := 1;
        ELSIF x =- 15235 THEN
            exp_f := 1;
        ELSIF x =- 15234 THEN
            exp_f := 1;
        ELSIF x =- 15233 THEN
            exp_f := 1;
        ELSIF x =- 15232 THEN
            exp_f := 1;
        ELSIF x =- 15231 THEN
            exp_f := 1;
        ELSIF x =- 15230 THEN
            exp_f := 1;
        ELSIF x =- 15229 THEN
            exp_f := 1;
        ELSIF x =- 15228 THEN
            exp_f := 1;
        ELSIF x =- 15227 THEN
            exp_f := 1;
        ELSIF x =- 15226 THEN
            exp_f := 1;
        ELSIF x =- 15225 THEN
            exp_f := 1;
        ELSIF x =- 15224 THEN
            exp_f := 1;
        ELSIF x =- 15223 THEN
            exp_f := 1;
        ELSIF x =- 15222 THEN
            exp_f := 1;
        ELSIF x =- 15221 THEN
            exp_f := 1;
        ELSIF x =- 15220 THEN
            exp_f := 1;
        ELSIF x =- 15219 THEN
            exp_f := 1;
        ELSIF x =- 15218 THEN
            exp_f := 1;
        ELSIF x =- 15217 THEN
            exp_f := 1;
        ELSIF x =- 15216 THEN
            exp_f := 1;
        ELSIF x =- 15215 THEN
            exp_f := 1;
        ELSIF x =- 15214 THEN
            exp_f := 1;
        ELSIF x =- 15213 THEN
            exp_f := 1;
        ELSIF x =- 15212 THEN
            exp_f := 1;
        ELSIF x =- 15211 THEN
            exp_f := 1;
        ELSIF x =- 15210 THEN
            exp_f := 1;
        ELSIF x =- 15209 THEN
            exp_f := 1;
        ELSIF x =- 15208 THEN
            exp_f := 1;
        ELSIF x =- 15207 THEN
            exp_f := 1;
        ELSIF x =- 15206 THEN
            exp_f := 1;
        ELSIF x =- 15205 THEN
            exp_f := 1;
        ELSIF x =- 15204 THEN
            exp_f := 1;
        ELSIF x =- 15203 THEN
            exp_f := 1;
        ELSIF x =- 15202 THEN
            exp_f := 1;
        ELSIF x =- 15201 THEN
            exp_f := 1;
        ELSIF x =- 15200 THEN
            exp_f := 1;
        ELSIF x =- 15199 THEN
            exp_f := 1;
        ELSIF x =- 15198 THEN
            exp_f := 1;
        ELSIF x =- 15197 THEN
            exp_f := 1;
        ELSIF x =- 15196 THEN
            exp_f := 1;
        ELSIF x =- 15195 THEN
            exp_f := 1;
        ELSIF x =- 15194 THEN
            exp_f := 1;
        ELSIF x =- 15193 THEN
            exp_f := 1;
        ELSIF x =- 15192 THEN
            exp_f := 1;
        ELSIF x =- 15191 THEN
            exp_f := 1;
        ELSIF x =- 15190 THEN
            exp_f := 1;
        ELSIF x =- 15189 THEN
            exp_f := 1;
        ELSIF x =- 15188 THEN
            exp_f := 1;
        ELSIF x =- 15187 THEN
            exp_f := 1;
        ELSIF x =- 15186 THEN
            exp_f := 1;
        ELSIF x =- 15185 THEN
            exp_f := 1;
        ELSIF x =- 15184 THEN
            exp_f := 1;
        ELSIF x =- 15183 THEN
            exp_f := 1;
        ELSIF x =- 15182 THEN
            exp_f := 1;
        ELSIF x =- 15181 THEN
            exp_f := 1;
        ELSIF x =- 15180 THEN
            exp_f := 1;
        ELSIF x =- 15179 THEN
            exp_f := 1;
        ELSIF x =- 15178 THEN
            exp_f := 1;
        ELSIF x =- 15177 THEN
            exp_f := 1;
        ELSIF x =- 15176 THEN
            exp_f := 1;
        ELSIF x =- 15175 THEN
            exp_f := 1;
        ELSIF x =- 15174 THEN
            exp_f := 1;
        ELSIF x =- 15173 THEN
            exp_f := 1;
        ELSIF x =- 15172 THEN
            exp_f := 1;
        ELSIF x =- 15171 THEN
            exp_f := 1;
        ELSIF x =- 15170 THEN
            exp_f := 1;
        ELSIF x =- 15169 THEN
            exp_f := 1;
        ELSIF x =- 15168 THEN
            exp_f := 1;
        ELSIF x =- 15167 THEN
            exp_f := 1;
        ELSIF x =- 15166 THEN
            exp_f := 1;
        ELSIF x =- 15165 THEN
            exp_f := 1;
        ELSIF x =- 15164 THEN
            exp_f := 1;
        ELSIF x =- 15163 THEN
            exp_f := 1;
        ELSIF x =- 15162 THEN
            exp_f := 1;
        ELSIF x =- 15161 THEN
            exp_f := 1;
        ELSIF x =- 15160 THEN
            exp_f := 1;
        ELSIF x =- 15159 THEN
            exp_f := 1;
        ELSIF x =- 15158 THEN
            exp_f := 1;
        ELSIF x =- 15157 THEN
            exp_f := 1;
        ELSIF x =- 15156 THEN
            exp_f := 1;
        ELSIF x =- 15155 THEN
            exp_f := 1;
        ELSIF x =- 15154 THEN
            exp_f := 1;
        ELSIF x =- 15153 THEN
            exp_f := 1;
        ELSIF x =- 15152 THEN
            exp_f := 1;
        ELSIF x =- 15151 THEN
            exp_f := 1;
        ELSIF x =- 15150 THEN
            exp_f := 1;
        ELSIF x =- 15149 THEN
            exp_f := 1;
        ELSIF x =- 15148 THEN
            exp_f := 1;
        ELSIF x =- 15147 THEN
            exp_f := 1;
        ELSIF x =- 15146 THEN
            exp_f := 1;
        ELSIF x =- 15145 THEN
            exp_f := 1;
        ELSIF x =- 15144 THEN
            exp_f := 1;
        ELSIF x =- 15143 THEN
            exp_f := 1;
        ELSIF x =- 15142 THEN
            exp_f := 1;
        ELSIF x =- 15141 THEN
            exp_f := 1;
        ELSIF x =- 15140 THEN
            exp_f := 1;
        ELSIF x =- 15139 THEN
            exp_f := 1;
        ELSIF x =- 15138 THEN
            exp_f := 1;
        ELSIF x =- 15137 THEN
            exp_f := 1;
        ELSIF x =- 15136 THEN
            exp_f := 1;
        ELSIF x =- 15135 THEN
            exp_f := 1;
        ELSIF x =- 15134 THEN
            exp_f := 1;
        ELSIF x =- 15133 THEN
            exp_f := 1;
        ELSIF x =- 15132 THEN
            exp_f := 1;
        ELSIF x =- 15131 THEN
            exp_f := 1;
        ELSIF x =- 15130 THEN
            exp_f := 1;
        ELSIF x =- 15129 THEN
            exp_f := 1;
        ELSIF x =- 15128 THEN
            exp_f := 1;
        ELSIF x =- 15127 THEN
            exp_f := 1;
        ELSIF x =- 15126 THEN
            exp_f := 1;
        ELSIF x =- 15125 THEN
            exp_f := 1;
        ELSIF x =- 15124 THEN
            exp_f := 1;
        ELSIF x =- 15123 THEN
            exp_f := 1;
        ELSIF x =- 15122 THEN
            exp_f := 1;
        ELSIF x =- 15121 THEN
            exp_f := 1;
        ELSIF x =- 15120 THEN
            exp_f := 1;
        ELSIF x =- 15119 THEN
            exp_f := 1;
        ELSIF x =- 15118 THEN
            exp_f := 1;
        ELSIF x =- 15117 THEN
            exp_f := 1;
        ELSIF x =- 15116 THEN
            exp_f := 1;
        ELSIF x =- 15115 THEN
            exp_f := 1;
        ELSIF x =- 15114 THEN
            exp_f := 1;
        ELSIF x =- 15113 THEN
            exp_f := 1;
        ELSIF x =- 15112 THEN
            exp_f := 1;
        ELSIF x =- 15111 THEN
            exp_f := 1;
        ELSIF x =- 15110 THEN
            exp_f := 1;
        ELSIF x =- 15109 THEN
            exp_f := 1;
        ELSIF x =- 15108 THEN
            exp_f := 1;
        ELSIF x =- 15107 THEN
            exp_f := 1;
        ELSIF x =- 15106 THEN
            exp_f := 1;
        ELSIF x =- 15105 THEN
            exp_f := 1;
        ELSIF x =- 15104 THEN
            exp_f := 1;
        ELSIF x =- 15103 THEN
            exp_f := 1;
        ELSIF x =- 15102 THEN
            exp_f := 1;
        ELSIF x =- 15101 THEN
            exp_f := 1;
        ELSIF x =- 15100 THEN
            exp_f := 1;
        ELSIF x =- 15099 THEN
            exp_f := 1;
        ELSIF x =- 15098 THEN
            exp_f := 1;
        ELSIF x =- 15097 THEN
            exp_f := 1;
        ELSIF x =- 15096 THEN
            exp_f := 1;
        ELSIF x =- 15095 THEN
            exp_f := 1;
        ELSIF x =- 15094 THEN
            exp_f := 1;
        ELSIF x =- 15093 THEN
            exp_f := 1;
        ELSIF x =- 15092 THEN
            exp_f := 1;
        ELSIF x =- 15091 THEN
            exp_f := 1;
        ELSIF x =- 15090 THEN
            exp_f := 1;
        ELSIF x =- 15089 THEN
            exp_f := 1;
        ELSIF x =- 15088 THEN
            exp_f := 1;
        ELSIF x =- 15087 THEN
            exp_f := 1;
        ELSIF x =- 15086 THEN
            exp_f := 1;
        ELSIF x =- 15085 THEN
            exp_f := 1;
        ELSIF x =- 15084 THEN
            exp_f := 1;
        ELSIF x =- 15083 THEN
            exp_f := 1;
        ELSIF x =- 15082 THEN
            exp_f := 1;
        ELSIF x =- 15081 THEN
            exp_f := 1;
        ELSIF x =- 15080 THEN
            exp_f := 1;
        ELSIF x =- 15079 THEN
            exp_f := 1;
        ELSIF x =- 15078 THEN
            exp_f := 1;
        ELSIF x =- 15077 THEN
            exp_f := 1;
        ELSIF x =- 15076 THEN
            exp_f := 1;
        ELSIF x =- 15075 THEN
            exp_f := 1;
        ELSIF x =- 15074 THEN
            exp_f := 1;
        ELSIF x =- 15073 THEN
            exp_f := 1;
        ELSIF x =- 15072 THEN
            exp_f := 1;
        ELSIF x =- 15071 THEN
            exp_f := 1;
        ELSIF x =- 15070 THEN
            exp_f := 1;
        ELSIF x =- 15069 THEN
            exp_f := 1;
        ELSIF x =- 15068 THEN
            exp_f := 1;
        ELSIF x =- 15067 THEN
            exp_f := 1;
        ELSIF x =- 15066 THEN
            exp_f := 1;
        ELSIF x =- 15065 THEN
            exp_f := 1;
        ELSIF x =- 15064 THEN
            exp_f := 1;
        ELSIF x =- 15063 THEN
            exp_f := 1;
        ELSIF x =- 15062 THEN
            exp_f := 1;
        ELSIF x =- 15061 THEN
            exp_f := 1;
        ELSIF x =- 15060 THEN
            exp_f := 1;
        ELSIF x =- 15059 THEN
            exp_f := 1;
        ELSIF x =- 15058 THEN
            exp_f := 1;
        ELSIF x =- 15057 THEN
            exp_f := 1;
        ELSIF x =- 15056 THEN
            exp_f := 1;
        ELSIF x =- 15055 THEN
            exp_f := 1;
        ELSIF x =- 15054 THEN
            exp_f := 1;
        ELSIF x =- 15053 THEN
            exp_f := 1;
        ELSIF x =- 15052 THEN
            exp_f := 1;
        ELSIF x =- 15051 THEN
            exp_f := 1;
        ELSIF x =- 15050 THEN
            exp_f := 1;
        ELSIF x =- 15049 THEN
            exp_f := 1;
        ELSIF x =- 15048 THEN
            exp_f := 1;
        ELSIF x =- 15047 THEN
            exp_f := 1;
        ELSIF x =- 15046 THEN
            exp_f := 1;
        ELSIF x =- 15045 THEN
            exp_f := 1;
        ELSIF x =- 15044 THEN
            exp_f := 1;
        ELSIF x =- 15043 THEN
            exp_f := 1;
        ELSIF x =- 15042 THEN
            exp_f := 1;
        ELSIF x =- 15041 THEN
            exp_f := 1;
        ELSIF x =- 15040 THEN
            exp_f := 1;
        ELSIF x =- 15039 THEN
            exp_f := 1;
        ELSIF x =- 15038 THEN
            exp_f := 1;
        ELSIF x =- 15037 THEN
            exp_f := 1;
        ELSIF x =- 15036 THEN
            exp_f := 1;
        ELSIF x =- 15035 THEN
            exp_f := 1;
        ELSIF x =- 15034 THEN
            exp_f := 1;
        ELSIF x =- 15033 THEN
            exp_f := 1;
        ELSIF x =- 15032 THEN
            exp_f := 1;
        ELSIF x =- 15031 THEN
            exp_f := 1;
        ELSIF x =- 15030 THEN
            exp_f := 1;
        ELSIF x =- 15029 THEN
            exp_f := 1;
        ELSIF x =- 15028 THEN
            exp_f := 1;
        ELSIF x =- 15027 THEN
            exp_f := 1;
        ELSIF x =- 15026 THEN
            exp_f := 1;
        ELSIF x =- 15025 THEN
            exp_f := 1;
        ELSIF x =- 15024 THEN
            exp_f := 1;
        ELSIF x =- 15023 THEN
            exp_f := 1;
        ELSIF x =- 15022 THEN
            exp_f := 1;
        ELSIF x =- 15021 THEN
            exp_f := 1;
        ELSIF x =- 15020 THEN
            exp_f := 1;
        ELSIF x =- 15019 THEN
            exp_f := 1;
        ELSIF x =- 15018 THEN
            exp_f := 1;
        ELSIF x =- 15017 THEN
            exp_f := 1;
        ELSIF x =- 15016 THEN
            exp_f := 1;
        ELSIF x =- 15015 THEN
            exp_f := 1;
        ELSIF x =- 15014 THEN
            exp_f := 1;
        ELSIF x =- 15013 THEN
            exp_f := 1;
        ELSIF x =- 15012 THEN
            exp_f := 1;
        ELSIF x =- 15011 THEN
            exp_f := 1;
        ELSIF x =- 15010 THEN
            exp_f := 1;
        ELSIF x =- 15009 THEN
            exp_f := 1;
        ELSIF x =- 15008 THEN
            exp_f := 1;
        ELSIF x =- 15007 THEN
            exp_f := 1;
        ELSIF x =- 15006 THEN
            exp_f := 1;
        ELSIF x =- 15005 THEN
            exp_f := 1;
        ELSIF x =- 15004 THEN
            exp_f := 1;
        ELSIF x =- 15003 THEN
            exp_f := 1;
        ELSIF x =- 15002 THEN
            exp_f := 1;
        ELSIF x =- 15001 THEN
            exp_f := 1;
        ELSIF x =- 15000 THEN
            exp_f := 1;
        ELSIF x =- 14999 THEN
            exp_f := 1;
        ELSIF x =- 14998 THEN
            exp_f := 1;
        ELSIF x =- 14997 THEN
            exp_f := 1;
        ELSIF x =- 14996 THEN
            exp_f := 1;
        ELSIF x =- 14995 THEN
            exp_f := 1;
        ELSIF x =- 14994 THEN
            exp_f := 1;
        ELSIF x =- 14993 THEN
            exp_f := 1;
        ELSIF x =- 14992 THEN
            exp_f := 1;
        ELSIF x =- 14991 THEN
            exp_f := 1;
        ELSIF x =- 14990 THEN
            exp_f := 1;
        ELSIF x =- 14989 THEN
            exp_f := 1;
        ELSIF x =- 14988 THEN
            exp_f := 1;
        ELSIF x =- 14987 THEN
            exp_f := 1;
        ELSIF x =- 14986 THEN
            exp_f := 1;
        ELSIF x =- 14985 THEN
            exp_f := 1;
        ELSIF x =- 14984 THEN
            exp_f := 1;
        ELSIF x =- 14983 THEN
            exp_f := 1;
        ELSIF x =- 14982 THEN
            exp_f := 1;
        ELSIF x =- 14981 THEN
            exp_f := 1;
        ELSIF x =- 14980 THEN
            exp_f := 1;
        ELSIF x =- 14979 THEN
            exp_f := 1;
        ELSIF x =- 14978 THEN
            exp_f := 1;
        ELSIF x =- 14977 THEN
            exp_f := 1;
        ELSIF x =- 14976 THEN
            exp_f := 1;
        ELSIF x =- 14975 THEN
            exp_f := 1;
        ELSIF x =- 14974 THEN
            exp_f := 1;
        ELSIF x =- 14973 THEN
            exp_f := 1;
        ELSIF x =- 14972 THEN
            exp_f := 1;
        ELSIF x =- 14971 THEN
            exp_f := 1;
        ELSIF x =- 14970 THEN
            exp_f := 1;
        ELSIF x =- 14969 THEN
            exp_f := 1;
        ELSIF x =- 14968 THEN
            exp_f := 1;
        ELSIF x =- 14967 THEN
            exp_f := 1;
        ELSIF x =- 14966 THEN
            exp_f := 1;
        ELSIF x =- 14965 THEN
            exp_f := 1;
        ELSIF x =- 14964 THEN
            exp_f := 1;
        ELSIF x =- 14963 THEN
            exp_f := 1;
        ELSIF x =- 14962 THEN
            exp_f := 1;
        ELSIF x =- 14961 THEN
            exp_f := 1;
        ELSIF x =- 14960 THEN
            exp_f := 1;
        ELSIF x =- 14959 THEN
            exp_f := 1;
        ELSIF x =- 14958 THEN
            exp_f := 1;
        ELSIF x =- 14957 THEN
            exp_f := 1;
        ELSIF x =- 14956 THEN
            exp_f := 1;
        ELSIF x =- 14955 THEN
            exp_f := 1;
        ELSIF x =- 14954 THEN
            exp_f := 1;
        ELSIF x =- 14953 THEN
            exp_f := 1;
        ELSIF x =- 14952 THEN
            exp_f := 1;
        ELSIF x =- 14951 THEN
            exp_f := 1;
        ELSIF x =- 14950 THEN
            exp_f := 1;
        ELSIF x =- 14949 THEN
            exp_f := 1;
        ELSIF x =- 14948 THEN
            exp_f := 1;
        ELSIF x =- 14947 THEN
            exp_f := 1;
        ELSIF x =- 14946 THEN
            exp_f := 1;
        ELSIF x =- 14945 THEN
            exp_f := 1;
        ELSIF x =- 14944 THEN
            exp_f := 1;
        ELSIF x =- 14943 THEN
            exp_f := 1;
        ELSIF x =- 14942 THEN
            exp_f := 1;
        ELSIF x =- 14941 THEN
            exp_f := 1;
        ELSIF x =- 14940 THEN
            exp_f := 1;
        ELSIF x =- 14939 THEN
            exp_f := 1;
        ELSIF x =- 14938 THEN
            exp_f := 1;
        ELSIF x =- 14937 THEN
            exp_f := 1;
        ELSIF x =- 14936 THEN
            exp_f := 1;
        ELSIF x =- 14935 THEN
            exp_f := 1;
        ELSIF x =- 14934 THEN
            exp_f := 1;
        ELSIF x =- 14933 THEN
            exp_f := 1;
        ELSIF x =- 14932 THEN
            exp_f := 1;
        ELSIF x =- 14931 THEN
            exp_f := 1;
        ELSIF x =- 14930 THEN
            exp_f := 1;
        ELSIF x =- 14929 THEN
            exp_f := 1;
        ELSIF x =- 14928 THEN
            exp_f := 1;
        ELSIF x =- 14927 THEN
            exp_f := 1;
        ELSIF x =- 14926 THEN
            exp_f := 1;
        ELSIF x =- 14925 THEN
            exp_f := 1;
        ELSIF x =- 14924 THEN
            exp_f := 1;
        ELSIF x =- 14923 THEN
            exp_f := 1;
        ELSIF x =- 14922 THEN
            exp_f := 1;
        ELSIF x =- 14921 THEN
            exp_f := 1;
        ELSIF x =- 14920 THEN
            exp_f := 1;
        ELSIF x =- 14919 THEN
            exp_f := 1;
        ELSIF x =- 14918 THEN
            exp_f := 1;
        ELSIF x =- 14917 THEN
            exp_f := 1;
        ELSIF x =- 14916 THEN
            exp_f := 1;
        ELSIF x =- 14915 THEN
            exp_f := 1;
        ELSIF x =- 14914 THEN
            exp_f := 1;
        ELSIF x =- 14913 THEN
            exp_f := 1;
        ELSIF x =- 14912 THEN
            exp_f := 1;
        ELSIF x =- 14911 THEN
            exp_f := 1;
        ELSIF x =- 14910 THEN
            exp_f := 1;
        ELSIF x =- 14909 THEN
            exp_f := 1;
        ELSIF x =- 14908 THEN
            exp_f := 1;
        ELSIF x =- 14907 THEN
            exp_f := 1;
        ELSIF x =- 14906 THEN
            exp_f := 1;
        ELSIF x =- 14905 THEN
            exp_f := 1;
        ELSIF x =- 14904 THEN
            exp_f := 1;
        ELSIF x =- 14903 THEN
            exp_f := 1;
        ELSIF x =- 14902 THEN
            exp_f := 1;
        ELSIF x =- 14901 THEN
            exp_f := 1;
        ELSIF x =- 14900 THEN
            exp_f := 1;
        ELSIF x =- 14899 THEN
            exp_f := 1;
        ELSIF x =- 14898 THEN
            exp_f := 1;
        ELSIF x =- 14897 THEN
            exp_f := 1;
        ELSIF x =- 14896 THEN
            exp_f := 1;
        ELSIF x =- 14895 THEN
            exp_f := 1;
        ELSIF x =- 14894 THEN
            exp_f := 1;
        ELSIF x =- 14893 THEN
            exp_f := 1;
        ELSIF x =- 14892 THEN
            exp_f := 1;
        ELSIF x =- 14891 THEN
            exp_f := 1;
        ELSIF x =- 14890 THEN
            exp_f := 1;
        ELSIF x =- 14889 THEN
            exp_f := 1;
        ELSIF x =- 14888 THEN
            exp_f := 1;
        ELSIF x =- 14887 THEN
            exp_f := 1;
        ELSIF x =- 14886 THEN
            exp_f := 1;
        ELSIF x =- 14885 THEN
            exp_f := 1;
        ELSIF x =- 14884 THEN
            exp_f := 1;
        ELSIF x =- 14883 THEN
            exp_f := 1;
        ELSIF x =- 14882 THEN
            exp_f := 1;
        ELSIF x =- 14881 THEN
            exp_f := 1;
        ELSIF x =- 14880 THEN
            exp_f := 1;
        ELSIF x =- 14879 THEN
            exp_f := 1;
        ELSIF x =- 14878 THEN
            exp_f := 1;
        ELSIF x =- 14877 THEN
            exp_f := 1;
        ELSIF x =- 14876 THEN
            exp_f := 1;
        ELSIF x =- 14875 THEN
            exp_f := 1;
        ELSIF x =- 14874 THEN
            exp_f := 1;
        ELSIF x =- 14873 THEN
            exp_f := 1;
        ELSIF x =- 14872 THEN
            exp_f := 1;
        ELSIF x =- 14871 THEN
            exp_f := 1;
        ELSIF x =- 14870 THEN
            exp_f := 1;
        ELSIF x =- 14869 THEN
            exp_f := 1;
        ELSIF x =- 14868 THEN
            exp_f := 1;
        ELSIF x =- 14867 THEN
            exp_f := 1;
        ELSIF x =- 14866 THEN
            exp_f := 1;
        ELSIF x =- 14865 THEN
            exp_f := 1;
        ELSIF x =- 14864 THEN
            exp_f := 1;
        ELSIF x =- 14863 THEN
            exp_f := 1;
        ELSIF x =- 14862 THEN
            exp_f := 1;
        ELSIF x =- 14861 THEN
            exp_f := 1;
        ELSIF x =- 14860 THEN
            exp_f := 1;
        ELSIF x =- 14859 THEN
            exp_f := 1;
        ELSIF x =- 14858 THEN
            exp_f := 1;
        ELSIF x =- 14857 THEN
            exp_f := 1;
        ELSIF x =- 14856 THEN
            exp_f := 1;
        ELSIF x =- 14855 THEN
            exp_f := 1;
        ELSIF x =- 14854 THEN
            exp_f := 1;
        ELSIF x =- 14853 THEN
            exp_f := 1;
        ELSIF x =- 14852 THEN
            exp_f := 1;
        ELSIF x =- 14851 THEN
            exp_f := 1;
        ELSIF x =- 14850 THEN
            exp_f := 1;
        ELSIF x =- 14849 THEN
            exp_f := 1;
        ELSIF x =- 14848 THEN
            exp_f := 1;
        ELSIF x =- 14847 THEN
            exp_f := 2;
        ELSIF x =- 14846 THEN
            exp_f := 2;
        ELSIF x =- 14845 THEN
            exp_f := 2;
        ELSIF x =- 14844 THEN
            exp_f := 2;
        ELSIF x =- 14843 THEN
            exp_f := 2;
        ELSIF x =- 14842 THEN
            exp_f := 2;
        ELSIF x =- 14841 THEN
            exp_f := 2;
        ELSIF x =- 14840 THEN
            exp_f := 2;
        ELSIF x =- 14839 THEN
            exp_f := 2;
        ELSIF x =- 14838 THEN
            exp_f := 2;
        ELSIF x =- 14837 THEN
            exp_f := 2;
        ELSIF x =- 14836 THEN
            exp_f := 2;
        ELSIF x =- 14835 THEN
            exp_f := 2;
        ELSIF x =- 14834 THEN
            exp_f := 2;
        ELSIF x =- 14833 THEN
            exp_f := 2;
        ELSIF x =- 14832 THEN
            exp_f := 2;
        ELSIF x =- 14831 THEN
            exp_f := 2;
        ELSIF x =- 14830 THEN
            exp_f := 2;
        ELSIF x =- 14829 THEN
            exp_f := 2;
        ELSIF x =- 14828 THEN
            exp_f := 2;
        ELSIF x =- 14827 THEN
            exp_f := 2;
        ELSIF x =- 14826 THEN
            exp_f := 2;
        ELSIF x =- 14825 THEN
            exp_f := 2;
        ELSIF x =- 14824 THEN
            exp_f := 2;
        ELSIF x =- 14823 THEN
            exp_f := 2;
        ELSIF x =- 14822 THEN
            exp_f := 2;
        ELSIF x =- 14821 THEN
            exp_f := 2;
        ELSIF x =- 14820 THEN
            exp_f := 2;
        ELSIF x =- 14819 THEN
            exp_f := 2;
        ELSIF x =- 14818 THEN
            exp_f := 2;
        ELSIF x =- 14817 THEN
            exp_f := 2;
        ELSIF x =- 14816 THEN
            exp_f := 2;
        ELSIF x =- 14815 THEN
            exp_f := 2;
        ELSIF x =- 14814 THEN
            exp_f := 2;
        ELSIF x =- 14813 THEN
            exp_f := 2;
        ELSIF x =- 14812 THEN
            exp_f := 2;
        ELSIF x =- 14811 THEN
            exp_f := 2;
        ELSIF x =- 14810 THEN
            exp_f := 2;
        ELSIF x =- 14809 THEN
            exp_f := 2;
        ELSIF x =- 14808 THEN
            exp_f := 2;
        ELSIF x =- 14807 THEN
            exp_f := 2;
        ELSIF x =- 14806 THEN
            exp_f := 2;
        ELSIF x =- 14805 THEN
            exp_f := 2;
        ELSIF x =- 14804 THEN
            exp_f := 2;
        ELSIF x =- 14803 THEN
            exp_f := 2;
        ELSIF x =- 14802 THEN
            exp_f := 2;
        ELSIF x =- 14801 THEN
            exp_f := 2;
        ELSIF x =- 14800 THEN
            exp_f := 2;
        ELSIF x =- 14799 THEN
            exp_f := 2;
        ELSIF x =- 14798 THEN
            exp_f := 2;
        ELSIF x =- 14797 THEN
            exp_f := 2;
        ELSIF x =- 14796 THEN
            exp_f := 2;
        ELSIF x =- 14795 THEN
            exp_f := 2;
        ELSIF x =- 14794 THEN
            exp_f := 2;
        ELSIF x =- 14793 THEN
            exp_f := 2;
        ELSIF x =- 14792 THEN
            exp_f := 2;
        ELSIF x =- 14791 THEN
            exp_f := 2;
        ELSIF x =- 14790 THEN
            exp_f := 2;
        ELSIF x =- 14789 THEN
            exp_f := 2;
        ELSIF x =- 14788 THEN
            exp_f := 2;
        ELSIF x =- 14787 THEN
            exp_f := 2;
        ELSIF x =- 14786 THEN
            exp_f := 2;
        ELSIF x =- 14785 THEN
            exp_f := 2;
        ELSIF x =- 14784 THEN
            exp_f := 2;
        ELSIF x =- 14783 THEN
            exp_f := 2;
        ELSIF x =- 14782 THEN
            exp_f := 2;
        ELSIF x =- 14781 THEN
            exp_f := 2;
        ELSIF x =- 14780 THEN
            exp_f := 2;
        ELSIF x =- 14779 THEN
            exp_f := 2;
        ELSIF x =- 14778 THEN
            exp_f := 2;
        ELSIF x =- 14777 THEN
            exp_f := 2;
        ELSIF x =- 14776 THEN
            exp_f := 2;
        ELSIF x =- 14775 THEN
            exp_f := 2;
        ELSIF x =- 14774 THEN
            exp_f := 2;
        ELSIF x =- 14773 THEN
            exp_f := 2;
        ELSIF x =- 14772 THEN
            exp_f := 2;
        ELSIF x =- 14771 THEN
            exp_f := 2;
        ELSIF x =- 14770 THEN
            exp_f := 2;
        ELSIF x =- 14769 THEN
            exp_f := 2;
        ELSIF x =- 14768 THEN
            exp_f := 2;
        ELSIF x =- 14767 THEN
            exp_f := 2;
        ELSIF x =- 14766 THEN
            exp_f := 2;
        ELSIF x =- 14765 THEN
            exp_f := 2;
        ELSIF x =- 14764 THEN
            exp_f := 2;
        ELSIF x =- 14763 THEN
            exp_f := 2;
        ELSIF x =- 14762 THEN
            exp_f := 2;
        ELSIF x =- 14761 THEN
            exp_f := 2;
        ELSIF x =- 14760 THEN
            exp_f := 2;
        ELSIF x =- 14759 THEN
            exp_f := 2;
        ELSIF x =- 14758 THEN
            exp_f := 2;
        ELSIF x =- 14757 THEN
            exp_f := 2;
        ELSIF x =- 14756 THEN
            exp_f := 2;
        ELSIF x =- 14755 THEN
            exp_f := 2;
        ELSIF x =- 14754 THEN
            exp_f := 2;
        ELSIF x =- 14753 THEN
            exp_f := 2;
        ELSIF x =- 14752 THEN
            exp_f := 2;
        ELSIF x =- 14751 THEN
            exp_f := 2;
        ELSIF x =- 14750 THEN
            exp_f := 2;
        ELSIF x =- 14749 THEN
            exp_f := 2;
        ELSIF x =- 14748 THEN
            exp_f := 2;
        ELSIF x =- 14747 THEN
            exp_f := 2;
        ELSIF x =- 14746 THEN
            exp_f := 2;
        ELSIF x =- 14745 THEN
            exp_f := 2;
        ELSIF x =- 14744 THEN
            exp_f := 2;
        ELSIF x =- 14743 THEN
            exp_f := 2;
        ELSIF x =- 14742 THEN
            exp_f := 2;
        ELSIF x =- 14741 THEN
            exp_f := 2;
        ELSIF x =- 14740 THEN
            exp_f := 2;
        ELSIF x =- 14739 THEN
            exp_f := 2;
        ELSIF x =- 14738 THEN
            exp_f := 2;
        ELSIF x =- 14737 THEN
            exp_f := 2;
        ELSIF x =- 14736 THEN
            exp_f := 2;
        ELSIF x =- 14735 THEN
            exp_f := 2;
        ELSIF x =- 14734 THEN
            exp_f := 2;
        ELSIF x =- 14733 THEN
            exp_f := 2;
        ELSIF x =- 14732 THEN
            exp_f := 2;
        ELSIF x =- 14731 THEN
            exp_f := 2;
        ELSIF x =- 14730 THEN
            exp_f := 2;
        ELSIF x =- 14729 THEN
            exp_f := 2;
        ELSIF x =- 14728 THEN
            exp_f := 2;
        ELSIF x =- 14727 THEN
            exp_f := 2;
        ELSIF x =- 14726 THEN
            exp_f := 2;
        ELSIF x =- 14725 THEN
            exp_f := 2;
        ELSIF x =- 14724 THEN
            exp_f := 2;
        ELSIF x =- 14723 THEN
            exp_f := 2;
        ELSIF x =- 14722 THEN
            exp_f := 2;
        ELSIF x =- 14721 THEN
            exp_f := 2;
        ELSIF x =- 14720 THEN
            exp_f := 2;
        ELSIF x =- 14719 THEN
            exp_f := 2;
        ELSIF x =- 14718 THEN
            exp_f := 2;
        ELSIF x =- 14717 THEN
            exp_f := 2;
        ELSIF x =- 14716 THEN
            exp_f := 2;
        ELSIF x =- 14715 THEN
            exp_f := 2;
        ELSIF x =- 14714 THEN
            exp_f := 2;
        ELSIF x =- 14713 THEN
            exp_f := 2;
        ELSIF x =- 14712 THEN
            exp_f := 2;
        ELSIF x =- 14711 THEN
            exp_f := 2;
        ELSIF x =- 14710 THEN
            exp_f := 2;
        ELSIF x =- 14709 THEN
            exp_f := 2;
        ELSIF x =- 14708 THEN
            exp_f := 2;
        ELSIF x =- 14707 THEN
            exp_f := 2;
        ELSIF x =- 14706 THEN
            exp_f := 2;
        ELSIF x =- 14705 THEN
            exp_f := 2;
        ELSIF x =- 14704 THEN
            exp_f := 2;
        ELSIF x =- 14703 THEN
            exp_f := 2;
        ELSIF x =- 14702 THEN
            exp_f := 2;
        ELSIF x =- 14701 THEN
            exp_f := 2;
        ELSIF x =- 14700 THEN
            exp_f := 2;
        ELSIF x =- 14699 THEN
            exp_f := 2;
        ELSIF x =- 14698 THEN
            exp_f := 2;
        ELSIF x =- 14697 THEN
            exp_f := 2;
        ELSIF x =- 14696 THEN
            exp_f := 2;
        ELSIF x =- 14695 THEN
            exp_f := 2;
        ELSIF x =- 14694 THEN
            exp_f := 2;
        ELSIF x =- 14693 THEN
            exp_f := 2;
        ELSIF x =- 14692 THEN
            exp_f := 2;
        ELSIF x =- 14691 THEN
            exp_f := 2;
        ELSIF x =- 14690 THEN
            exp_f := 2;
        ELSIF x =- 14689 THEN
            exp_f := 2;
        ELSIF x =- 14688 THEN
            exp_f := 2;
        ELSIF x =- 14687 THEN
            exp_f := 2;
        ELSIF x =- 14686 THEN
            exp_f := 2;
        ELSIF x =- 14685 THEN
            exp_f := 2;
        ELSIF x =- 14684 THEN
            exp_f := 2;
        ELSIF x =- 14683 THEN
            exp_f := 2;
        ELSIF x =- 14682 THEN
            exp_f := 2;
        ELSIF x =- 14681 THEN
            exp_f := 2;
        ELSIF x =- 14680 THEN
            exp_f := 2;
        ELSIF x =- 14679 THEN
            exp_f := 2;
        ELSIF x =- 14678 THEN
            exp_f := 2;
        ELSIF x =- 14677 THEN
            exp_f := 2;
        ELSIF x =- 14676 THEN
            exp_f := 2;
        ELSIF x =- 14675 THEN
            exp_f := 2;
        ELSIF x =- 14674 THEN
            exp_f := 2;
        ELSIF x =- 14673 THEN
            exp_f := 2;
        ELSIF x =- 14672 THEN
            exp_f := 2;
        ELSIF x =- 14671 THEN
            exp_f := 2;
        ELSIF x =- 14670 THEN
            exp_f := 2;
        ELSIF x =- 14669 THEN
            exp_f := 2;
        ELSIF x =- 14668 THEN
            exp_f := 2;
        ELSIF x =- 14667 THEN
            exp_f := 2;
        ELSIF x =- 14666 THEN
            exp_f := 2;
        ELSIF x =- 14665 THEN
            exp_f := 2;
        ELSIF x =- 14664 THEN
            exp_f := 2;
        ELSIF x =- 14663 THEN
            exp_f := 2;
        ELSIF x =- 14662 THEN
            exp_f := 2;
        ELSIF x =- 14661 THEN
            exp_f := 2;
        ELSIF x =- 14660 THEN
            exp_f := 2;
        ELSIF x =- 14659 THEN
            exp_f := 2;
        ELSIF x =- 14658 THEN
            exp_f := 2;
        ELSIF x =- 14657 THEN
            exp_f := 2;
        ELSIF x =- 14656 THEN
            exp_f := 2;
        ELSIF x =- 14655 THEN
            exp_f := 2;
        ELSIF x =- 14654 THEN
            exp_f := 2;
        ELSIF x =- 14653 THEN
            exp_f := 2;
        ELSIF x =- 14652 THEN
            exp_f := 2;
        ELSIF x =- 14651 THEN
            exp_f := 2;
        ELSIF x =- 14650 THEN
            exp_f := 2;
        ELSIF x =- 14649 THEN
            exp_f := 2;
        ELSIF x =- 14648 THEN
            exp_f := 2;
        ELSIF x =- 14647 THEN
            exp_f := 2;
        ELSIF x =- 14646 THEN
            exp_f := 2;
        ELSIF x =- 14645 THEN
            exp_f := 2;
        ELSIF x =- 14644 THEN
            exp_f := 2;
        ELSIF x =- 14643 THEN
            exp_f := 2;
        ELSIF x =- 14642 THEN
            exp_f := 2;
        ELSIF x =- 14641 THEN
            exp_f := 2;
        ELSIF x =- 14640 THEN
            exp_f := 2;
        ELSIF x =- 14639 THEN
            exp_f := 2;
        ELSIF x =- 14638 THEN
            exp_f := 2;
        ELSIF x =- 14637 THEN
            exp_f := 2;
        ELSIF x =- 14636 THEN
            exp_f := 2;
        ELSIF x =- 14635 THEN
            exp_f := 2;
        ELSIF x =- 14634 THEN
            exp_f := 2;
        ELSIF x =- 14633 THEN
            exp_f := 2;
        ELSIF x =- 14632 THEN
            exp_f := 2;
        ELSIF x =- 14631 THEN
            exp_f := 2;
        ELSIF x =- 14630 THEN
            exp_f := 2;
        ELSIF x =- 14629 THEN
            exp_f := 2;
        ELSIF x =- 14628 THEN
            exp_f := 2;
        ELSIF x =- 14627 THEN
            exp_f := 2;
        ELSIF x =- 14626 THEN
            exp_f := 2;
        ELSIF x =- 14625 THEN
            exp_f := 2;
        ELSIF x =- 14624 THEN
            exp_f := 2;
        ELSIF x =- 14623 THEN
            exp_f := 2;
        ELSIF x =- 14622 THEN
            exp_f := 2;
        ELSIF x =- 14621 THEN
            exp_f := 2;
        ELSIF x =- 14620 THEN
            exp_f := 2;
        ELSIF x =- 14619 THEN
            exp_f := 2;
        ELSIF x =- 14618 THEN
            exp_f := 2;
        ELSIF x =- 14617 THEN
            exp_f := 2;
        ELSIF x =- 14616 THEN
            exp_f := 2;
        ELSIF x =- 14615 THEN
            exp_f := 2;
        ELSIF x =- 14614 THEN
            exp_f := 2;
        ELSIF x =- 14613 THEN
            exp_f := 2;
        ELSIF x =- 14612 THEN
            exp_f := 2;
        ELSIF x =- 14611 THEN
            exp_f := 2;
        ELSIF x =- 14610 THEN
            exp_f := 2;
        ELSIF x =- 14609 THEN
            exp_f := 2;
        ELSIF x =- 14608 THEN
            exp_f := 2;
        ELSIF x =- 14607 THEN
            exp_f := 2;
        ELSIF x =- 14606 THEN
            exp_f := 2;
        ELSIF x =- 14605 THEN
            exp_f := 2;
        ELSIF x =- 14604 THEN
            exp_f := 2;
        ELSIF x =- 14603 THEN
            exp_f := 2;
        ELSIF x =- 14602 THEN
            exp_f := 2;
        ELSIF x =- 14601 THEN
            exp_f := 2;
        ELSIF x =- 14600 THEN
            exp_f := 2;
        ELSIF x =- 14599 THEN
            exp_f := 2;
        ELSIF x =- 14598 THEN
            exp_f := 2;
        ELSIF x =- 14597 THEN
            exp_f := 2;
        ELSIF x =- 14596 THEN
            exp_f := 2;
        ELSIF x =- 14595 THEN
            exp_f := 2;
        ELSIF x =- 14594 THEN
            exp_f := 2;
        ELSIF x =- 14593 THEN
            exp_f := 2;
        ELSIF x =- 14592 THEN
            exp_f := 2;
        ELSIF x =- 14591 THEN
            exp_f := 2;
        ELSIF x =- 14590 THEN
            exp_f := 2;
        ELSIF x =- 14589 THEN
            exp_f := 2;
        ELSIF x =- 14588 THEN
            exp_f := 2;
        ELSIF x =- 14587 THEN
            exp_f := 2;
        ELSIF x =- 14586 THEN
            exp_f := 2;
        ELSIF x =- 14585 THEN
            exp_f := 2;
        ELSIF x =- 14584 THEN
            exp_f := 2;
        ELSIF x =- 14583 THEN
            exp_f := 2;
        ELSIF x =- 14582 THEN
            exp_f := 2;
        ELSIF x =- 14581 THEN
            exp_f := 2;
        ELSIF x =- 14580 THEN
            exp_f := 2;
        ELSIF x =- 14579 THEN
            exp_f := 2;
        ELSIF x =- 14578 THEN
            exp_f := 2;
        ELSIF x =- 14577 THEN
            exp_f := 2;
        ELSIF x =- 14576 THEN
            exp_f := 2;
        ELSIF x =- 14575 THEN
            exp_f := 2;
        ELSIF x =- 14574 THEN
            exp_f := 2;
        ELSIF x =- 14573 THEN
            exp_f := 2;
        ELSIF x =- 14572 THEN
            exp_f := 2;
        ELSIF x =- 14571 THEN
            exp_f := 2;
        ELSIF x =- 14570 THEN
            exp_f := 2;
        ELSIF x =- 14569 THEN
            exp_f := 2;
        ELSIF x =- 14568 THEN
            exp_f := 2;
        ELSIF x =- 14567 THEN
            exp_f := 2;
        ELSIF x =- 14566 THEN
            exp_f := 2;
        ELSIF x =- 14565 THEN
            exp_f := 2;
        ELSIF x =- 14564 THEN
            exp_f := 2;
        ELSIF x =- 14563 THEN
            exp_f := 2;
        ELSIF x =- 14562 THEN
            exp_f := 2;
        ELSIF x =- 14561 THEN
            exp_f := 2;
        ELSIF x =- 14560 THEN
            exp_f := 2;
        ELSIF x =- 14559 THEN
            exp_f := 2;
        ELSIF x =- 14558 THEN
            exp_f := 2;
        ELSIF x =- 14557 THEN
            exp_f := 2;
        ELSIF x =- 14556 THEN
            exp_f := 2;
        ELSIF x =- 14555 THEN
            exp_f := 2;
        ELSIF x =- 14554 THEN
            exp_f := 2;
        ELSIF x =- 14553 THEN
            exp_f := 2;
        ELSIF x =- 14552 THEN
            exp_f := 2;
        ELSIF x =- 14551 THEN
            exp_f := 2;
        ELSIF x =- 14550 THEN
            exp_f := 2;
        ELSIF x =- 14549 THEN
            exp_f := 2;
        ELSIF x =- 14548 THEN
            exp_f := 2;
        ELSIF x =- 14547 THEN
            exp_f := 2;
        ELSIF x =- 14546 THEN
            exp_f := 2;
        ELSIF x =- 14545 THEN
            exp_f := 2;
        ELSIF x =- 14544 THEN
            exp_f := 2;
        ELSIF x =- 14543 THEN
            exp_f := 2;
        ELSIF x =- 14542 THEN
            exp_f := 2;
        ELSIF x =- 14541 THEN
            exp_f := 2;
        ELSIF x =- 14540 THEN
            exp_f := 2;
        ELSIF x =- 14539 THEN
            exp_f := 2;
        ELSIF x =- 14538 THEN
            exp_f := 2;
        ELSIF x =- 14537 THEN
            exp_f := 2;
        ELSIF x =- 14536 THEN
            exp_f := 2;
        ELSIF x =- 14535 THEN
            exp_f := 2;
        ELSIF x =- 14534 THEN
            exp_f := 2;
        ELSIF x =- 14533 THEN
            exp_f := 2;
        ELSIF x =- 14532 THEN
            exp_f := 2;
        ELSIF x =- 14531 THEN
            exp_f := 2;
        ELSIF x =- 14530 THEN
            exp_f := 2;
        ELSIF x =- 14529 THEN
            exp_f := 2;
        ELSIF x =- 14528 THEN
            exp_f := 2;
        ELSIF x =- 14527 THEN
            exp_f := 2;
        ELSIF x =- 14526 THEN
            exp_f := 2;
        ELSIF x =- 14525 THEN
            exp_f := 2;
        ELSIF x =- 14524 THEN
            exp_f := 2;
        ELSIF x =- 14523 THEN
            exp_f := 2;
        ELSIF x =- 14522 THEN
            exp_f := 2;
        ELSIF x =- 14521 THEN
            exp_f := 2;
        ELSIF x =- 14520 THEN
            exp_f := 2;
        ELSIF x =- 14519 THEN
            exp_f := 2;
        ELSIF x =- 14518 THEN
            exp_f := 2;
        ELSIF x =- 14517 THEN
            exp_f := 2;
        ELSIF x =- 14516 THEN
            exp_f := 2;
        ELSIF x =- 14515 THEN
            exp_f := 2;
        ELSIF x =- 14514 THEN
            exp_f := 2;
        ELSIF x =- 14513 THEN
            exp_f := 2;
        ELSIF x =- 14512 THEN
            exp_f := 2;
        ELSIF x =- 14511 THEN
            exp_f := 2;
        ELSIF x =- 14510 THEN
            exp_f := 2;
        ELSIF x =- 14509 THEN
            exp_f := 2;
        ELSIF x =- 14508 THEN
            exp_f := 2;
        ELSIF x =- 14507 THEN
            exp_f := 2;
        ELSIF x =- 14506 THEN
            exp_f := 2;
        ELSIF x =- 14505 THEN
            exp_f := 2;
        ELSIF x =- 14504 THEN
            exp_f := 2;
        ELSIF x =- 14503 THEN
            exp_f := 2;
        ELSIF x =- 14502 THEN
            exp_f := 2;
        ELSIF x =- 14501 THEN
            exp_f := 2;
        ELSIF x =- 14500 THEN
            exp_f := 2;
        ELSIF x =- 14499 THEN
            exp_f := 2;
        ELSIF x =- 14498 THEN
            exp_f := 2;
        ELSIF x =- 14497 THEN
            exp_f := 2;
        ELSIF x =- 14496 THEN
            exp_f := 2;
        ELSIF x =- 14495 THEN
            exp_f := 2;
        ELSIF x =- 14494 THEN
            exp_f := 2;
        ELSIF x =- 14493 THEN
            exp_f := 2;
        ELSIF x =- 14492 THEN
            exp_f := 2;
        ELSIF x =- 14491 THEN
            exp_f := 2;
        ELSIF x =- 14490 THEN
            exp_f := 2;
        ELSIF x =- 14489 THEN
            exp_f := 2;
        ELSIF x =- 14488 THEN
            exp_f := 2;
        ELSIF x =- 14487 THEN
            exp_f := 2;
        ELSIF x =- 14486 THEN
            exp_f := 2;
        ELSIF x =- 14485 THEN
            exp_f := 2;
        ELSIF x =- 14484 THEN
            exp_f := 2;
        ELSIF x =- 14483 THEN
            exp_f := 2;
        ELSIF x =- 14482 THEN
            exp_f := 2;
        ELSIF x =- 14481 THEN
            exp_f := 2;
        ELSIF x =- 14480 THEN
            exp_f := 2;
        ELSIF x =- 14479 THEN
            exp_f := 2;
        ELSIF x =- 14478 THEN
            exp_f := 2;
        ELSIF x =- 14477 THEN
            exp_f := 2;
        ELSIF x =- 14476 THEN
            exp_f := 2;
        ELSIF x =- 14475 THEN
            exp_f := 2;
        ELSIF x =- 14474 THEN
            exp_f := 2;
        ELSIF x =- 14473 THEN
            exp_f := 2;
        ELSIF x =- 14472 THEN
            exp_f := 2;
        ELSIF x =- 14471 THEN
            exp_f := 2;
        ELSIF x =- 14470 THEN
            exp_f := 2;
        ELSIF x =- 14469 THEN
            exp_f := 2;
        ELSIF x =- 14468 THEN
            exp_f := 2;
        ELSIF x =- 14467 THEN
            exp_f := 2;
        ELSIF x =- 14466 THEN
            exp_f := 2;
        ELSIF x =- 14465 THEN
            exp_f := 2;
        ELSIF x =- 14464 THEN
            exp_f := 2;
        ELSIF x =- 14463 THEN
            exp_f := 2;
        ELSIF x =- 14462 THEN
            exp_f := 2;
        ELSIF x =- 14461 THEN
            exp_f := 2;
        ELSIF x =- 14460 THEN
            exp_f := 2;
        ELSIF x =- 14459 THEN
            exp_f := 2;
        ELSIF x =- 14458 THEN
            exp_f := 2;
        ELSIF x =- 14457 THEN
            exp_f := 2;
        ELSIF x =- 14456 THEN
            exp_f := 2;
        ELSIF x =- 14455 THEN
            exp_f := 2;
        ELSIF x =- 14454 THEN
            exp_f := 2;
        ELSIF x =- 14453 THEN
            exp_f := 2;
        ELSIF x =- 14452 THEN
            exp_f := 2;
        ELSIF x =- 14451 THEN
            exp_f := 2;
        ELSIF x =- 14450 THEN
            exp_f := 2;
        ELSIF x =- 14449 THEN
            exp_f := 2;
        ELSIF x =- 14448 THEN
            exp_f := 2;
        ELSIF x =- 14447 THEN
            exp_f := 2;
        ELSIF x =- 14446 THEN
            exp_f := 2;
        ELSIF x =- 14445 THEN
            exp_f := 2;
        ELSIF x =- 14444 THEN
            exp_f := 2;
        ELSIF x =- 14443 THEN
            exp_f := 2;
        ELSIF x =- 14442 THEN
            exp_f := 2;
        ELSIF x =- 14441 THEN
            exp_f := 2;
        ELSIF x =- 14440 THEN
            exp_f := 2;
        ELSIF x =- 14439 THEN
            exp_f := 2;
        ELSIF x =- 14438 THEN
            exp_f := 2;
        ELSIF x =- 14437 THEN
            exp_f := 2;
        ELSIF x =- 14436 THEN
            exp_f := 2;
        ELSIF x =- 14435 THEN
            exp_f := 2;
        ELSIF x =- 14434 THEN
            exp_f := 2;
        ELSIF x =- 14433 THEN
            exp_f := 2;
        ELSIF x =- 14432 THEN
            exp_f := 2;
        ELSIF x =- 14431 THEN
            exp_f := 2;
        ELSIF x =- 14430 THEN
            exp_f := 2;
        ELSIF x =- 14429 THEN
            exp_f := 2;
        ELSIF x =- 14428 THEN
            exp_f := 2;
        ELSIF x =- 14427 THEN
            exp_f := 2;
        ELSIF x =- 14426 THEN
            exp_f := 2;
        ELSIF x =- 14425 THEN
            exp_f := 2;
        ELSIF x =- 14424 THEN
            exp_f := 2;
        ELSIF x =- 14423 THEN
            exp_f := 2;
        ELSIF x =- 14422 THEN
            exp_f := 2;
        ELSIF x =- 14421 THEN
            exp_f := 2;
        ELSIF x =- 14420 THEN
            exp_f := 2;
        ELSIF x =- 14419 THEN
            exp_f := 2;
        ELSIF x =- 14418 THEN
            exp_f := 2;
        ELSIF x =- 14417 THEN
            exp_f := 2;
        ELSIF x =- 14416 THEN
            exp_f := 2;
        ELSIF x =- 14415 THEN
            exp_f := 2;
        ELSIF x =- 14414 THEN
            exp_f := 2;
        ELSIF x =- 14413 THEN
            exp_f := 2;
        ELSIF x =- 14412 THEN
            exp_f := 2;
        ELSIF x =- 14411 THEN
            exp_f := 2;
        ELSIF x =- 14410 THEN
            exp_f := 2;
        ELSIF x =- 14409 THEN
            exp_f := 2;
        ELSIF x =- 14408 THEN
            exp_f := 2;
        ELSIF x =- 14407 THEN
            exp_f := 2;
        ELSIF x =- 14406 THEN
            exp_f := 2;
        ELSIF x =- 14405 THEN
            exp_f := 2;
        ELSIF x =- 14404 THEN
            exp_f := 2;
        ELSIF x =- 14403 THEN
            exp_f := 2;
        ELSIF x =- 14402 THEN
            exp_f := 2;
        ELSIF x =- 14401 THEN
            exp_f := 2;
        ELSIF x =- 14400 THEN
            exp_f := 2;
        ELSIF x =- 14399 THEN
            exp_f := 2;
        ELSIF x =- 14398 THEN
            exp_f := 2;
        ELSIF x =- 14397 THEN
            exp_f := 2;
        ELSIF x =- 14396 THEN
            exp_f := 2;
        ELSIF x =- 14395 THEN
            exp_f := 2;
        ELSIF x =- 14394 THEN
            exp_f := 2;
        ELSIF x =- 14393 THEN
            exp_f := 2;
        ELSIF x =- 14392 THEN
            exp_f := 2;
        ELSIF x =- 14391 THEN
            exp_f := 2;
        ELSIF x =- 14390 THEN
            exp_f := 2;
        ELSIF x =- 14389 THEN
            exp_f := 2;
        ELSIF x =- 14388 THEN
            exp_f := 2;
        ELSIF x =- 14387 THEN
            exp_f := 2;
        ELSIF x =- 14386 THEN
            exp_f := 2;
        ELSIF x =- 14385 THEN
            exp_f := 2;
        ELSIF x =- 14384 THEN
            exp_f := 2;
        ELSIF x =- 14383 THEN
            exp_f := 2;
        ELSIF x =- 14382 THEN
            exp_f := 2;
        ELSIF x =- 14381 THEN
            exp_f := 2;
        ELSIF x =- 14380 THEN
            exp_f := 2;
        ELSIF x =- 14379 THEN
            exp_f := 2;
        ELSIF x =- 14378 THEN
            exp_f := 2;
        ELSIF x =- 14377 THEN
            exp_f := 2;
        ELSIF x =- 14376 THEN
            exp_f := 2;
        ELSIF x =- 14375 THEN
            exp_f := 2;
        ELSIF x =- 14374 THEN
            exp_f := 2;
        ELSIF x =- 14373 THEN
            exp_f := 2;
        ELSIF x =- 14372 THEN
            exp_f := 2;
        ELSIF x =- 14371 THEN
            exp_f := 2;
        ELSIF x =- 14370 THEN
            exp_f := 2;
        ELSIF x =- 14369 THEN
            exp_f := 2;
        ELSIF x =- 14368 THEN
            exp_f := 2;
        ELSIF x =- 14367 THEN
            exp_f := 2;
        ELSIF x =- 14366 THEN
            exp_f := 2;
        ELSIF x =- 14365 THEN
            exp_f := 2;
        ELSIF x =- 14364 THEN
            exp_f := 2;
        ELSIF x =- 14363 THEN
            exp_f := 2;
        ELSIF x =- 14362 THEN
            exp_f := 2;
        ELSIF x =- 14361 THEN
            exp_f := 2;
        ELSIF x =- 14360 THEN
            exp_f := 2;
        ELSIF x =- 14359 THEN
            exp_f := 2;
        ELSIF x =- 14358 THEN
            exp_f := 2;
        ELSIF x =- 14357 THEN
            exp_f := 2;
        ELSIF x =- 14356 THEN
            exp_f := 2;
        ELSIF x =- 14355 THEN
            exp_f := 2;
        ELSIF x =- 14354 THEN
            exp_f := 2;
        ELSIF x =- 14353 THEN
            exp_f := 2;
        ELSIF x =- 14352 THEN
            exp_f := 2;
        ELSIF x =- 14351 THEN
            exp_f := 2;
        ELSIF x =- 14350 THEN
            exp_f := 2;
        ELSIF x =- 14349 THEN
            exp_f := 2;
        ELSIF x =- 14348 THEN
            exp_f := 2;
        ELSIF x =- 14347 THEN
            exp_f := 2;
        ELSIF x =- 14346 THEN
            exp_f := 2;
        ELSIF x =- 14345 THEN
            exp_f := 2;
        ELSIF x =- 14344 THEN
            exp_f := 2;
        ELSIF x =- 14343 THEN
            exp_f := 2;
        ELSIF x =- 14342 THEN
            exp_f := 2;
        ELSIF x =- 14341 THEN
            exp_f := 2;
        ELSIF x =- 14340 THEN
            exp_f := 2;
        ELSIF x =- 14339 THEN
            exp_f := 2;
        ELSIF x =- 14338 THEN
            exp_f := 2;
        ELSIF x =- 14337 THEN
            exp_f := 2;
        ELSIF x =- 14336 THEN
            exp_f := 2;
        ELSIF x =- 14335 THEN
            exp_f := 2;
        ELSIF x =- 14334 THEN
            exp_f := 2;
        ELSIF x =- 14333 THEN
            exp_f := 2;
        ELSIF x =- 14332 THEN
            exp_f := 2;
        ELSIF x =- 14331 THEN
            exp_f := 2;
        ELSIF x =- 14330 THEN
            exp_f := 2;
        ELSIF x =- 14329 THEN
            exp_f := 2;
        ELSIF x =- 14328 THEN
            exp_f := 2;
        ELSIF x =- 14327 THEN
            exp_f := 2;
        ELSIF x =- 14326 THEN
            exp_f := 2;
        ELSIF x =- 14325 THEN
            exp_f := 2;
        ELSIF x =- 14324 THEN
            exp_f := 2;
        ELSIF x =- 14323 THEN
            exp_f := 2;
        ELSIF x =- 14322 THEN
            exp_f := 2;
        ELSIF x =- 14321 THEN
            exp_f := 2;
        ELSIF x =- 14320 THEN
            exp_f := 2;
        ELSIF x =- 14319 THEN
            exp_f := 2;
        ELSIF x =- 14318 THEN
            exp_f := 2;
        ELSIF x =- 14317 THEN
            exp_f := 2;
        ELSIF x =- 14316 THEN
            exp_f := 2;
        ELSIF x =- 14315 THEN
            exp_f := 2;
        ELSIF x =- 14314 THEN
            exp_f := 2;
        ELSIF x =- 14313 THEN
            exp_f := 2;
        ELSIF x =- 14312 THEN
            exp_f := 2;
        ELSIF x =- 14311 THEN
            exp_f := 2;
        ELSIF x =- 14310 THEN
            exp_f := 2;
        ELSIF x =- 14309 THEN
            exp_f := 2;
        ELSIF x =- 14308 THEN
            exp_f := 2;
        ELSIF x =- 14307 THEN
            exp_f := 2;
        ELSIF x =- 14306 THEN
            exp_f := 2;
        ELSIF x =- 14305 THEN
            exp_f := 2;
        ELSIF x =- 14304 THEN
            exp_f := 2;
        ELSIF x =- 14303 THEN
            exp_f := 2;
        ELSIF x =- 14302 THEN
            exp_f := 2;
        ELSIF x =- 14301 THEN
            exp_f := 2;
        ELSIF x =- 14300 THEN
            exp_f := 2;
        ELSIF x =- 14299 THEN
            exp_f := 2;
        ELSIF x =- 14298 THEN
            exp_f := 2;
        ELSIF x =- 14297 THEN
            exp_f := 2;
        ELSIF x =- 14296 THEN
            exp_f := 2;
        ELSIF x =- 14295 THEN
            exp_f := 2;
        ELSIF x =- 14294 THEN
            exp_f := 2;
        ELSIF x =- 14293 THEN
            exp_f := 2;
        ELSIF x =- 14292 THEN
            exp_f := 2;
        ELSIF x =- 14291 THEN
            exp_f := 2;
        ELSIF x =- 14290 THEN
            exp_f := 2;
        ELSIF x =- 14289 THEN
            exp_f := 2;
        ELSIF x =- 14288 THEN
            exp_f := 2;
        ELSIF x =- 14287 THEN
            exp_f := 2;
        ELSIF x =- 14286 THEN
            exp_f := 2;
        ELSIF x =- 14285 THEN
            exp_f := 2;
        ELSIF x =- 14284 THEN
            exp_f := 2;
        ELSIF x =- 14283 THEN
            exp_f := 2;
        ELSIF x =- 14282 THEN
            exp_f := 2;
        ELSIF x =- 14281 THEN
            exp_f := 2;
        ELSIF x =- 14280 THEN
            exp_f := 2;
        ELSIF x =- 14279 THEN
            exp_f := 2;
        ELSIF x =- 14278 THEN
            exp_f := 2;
        ELSIF x =- 14277 THEN
            exp_f := 2;
        ELSIF x =- 14276 THEN
            exp_f := 2;
        ELSIF x =- 14275 THEN
            exp_f := 2;
        ELSIF x =- 14274 THEN
            exp_f := 2;
        ELSIF x =- 14273 THEN
            exp_f := 2;
        ELSIF x =- 14272 THEN
            exp_f := 2;
        ELSIF x =- 14271 THEN
            exp_f := 2;
        ELSIF x =- 14270 THEN
            exp_f := 2;
        ELSIF x =- 14269 THEN
            exp_f := 2;
        ELSIF x =- 14268 THEN
            exp_f := 2;
        ELSIF x =- 14267 THEN
            exp_f := 2;
        ELSIF x =- 14266 THEN
            exp_f := 2;
        ELSIF x =- 14265 THEN
            exp_f := 2;
        ELSIF x =- 14264 THEN
            exp_f := 2;
        ELSIF x =- 14263 THEN
            exp_f := 2;
        ELSIF x =- 14262 THEN
            exp_f := 2;
        ELSIF x =- 14261 THEN
            exp_f := 2;
        ELSIF x =- 14260 THEN
            exp_f := 2;
        ELSIF x =- 14259 THEN
            exp_f := 2;
        ELSIF x =- 14258 THEN
            exp_f := 2;
        ELSIF x =- 14257 THEN
            exp_f := 2;
        ELSIF x =- 14256 THEN
            exp_f := 2;
        ELSIF x =- 14255 THEN
            exp_f := 2;
        ELSIF x =- 14254 THEN
            exp_f := 2;
        ELSIF x =- 14253 THEN
            exp_f := 2;
        ELSIF x =- 14252 THEN
            exp_f := 2;
        ELSIF x =- 14251 THEN
            exp_f := 2;
        ELSIF x =- 14250 THEN
            exp_f := 2;
        ELSIF x =- 14249 THEN
            exp_f := 2;
        ELSIF x =- 14248 THEN
            exp_f := 2;
        ELSIF x =- 14247 THEN
            exp_f := 2;
        ELSIF x =- 14246 THEN
            exp_f := 2;
        ELSIF x =- 14245 THEN
            exp_f := 2;
        ELSIF x =- 14244 THEN
            exp_f := 2;
        ELSIF x =- 14243 THEN
            exp_f := 2;
        ELSIF x =- 14242 THEN
            exp_f := 2;
        ELSIF x =- 14241 THEN
            exp_f := 2;
        ELSIF x =- 14240 THEN
            exp_f := 2;
        ELSIF x =- 14239 THEN
            exp_f := 2;
        ELSIF x =- 14238 THEN
            exp_f := 2;
        ELSIF x =- 14237 THEN
            exp_f := 2;
        ELSIF x =- 14236 THEN
            exp_f := 2;
        ELSIF x =- 14235 THEN
            exp_f := 2;
        ELSIF x =- 14234 THEN
            exp_f := 2;
        ELSIF x =- 14233 THEN
            exp_f := 2;
        ELSIF x =- 14232 THEN
            exp_f := 2;
        ELSIF x =- 14231 THEN
            exp_f := 2;
        ELSIF x =- 14230 THEN
            exp_f := 2;
        ELSIF x =- 14229 THEN
            exp_f := 2;
        ELSIF x =- 14228 THEN
            exp_f := 2;
        ELSIF x =- 14227 THEN
            exp_f := 2;
        ELSIF x =- 14226 THEN
            exp_f := 2;
        ELSIF x =- 14225 THEN
            exp_f := 2;
        ELSIF x =- 14224 THEN
            exp_f := 2;
        ELSIF x =- 14223 THEN
            exp_f := 2;
        ELSIF x =- 14222 THEN
            exp_f := 2;
        ELSIF x =- 14221 THEN
            exp_f := 2;
        ELSIF x =- 14220 THEN
            exp_f := 2;
        ELSIF x =- 14219 THEN
            exp_f := 2;
        ELSIF x =- 14218 THEN
            exp_f := 2;
        ELSIF x =- 14217 THEN
            exp_f := 2;
        ELSIF x =- 14216 THEN
            exp_f := 2;
        ELSIF x =- 14215 THEN
            exp_f := 2;
        ELSIF x =- 14214 THEN
            exp_f := 2;
        ELSIF x =- 14213 THEN
            exp_f := 2;
        ELSIF x =- 14212 THEN
            exp_f := 2;
        ELSIF x =- 14211 THEN
            exp_f := 2;
        ELSIF x =- 14210 THEN
            exp_f := 2;
        ELSIF x =- 14209 THEN
            exp_f := 2;
        ELSIF x =- 14208 THEN
            exp_f := 2;
        ELSIF x =- 14207 THEN
            exp_f := 2;
        ELSIF x =- 14206 THEN
            exp_f := 2;
        ELSIF x =- 14205 THEN
            exp_f := 2;
        ELSIF x =- 14204 THEN
            exp_f := 2;
        ELSIF x =- 14203 THEN
            exp_f := 2;
        ELSIF x =- 14202 THEN
            exp_f := 2;
        ELSIF x =- 14201 THEN
            exp_f := 2;
        ELSIF x =- 14200 THEN
            exp_f := 2;
        ELSIF x =- 14199 THEN
            exp_f := 2;
        ELSIF x =- 14198 THEN
            exp_f := 2;
        ELSIF x =- 14197 THEN
            exp_f := 2;
        ELSIF x =- 14196 THEN
            exp_f := 2;
        ELSIF x =- 14195 THEN
            exp_f := 2;
        ELSIF x =- 14194 THEN
            exp_f := 2;
        ELSIF x =- 14193 THEN
            exp_f := 2;
        ELSIF x =- 14192 THEN
            exp_f := 2;
        ELSIF x =- 14191 THEN
            exp_f := 2;
        ELSIF x =- 14190 THEN
            exp_f := 2;
        ELSIF x =- 14189 THEN
            exp_f := 2;
        ELSIF x =- 14188 THEN
            exp_f := 2;
        ELSIF x =- 14187 THEN
            exp_f := 2;
        ELSIF x =- 14186 THEN
            exp_f := 2;
        ELSIF x =- 14185 THEN
            exp_f := 2;
        ELSIF x =- 14184 THEN
            exp_f := 2;
        ELSIF x =- 14183 THEN
            exp_f := 2;
        ELSIF x =- 14182 THEN
            exp_f := 2;
        ELSIF x =- 14181 THEN
            exp_f := 2;
        ELSIF x =- 14180 THEN
            exp_f := 2;
        ELSIF x =- 14179 THEN
            exp_f := 2;
        ELSIF x =- 14178 THEN
            exp_f := 2;
        ELSIF x =- 14177 THEN
            exp_f := 2;
        ELSIF x =- 14176 THEN
            exp_f := 2;
        ELSIF x =- 14175 THEN
            exp_f := 2;
        ELSIF x =- 14174 THEN
            exp_f := 2;
        ELSIF x =- 14173 THEN
            exp_f := 2;
        ELSIF x =- 14172 THEN
            exp_f := 2;
        ELSIF x =- 14171 THEN
            exp_f := 2;
        ELSIF x =- 14170 THEN
            exp_f := 2;
        ELSIF x =- 14169 THEN
            exp_f := 2;
        ELSIF x =- 14168 THEN
            exp_f := 2;
        ELSIF x =- 14167 THEN
            exp_f := 2;
        ELSIF x =- 14166 THEN
            exp_f := 2;
        ELSIF x =- 14165 THEN
            exp_f := 2;
        ELSIF x =- 14164 THEN
            exp_f := 2;
        ELSIF x =- 14163 THEN
            exp_f := 2;
        ELSIF x =- 14162 THEN
            exp_f := 2;
        ELSIF x =- 14161 THEN
            exp_f := 2;
        ELSIF x =- 14160 THEN
            exp_f := 2;
        ELSIF x =- 14159 THEN
            exp_f := 2;
        ELSIF x =- 14158 THEN
            exp_f := 2;
        ELSIF x =- 14157 THEN
            exp_f := 2;
        ELSIF x =- 14156 THEN
            exp_f := 2;
        ELSIF x =- 14155 THEN
            exp_f := 2;
        ELSIF x =- 14154 THEN
            exp_f := 2;
        ELSIF x =- 14153 THEN
            exp_f := 2;
        ELSIF x =- 14152 THEN
            exp_f := 2;
        ELSIF x =- 14151 THEN
            exp_f := 2;
        ELSIF x =- 14150 THEN
            exp_f := 2;
        ELSIF x =- 14149 THEN
            exp_f := 2;
        ELSIF x =- 14148 THEN
            exp_f := 2;
        ELSIF x =- 14147 THEN
            exp_f := 2;
        ELSIF x =- 14146 THEN
            exp_f := 2;
        ELSIF x =- 14145 THEN
            exp_f := 2;
        ELSIF x =- 14144 THEN
            exp_f := 2;
        ELSIF x =- 14143 THEN
            exp_f := 2;
        ELSIF x =- 14142 THEN
            exp_f := 2;
        ELSIF x =- 14141 THEN
            exp_f := 2;
        ELSIF x =- 14140 THEN
            exp_f := 2;
        ELSIF x =- 14139 THEN
            exp_f := 2;
        ELSIF x =- 14138 THEN
            exp_f := 2;
        ELSIF x =- 14137 THEN
            exp_f := 2;
        ELSIF x =- 14136 THEN
            exp_f := 2;
        ELSIF x =- 14135 THEN
            exp_f := 2;
        ELSIF x =- 14134 THEN
            exp_f := 2;
        ELSIF x =- 14133 THEN
            exp_f := 2;
        ELSIF x =- 14132 THEN
            exp_f := 2;
        ELSIF x =- 14131 THEN
            exp_f := 2;
        ELSIF x =- 14130 THEN
            exp_f := 2;
        ELSIF x =- 14129 THEN
            exp_f := 2;
        ELSIF x =- 14128 THEN
            exp_f := 2;
        ELSIF x =- 14127 THEN
            exp_f := 2;
        ELSIF x =- 14126 THEN
            exp_f := 2;
        ELSIF x =- 14125 THEN
            exp_f := 2;
        ELSIF x =- 14124 THEN
            exp_f := 2;
        ELSIF x =- 14123 THEN
            exp_f := 2;
        ELSIF x =- 14122 THEN
            exp_f := 2;
        ELSIF x =- 14121 THEN
            exp_f := 2;
        ELSIF x =- 14120 THEN
            exp_f := 2;
        ELSIF x =- 14119 THEN
            exp_f := 2;
        ELSIF x =- 14118 THEN
            exp_f := 2;
        ELSIF x =- 14117 THEN
            exp_f := 2;
        ELSIF x =- 14116 THEN
            exp_f := 2;
        ELSIF x =- 14115 THEN
            exp_f := 2;
        ELSIF x =- 14114 THEN
            exp_f := 2;
        ELSIF x =- 14113 THEN
            exp_f := 2;
        ELSIF x =- 14112 THEN
            exp_f := 2;
        ELSIF x =- 14111 THEN
            exp_f := 2;
        ELSIF x =- 14110 THEN
            exp_f := 2;
        ELSIF x =- 14109 THEN
            exp_f := 2;
        ELSIF x =- 14108 THEN
            exp_f := 2;
        ELSIF x =- 14107 THEN
            exp_f := 2;
        ELSIF x =- 14106 THEN
            exp_f := 2;
        ELSIF x =- 14105 THEN
            exp_f := 2;
        ELSIF x =- 14104 THEN
            exp_f := 2;
        ELSIF x =- 14103 THEN
            exp_f := 2;
        ELSIF x =- 14102 THEN
            exp_f := 2;
        ELSIF x =- 14101 THEN
            exp_f := 2;
        ELSIF x =- 14100 THEN
            exp_f := 2;
        ELSIF x =- 14099 THEN
            exp_f := 2;
        ELSIF x =- 14098 THEN
            exp_f := 2;
        ELSIF x =- 14097 THEN
            exp_f := 2;
        ELSIF x =- 14096 THEN
            exp_f := 2;
        ELSIF x =- 14095 THEN
            exp_f := 2;
        ELSIF x =- 14094 THEN
            exp_f := 2;
        ELSIF x =- 14093 THEN
            exp_f := 2;
        ELSIF x =- 14092 THEN
            exp_f := 2;
        ELSIF x =- 14091 THEN
            exp_f := 2;
        ELSIF x =- 14090 THEN
            exp_f := 2;
        ELSIF x =- 14089 THEN
            exp_f := 2;
        ELSIF x =- 14088 THEN
            exp_f := 2;
        ELSIF x =- 14087 THEN
            exp_f := 2;
        ELSIF x =- 14086 THEN
            exp_f := 2;
        ELSIF x =- 14085 THEN
            exp_f := 2;
        ELSIF x =- 14084 THEN
            exp_f := 2;
        ELSIF x =- 14083 THEN
            exp_f := 2;
        ELSIF x =- 14082 THEN
            exp_f := 2;
        ELSIF x =- 14081 THEN
            exp_f := 2;
        ELSIF x =- 14080 THEN
            exp_f := 2;
        ELSIF x =- 14079 THEN
            exp_f := 2;
        ELSIF x =- 14078 THEN
            exp_f := 2;
        ELSIF x =- 14077 THEN
            exp_f := 2;
        ELSIF x =- 14076 THEN
            exp_f := 2;
        ELSIF x =- 14075 THEN
            exp_f := 2;
        ELSIF x =- 14074 THEN
            exp_f := 2;
        ELSIF x =- 14073 THEN
            exp_f := 2;
        ELSIF x =- 14072 THEN
            exp_f := 2;
        ELSIF x =- 14071 THEN
            exp_f := 2;
        ELSIF x =- 14070 THEN
            exp_f := 2;
        ELSIF x =- 14069 THEN
            exp_f := 2;
        ELSIF x =- 14068 THEN
            exp_f := 2;
        ELSIF x =- 14067 THEN
            exp_f := 2;
        ELSIF x =- 14066 THEN
            exp_f := 2;
        ELSIF x =- 14065 THEN
            exp_f := 2;
        ELSIF x =- 14064 THEN
            exp_f := 2;
        ELSIF x =- 14063 THEN
            exp_f := 2;
        ELSIF x =- 14062 THEN
            exp_f := 2;
        ELSIF x =- 14061 THEN
            exp_f := 2;
        ELSIF x =- 14060 THEN
            exp_f := 2;
        ELSIF x =- 14059 THEN
            exp_f := 2;
        ELSIF x =- 14058 THEN
            exp_f := 2;
        ELSIF x =- 14057 THEN
            exp_f := 2;
        ELSIF x =- 14056 THEN
            exp_f := 2;
        ELSIF x =- 14055 THEN
            exp_f := 2;
        ELSIF x =- 14054 THEN
            exp_f := 2;
        ELSIF x =- 14053 THEN
            exp_f := 2;
        ELSIF x =- 14052 THEN
            exp_f := 2;
        ELSIF x =- 14051 THEN
            exp_f := 2;
        ELSIF x =- 14050 THEN
            exp_f := 2;
        ELSIF x =- 14049 THEN
            exp_f := 2;
        ELSIF x =- 14048 THEN
            exp_f := 2;
        ELSIF x =- 14047 THEN
            exp_f := 2;
        ELSIF x =- 14046 THEN
            exp_f := 2;
        ELSIF x =- 14045 THEN
            exp_f := 2;
        ELSIF x =- 14044 THEN
            exp_f := 2;
        ELSIF x =- 14043 THEN
            exp_f := 2;
        ELSIF x =- 14042 THEN
            exp_f := 2;
        ELSIF x =- 14041 THEN
            exp_f := 2;
        ELSIF x =- 14040 THEN
            exp_f := 2;
        ELSIF x =- 14039 THEN
            exp_f := 2;
        ELSIF x =- 14038 THEN
            exp_f := 2;
        ELSIF x =- 14037 THEN
            exp_f := 2;
        ELSIF x =- 14036 THEN
            exp_f := 2;
        ELSIF x =- 14035 THEN
            exp_f := 2;
        ELSIF x =- 14034 THEN
            exp_f := 2;
        ELSIF x =- 14033 THEN
            exp_f := 2;
        ELSIF x =- 14032 THEN
            exp_f := 2;
        ELSIF x =- 14031 THEN
            exp_f := 2;
        ELSIF x =- 14030 THEN
            exp_f := 2;
        ELSIF x =- 14029 THEN
            exp_f := 2;
        ELSIF x =- 14028 THEN
            exp_f := 2;
        ELSIF x =- 14027 THEN
            exp_f := 2;
        ELSIF x =- 14026 THEN
            exp_f := 2;
        ELSIF x =- 14025 THEN
            exp_f := 2;
        ELSIF x =- 14024 THEN
            exp_f := 2;
        ELSIF x =- 14023 THEN
            exp_f := 2;
        ELSIF x =- 14022 THEN
            exp_f := 2;
        ELSIF x =- 14021 THEN
            exp_f := 2;
        ELSIF x =- 14020 THEN
            exp_f := 2;
        ELSIF x =- 14019 THEN
            exp_f := 2;
        ELSIF x =- 14018 THEN
            exp_f := 2;
        ELSIF x =- 14017 THEN
            exp_f := 2;
        ELSIF x =- 14016 THEN
            exp_f := 2;
        ELSIF x =- 14015 THEN
            exp_f := 2;
        ELSIF x =- 14014 THEN
            exp_f := 2;
        ELSIF x =- 14013 THEN
            exp_f := 2;
        ELSIF x =- 14012 THEN
            exp_f := 2;
        ELSIF x =- 14011 THEN
            exp_f := 2;
        ELSIF x =- 14010 THEN
            exp_f := 2;
        ELSIF x =- 14009 THEN
            exp_f := 2;
        ELSIF x =- 14008 THEN
            exp_f := 2;
        ELSIF x =- 14007 THEN
            exp_f := 2;
        ELSIF x =- 14006 THEN
            exp_f := 2;
        ELSIF x =- 14005 THEN
            exp_f := 2;
        ELSIF x =- 14004 THEN
            exp_f := 2;
        ELSIF x =- 14003 THEN
            exp_f := 2;
        ELSIF x =- 14002 THEN
            exp_f := 2;
        ELSIF x =- 14001 THEN
            exp_f := 2;
        ELSIF x =- 14000 THEN
            exp_f := 2;
        ELSIF x =- 13999 THEN
            exp_f := 2;
        ELSIF x =- 13998 THEN
            exp_f := 2;
        ELSIF x =- 13997 THEN
            exp_f := 2;
        ELSIF x =- 13996 THEN
            exp_f := 2;
        ELSIF x =- 13995 THEN
            exp_f := 2;
        ELSIF x =- 13994 THEN
            exp_f := 2;
        ELSIF x =- 13993 THEN
            exp_f := 2;
        ELSIF x =- 13992 THEN
            exp_f := 2;
        ELSIF x =- 13991 THEN
            exp_f := 2;
        ELSIF x =- 13990 THEN
            exp_f := 2;
        ELSIF x =- 13989 THEN
            exp_f := 2;
        ELSIF x =- 13988 THEN
            exp_f := 2;
        ELSIF x =- 13987 THEN
            exp_f := 2;
        ELSIF x =- 13986 THEN
            exp_f := 2;
        ELSIF x =- 13985 THEN
            exp_f := 2;
        ELSIF x =- 13984 THEN
            exp_f := 2;
        ELSIF x =- 13983 THEN
            exp_f := 2;
        ELSIF x =- 13982 THEN
            exp_f := 2;
        ELSIF x =- 13981 THEN
            exp_f := 2;
        ELSIF x =- 13980 THEN
            exp_f := 2;
        ELSIF x =- 13979 THEN
            exp_f := 2;
        ELSIF x =- 13978 THEN
            exp_f := 2;
        ELSIF x =- 13977 THEN
            exp_f := 2;
        ELSIF x =- 13976 THEN
            exp_f := 2;
        ELSIF x =- 13975 THEN
            exp_f := 2;
        ELSIF x =- 13974 THEN
            exp_f := 2;
        ELSIF x =- 13973 THEN
            exp_f := 2;
        ELSIF x =- 13972 THEN
            exp_f := 2;
        ELSIF x =- 13971 THEN
            exp_f := 2;
        ELSIF x =- 13970 THEN
            exp_f := 2;
        ELSIF x =- 13969 THEN
            exp_f := 2;
        ELSIF x =- 13968 THEN
            exp_f := 2;
        ELSIF x =- 13967 THEN
            exp_f := 2;
        ELSIF x =- 13966 THEN
            exp_f := 2;
        ELSIF x =- 13965 THEN
            exp_f := 2;
        ELSIF x =- 13964 THEN
            exp_f := 2;
        ELSIF x =- 13963 THEN
            exp_f := 2;
        ELSIF x =- 13962 THEN
            exp_f := 2;
        ELSIF x =- 13961 THEN
            exp_f := 2;
        ELSIF x =- 13960 THEN
            exp_f := 2;
        ELSIF x =- 13959 THEN
            exp_f := 2;
        ELSIF x =- 13958 THEN
            exp_f := 2;
        ELSIF x =- 13957 THEN
            exp_f := 2;
        ELSIF x =- 13956 THEN
            exp_f := 2;
        ELSIF x =- 13955 THEN
            exp_f := 2;
        ELSIF x =- 13954 THEN
            exp_f := 2;
        ELSIF x =- 13953 THEN
            exp_f := 2;
        ELSIF x =- 13952 THEN
            exp_f := 2;
        ELSIF x =- 13951 THEN
            exp_f := 2;
        ELSIF x =- 13950 THEN
            exp_f := 2;
        ELSIF x =- 13949 THEN
            exp_f := 2;
        ELSIF x =- 13948 THEN
            exp_f := 2;
        ELSIF x =- 13947 THEN
            exp_f := 2;
        ELSIF x =- 13946 THEN
            exp_f := 2;
        ELSIF x =- 13945 THEN
            exp_f := 2;
        ELSIF x =- 13944 THEN
            exp_f := 2;
        ELSIF x =- 13943 THEN
            exp_f := 2;
        ELSIF x =- 13942 THEN
            exp_f := 2;
        ELSIF x =- 13941 THEN
            exp_f := 2;
        ELSIF x =- 13940 THEN
            exp_f := 2;
        ELSIF x =- 13939 THEN
            exp_f := 2;
        ELSIF x =- 13938 THEN
            exp_f := 2;
        ELSIF x =- 13937 THEN
            exp_f := 2;
        ELSIF x =- 13936 THEN
            exp_f := 2;
        ELSIF x =- 13935 THEN
            exp_f := 2;
        ELSIF x =- 13934 THEN
            exp_f := 2;
        ELSIF x =- 13933 THEN
            exp_f := 2;
        ELSIF x =- 13932 THEN
            exp_f := 2;
        ELSIF x =- 13931 THEN
            exp_f := 2;
        ELSIF x =- 13930 THEN
            exp_f := 2;
        ELSIF x =- 13929 THEN
            exp_f := 2;
        ELSIF x =- 13928 THEN
            exp_f := 2;
        ELSIF x =- 13927 THEN
            exp_f := 2;
        ELSIF x =- 13926 THEN
            exp_f := 2;
        ELSIF x =- 13925 THEN
            exp_f := 2;
        ELSIF x =- 13924 THEN
            exp_f := 2;
        ELSIF x =- 13923 THEN
            exp_f := 2;
        ELSIF x =- 13922 THEN
            exp_f := 2;
        ELSIF x =- 13921 THEN
            exp_f := 2;
        ELSIF x =- 13920 THEN
            exp_f := 2;
        ELSIF x =- 13919 THEN
            exp_f := 2;
        ELSIF x =- 13918 THEN
            exp_f := 2;
        ELSIF x =- 13917 THEN
            exp_f := 2;
        ELSIF x =- 13916 THEN
            exp_f := 2;
        ELSIF x =- 13915 THEN
            exp_f := 2;
        ELSIF x =- 13914 THEN
            exp_f := 2;
        ELSIF x =- 13913 THEN
            exp_f := 2;
        ELSIF x =- 13912 THEN
            exp_f := 2;
        ELSIF x =- 13911 THEN
            exp_f := 2;
        ELSIF x =- 13910 THEN
            exp_f := 2;
        ELSIF x =- 13909 THEN
            exp_f := 2;
        ELSIF x =- 13908 THEN
            exp_f := 2;
        ELSIF x =- 13907 THEN
            exp_f := 2;
        ELSIF x =- 13906 THEN
            exp_f := 2;
        ELSIF x =- 13905 THEN
            exp_f := 2;
        ELSIF x =- 13904 THEN
            exp_f := 2;
        ELSIF x =- 13903 THEN
            exp_f := 2;
        ELSIF x =- 13902 THEN
            exp_f := 2;
        ELSIF x =- 13901 THEN
            exp_f := 2;
        ELSIF x =- 13900 THEN
            exp_f := 2;
        ELSIF x =- 13899 THEN
            exp_f := 2;
        ELSIF x =- 13898 THEN
            exp_f := 2;
        ELSIF x =- 13897 THEN
            exp_f := 2;
        ELSIF x =- 13896 THEN
            exp_f := 2;
        ELSIF x =- 13895 THEN
            exp_f := 2;
        ELSIF x =- 13894 THEN
            exp_f := 2;
        ELSIF x =- 13893 THEN
            exp_f := 2;
        ELSIF x =- 13892 THEN
            exp_f := 2;
        ELSIF x =- 13891 THEN
            exp_f := 2;
        ELSIF x =- 13890 THEN
            exp_f := 2;
        ELSIF x =- 13889 THEN
            exp_f := 2;
        ELSIF x =- 13888 THEN
            exp_f := 2;
        ELSIF x =- 13887 THEN
            exp_f := 2;
        ELSIF x =- 13886 THEN
            exp_f := 2;
        ELSIF x =- 13885 THEN
            exp_f := 2;
        ELSIF x =- 13884 THEN
            exp_f := 2;
        ELSIF x =- 13883 THEN
            exp_f := 2;
        ELSIF x =- 13882 THEN
            exp_f := 2;
        ELSIF x =- 13881 THEN
            exp_f := 2;
        ELSIF x =- 13880 THEN
            exp_f := 2;
        ELSIF x =- 13879 THEN
            exp_f := 2;
        ELSIF x =- 13878 THEN
            exp_f := 2;
        ELSIF x =- 13877 THEN
            exp_f := 2;
        ELSIF x =- 13876 THEN
            exp_f := 2;
        ELSIF x =- 13875 THEN
            exp_f := 2;
        ELSIF x =- 13874 THEN
            exp_f := 2;
        ELSIF x =- 13873 THEN
            exp_f := 2;
        ELSIF x =- 13872 THEN
            exp_f := 2;
        ELSIF x =- 13871 THEN
            exp_f := 2;
        ELSIF x =- 13870 THEN
            exp_f := 2;
        ELSIF x =- 13869 THEN
            exp_f := 2;
        ELSIF x =- 13868 THEN
            exp_f := 2;
        ELSIF x =- 13867 THEN
            exp_f := 2;
        ELSIF x =- 13866 THEN
            exp_f := 2;
        ELSIF x =- 13865 THEN
            exp_f := 2;
        ELSIF x =- 13864 THEN
            exp_f := 2;
        ELSIF x =- 13863 THEN
            exp_f := 2;
        ELSIF x =- 13862 THEN
            exp_f := 2;
        ELSIF x =- 13861 THEN
            exp_f := 2;
        ELSIF x =- 13860 THEN
            exp_f := 2;
        ELSIF x =- 13859 THEN
            exp_f := 2;
        ELSIF x =- 13858 THEN
            exp_f := 2;
        ELSIF x =- 13857 THEN
            exp_f := 2;
        ELSIF x =- 13856 THEN
            exp_f := 2;
        ELSIF x =- 13855 THEN
            exp_f := 2;
        ELSIF x =- 13854 THEN
            exp_f := 2;
        ELSIF x =- 13853 THEN
            exp_f := 2;
        ELSIF x =- 13852 THEN
            exp_f := 2;
        ELSIF x =- 13851 THEN
            exp_f := 2;
        ELSIF x =- 13850 THEN
            exp_f := 2;
        ELSIF x =- 13849 THEN
            exp_f := 2;
        ELSIF x =- 13848 THEN
            exp_f := 2;
        ELSIF x =- 13847 THEN
            exp_f := 2;
        ELSIF x =- 13846 THEN
            exp_f := 2;
        ELSIF x =- 13845 THEN
            exp_f := 2;
        ELSIF x =- 13844 THEN
            exp_f := 2;
        ELSIF x =- 13843 THEN
            exp_f := 2;
        ELSIF x =- 13842 THEN
            exp_f := 2;
        ELSIF x =- 13841 THEN
            exp_f := 2;
        ELSIF x =- 13840 THEN
            exp_f := 2;
        ELSIF x =- 13839 THEN
            exp_f := 2;
        ELSIF x =- 13838 THEN
            exp_f := 2;
        ELSIF x =- 13837 THEN
            exp_f := 2;
        ELSIF x =- 13836 THEN
            exp_f := 2;
        ELSIF x =- 13835 THEN
            exp_f := 2;
        ELSIF x =- 13834 THEN
            exp_f := 2;
        ELSIF x =- 13833 THEN
            exp_f := 2;
        ELSIF x =- 13832 THEN
            exp_f := 2;
        ELSIF x =- 13831 THEN
            exp_f := 2;
        ELSIF x =- 13830 THEN
            exp_f := 2;
        ELSIF x =- 13829 THEN
            exp_f := 2;
        ELSIF x =- 13828 THEN
            exp_f := 2;
        ELSIF x =- 13827 THEN
            exp_f := 2;
        ELSIF x =- 13826 THEN
            exp_f := 2;
        ELSIF x =- 13825 THEN
            exp_f := 2;
        ELSIF x =- 13824 THEN
            exp_f := 2;
        ELSIF x =- 13823 THEN
            exp_f := 3;
        ELSIF x =- 13822 THEN
            exp_f := 3;
        ELSIF x =- 13821 THEN
            exp_f := 3;
        ELSIF x =- 13820 THEN
            exp_f := 3;
        ELSIF x =- 13819 THEN
            exp_f := 3;
        ELSIF x =- 13818 THEN
            exp_f := 3;
        ELSIF x =- 13817 THEN
            exp_f := 3;
        ELSIF x =- 13816 THEN
            exp_f := 3;
        ELSIF x =- 13815 THEN
            exp_f := 3;
        ELSIF x =- 13814 THEN
            exp_f := 3;
        ELSIF x =- 13813 THEN
            exp_f := 3;
        ELSIF x =- 13812 THEN
            exp_f := 3;
        ELSIF x =- 13811 THEN
            exp_f := 3;
        ELSIF x =- 13810 THEN
            exp_f := 3;
        ELSIF x =- 13809 THEN
            exp_f := 3;
        ELSIF x =- 13808 THEN
            exp_f := 3;
        ELSIF x =- 13807 THEN
            exp_f := 3;
        ELSIF x =- 13806 THEN
            exp_f := 3;
        ELSIF x =- 13805 THEN
            exp_f := 3;
        ELSIF x =- 13804 THEN
            exp_f := 3;
        ELSIF x =- 13803 THEN
            exp_f := 3;
        ELSIF x =- 13802 THEN
            exp_f := 3;
        ELSIF x =- 13801 THEN
            exp_f := 3;
        ELSIF x =- 13800 THEN
            exp_f := 3;
        ELSIF x =- 13799 THEN
            exp_f := 3;
        ELSIF x =- 13798 THEN
            exp_f := 3;
        ELSIF x =- 13797 THEN
            exp_f := 3;
        ELSIF x =- 13796 THEN
            exp_f := 3;
        ELSIF x =- 13795 THEN
            exp_f := 3;
        ELSIF x =- 13794 THEN
            exp_f := 3;
        ELSIF x =- 13793 THEN
            exp_f := 3;
        ELSIF x =- 13792 THEN
            exp_f := 3;
        ELSIF x =- 13791 THEN
            exp_f := 3;
        ELSIF x =- 13790 THEN
            exp_f := 3;
        ELSIF x =- 13789 THEN
            exp_f := 3;
        ELSIF x =- 13788 THEN
            exp_f := 3;
        ELSIF x =- 13787 THEN
            exp_f := 3;
        ELSIF x =- 13786 THEN
            exp_f := 3;
        ELSIF x =- 13785 THEN
            exp_f := 3;
        ELSIF x =- 13784 THEN
            exp_f := 3;
        ELSIF x =- 13783 THEN
            exp_f := 3;
        ELSIF x =- 13782 THEN
            exp_f := 3;
        ELSIF x =- 13781 THEN
            exp_f := 3;
        ELSIF x =- 13780 THEN
            exp_f := 3;
        ELSIF x =- 13779 THEN
            exp_f := 3;
        ELSIF x =- 13778 THEN
            exp_f := 3;
        ELSIF x =- 13777 THEN
            exp_f := 3;
        ELSIF x =- 13776 THEN
            exp_f := 3;
        ELSIF x =- 13775 THEN
            exp_f := 3;
        ELSIF x =- 13774 THEN
            exp_f := 3;
        ELSIF x =- 13773 THEN
            exp_f := 3;
        ELSIF x =- 13772 THEN
            exp_f := 3;
        ELSIF x =- 13771 THEN
            exp_f := 3;
        ELSIF x =- 13770 THEN
            exp_f := 3;
        ELSIF x =- 13769 THEN
            exp_f := 3;
        ELSIF x =- 13768 THEN
            exp_f := 3;
        ELSIF x =- 13767 THEN
            exp_f := 3;
        ELSIF x =- 13766 THEN
            exp_f := 3;
        ELSIF x =- 13765 THEN
            exp_f := 3;
        ELSIF x =- 13764 THEN
            exp_f := 3;
        ELSIF x =- 13763 THEN
            exp_f := 3;
        ELSIF x =- 13762 THEN
            exp_f := 3;
        ELSIF x =- 13761 THEN
            exp_f := 3;
        ELSIF x =- 13760 THEN
            exp_f := 3;
        ELSIF x =- 13759 THEN
            exp_f := 3;
        ELSIF x =- 13758 THEN
            exp_f := 3;
        ELSIF x =- 13757 THEN
            exp_f := 3;
        ELSIF x =- 13756 THEN
            exp_f := 3;
        ELSIF x =- 13755 THEN
            exp_f := 3;
        ELSIF x =- 13754 THEN
            exp_f := 3;
        ELSIF x =- 13753 THEN
            exp_f := 3;
        ELSIF x =- 13752 THEN
            exp_f := 3;
        ELSIF x =- 13751 THEN
            exp_f := 3;
        ELSIF x =- 13750 THEN
            exp_f := 3;
        ELSIF x =- 13749 THEN
            exp_f := 3;
        ELSIF x =- 13748 THEN
            exp_f := 3;
        ELSIF x =- 13747 THEN
            exp_f := 3;
        ELSIF x =- 13746 THEN
            exp_f := 3;
        ELSIF x =- 13745 THEN
            exp_f := 3;
        ELSIF x =- 13744 THEN
            exp_f := 3;
        ELSIF x =- 13743 THEN
            exp_f := 3;
        ELSIF x =- 13742 THEN
            exp_f := 3;
        ELSIF x =- 13741 THEN
            exp_f := 3;
        ELSIF x =- 13740 THEN
            exp_f := 3;
        ELSIF x =- 13739 THEN
            exp_f := 3;
        ELSIF x =- 13738 THEN
            exp_f := 3;
        ELSIF x =- 13737 THEN
            exp_f := 3;
        ELSIF x =- 13736 THEN
            exp_f := 3;
        ELSIF x =- 13735 THEN
            exp_f := 3;
        ELSIF x =- 13734 THEN
            exp_f := 3;
        ELSIF x =- 13733 THEN
            exp_f := 3;
        ELSIF x =- 13732 THEN
            exp_f := 3;
        ELSIF x =- 13731 THEN
            exp_f := 3;
        ELSIF x =- 13730 THEN
            exp_f := 3;
        ELSIF x =- 13729 THEN
            exp_f := 3;
        ELSIF x =- 13728 THEN
            exp_f := 3;
        ELSIF x =- 13727 THEN
            exp_f := 3;
        ELSIF x =- 13726 THEN
            exp_f := 3;
        ELSIF x =- 13725 THEN
            exp_f := 3;
        ELSIF x =- 13724 THEN
            exp_f := 3;
        ELSIF x =- 13723 THEN
            exp_f := 3;
        ELSIF x =- 13722 THEN
            exp_f := 3;
        ELSIF x =- 13721 THEN
            exp_f := 3;
        ELSIF x =- 13720 THEN
            exp_f := 3;
        ELSIF x =- 13719 THEN
            exp_f := 3;
        ELSIF x =- 13718 THEN
            exp_f := 3;
        ELSIF x =- 13717 THEN
            exp_f := 3;
        ELSIF x =- 13716 THEN
            exp_f := 3;
        ELSIF x =- 13715 THEN
            exp_f := 3;
        ELSIF x =- 13714 THEN
            exp_f := 3;
        ELSIF x =- 13713 THEN
            exp_f := 3;
        ELSIF x =- 13712 THEN
            exp_f := 3;
        ELSIF x =- 13711 THEN
            exp_f := 3;
        ELSIF x =- 13710 THEN
            exp_f := 3;
        ELSIF x =- 13709 THEN
            exp_f := 3;
        ELSIF x =- 13708 THEN
            exp_f := 3;
        ELSIF x =- 13707 THEN
            exp_f := 3;
        ELSIF x =- 13706 THEN
            exp_f := 3;
        ELSIF x =- 13705 THEN
            exp_f := 3;
        ELSIF x =- 13704 THEN
            exp_f := 3;
        ELSIF x =- 13703 THEN
            exp_f := 3;
        ELSIF x =- 13702 THEN
            exp_f := 3;
        ELSIF x =- 13701 THEN
            exp_f := 3;
        ELSIF x =- 13700 THEN
            exp_f := 3;
        ELSIF x =- 13699 THEN
            exp_f := 3;
        ELSIF x =- 13698 THEN
            exp_f := 3;
        ELSIF x =- 13697 THEN
            exp_f := 3;
        ELSIF x =- 13696 THEN
            exp_f := 3;
        ELSIF x =- 13695 THEN
            exp_f := 3;
        ELSIF x =- 13694 THEN
            exp_f := 3;
        ELSIF x =- 13693 THEN
            exp_f := 3;
        ELSIF x =- 13692 THEN
            exp_f := 3;
        ELSIF x =- 13691 THEN
            exp_f := 3;
        ELSIF x =- 13690 THEN
            exp_f := 3;
        ELSIF x =- 13689 THEN
            exp_f := 3;
        ELSIF x =- 13688 THEN
            exp_f := 3;
        ELSIF x =- 13687 THEN
            exp_f := 3;
        ELSIF x =- 13686 THEN
            exp_f := 3;
        ELSIF x =- 13685 THEN
            exp_f := 3;
        ELSIF x =- 13684 THEN
            exp_f := 3;
        ELSIF x =- 13683 THEN
            exp_f := 3;
        ELSIF x =- 13682 THEN
            exp_f := 3;
        ELSIF x =- 13681 THEN
            exp_f := 3;
        ELSIF x =- 13680 THEN
            exp_f := 3;
        ELSIF x =- 13679 THEN
            exp_f := 3;
        ELSIF x =- 13678 THEN
            exp_f := 3;
        ELSIF x =- 13677 THEN
            exp_f := 3;
        ELSIF x =- 13676 THEN
            exp_f := 3;
        ELSIF x =- 13675 THEN
            exp_f := 3;
        ELSIF x =- 13674 THEN
            exp_f := 3;
        ELSIF x =- 13673 THEN
            exp_f := 3;
        ELSIF x =- 13672 THEN
            exp_f := 3;
        ELSIF x =- 13671 THEN
            exp_f := 3;
        ELSIF x =- 13670 THEN
            exp_f := 3;
        ELSIF x =- 13669 THEN
            exp_f := 3;
        ELSIF x =- 13668 THEN
            exp_f := 3;
        ELSIF x =- 13667 THEN
            exp_f := 3;
        ELSIF x =- 13666 THEN
            exp_f := 3;
        ELSIF x =- 13665 THEN
            exp_f := 3;
        ELSIF x =- 13664 THEN
            exp_f := 3;
        ELSIF x =- 13663 THEN
            exp_f := 3;
        ELSIF x =- 13662 THEN
            exp_f := 3;
        ELSIF x =- 13661 THEN
            exp_f := 3;
        ELSIF x =- 13660 THEN
            exp_f := 3;
        ELSIF x =- 13659 THEN
            exp_f := 3;
        ELSIF x =- 13658 THEN
            exp_f := 3;
        ELSIF x =- 13657 THEN
            exp_f := 3;
        ELSIF x =- 13656 THEN
            exp_f := 3;
        ELSIF x =- 13655 THEN
            exp_f := 3;
        ELSIF x =- 13654 THEN
            exp_f := 3;
        ELSIF x =- 13653 THEN
            exp_f := 3;
        ELSIF x =- 13652 THEN
            exp_f := 3;
        ELSIF x =- 13651 THEN
            exp_f := 3;
        ELSIF x =- 13650 THEN
            exp_f := 3;
        ELSIF x =- 13649 THEN
            exp_f := 3;
        ELSIF x =- 13648 THEN
            exp_f := 3;
        ELSIF x =- 13647 THEN
            exp_f := 3;
        ELSIF x =- 13646 THEN
            exp_f := 3;
        ELSIF x =- 13645 THEN
            exp_f := 3;
        ELSIF x =- 13644 THEN
            exp_f := 3;
        ELSIF x =- 13643 THEN
            exp_f := 3;
        ELSIF x =- 13642 THEN
            exp_f := 3;
        ELSIF x =- 13641 THEN
            exp_f := 3;
        ELSIF x =- 13640 THEN
            exp_f := 3;
        ELSIF x =- 13639 THEN
            exp_f := 3;
        ELSIF x =- 13638 THEN
            exp_f := 3;
        ELSIF x =- 13637 THEN
            exp_f := 3;
        ELSIF x =- 13636 THEN
            exp_f := 3;
        ELSIF x =- 13635 THEN
            exp_f := 3;
        ELSIF x =- 13634 THEN
            exp_f := 3;
        ELSIF x =- 13633 THEN
            exp_f := 3;
        ELSIF x =- 13632 THEN
            exp_f := 3;
        ELSIF x =- 13631 THEN
            exp_f := 3;
        ELSIF x =- 13630 THEN
            exp_f := 3;
        ELSIF x =- 13629 THEN
            exp_f := 3;
        ELSIF x =- 13628 THEN
            exp_f := 3;
        ELSIF x =- 13627 THEN
            exp_f := 3;
        ELSIF x =- 13626 THEN
            exp_f := 3;
        ELSIF x =- 13625 THEN
            exp_f := 3;
        ELSIF x =- 13624 THEN
            exp_f := 3;
        ELSIF x =- 13623 THEN
            exp_f := 3;
        ELSIF x =- 13622 THEN
            exp_f := 3;
        ELSIF x =- 13621 THEN
            exp_f := 3;
        ELSIF x =- 13620 THEN
            exp_f := 3;
        ELSIF x =- 13619 THEN
            exp_f := 3;
        ELSIF x =- 13618 THEN
            exp_f := 3;
        ELSIF x =- 13617 THEN
            exp_f := 3;
        ELSIF x =- 13616 THEN
            exp_f := 3;
        ELSIF x =- 13615 THEN
            exp_f := 3;
        ELSIF x =- 13614 THEN
            exp_f := 3;
        ELSIF x =- 13613 THEN
            exp_f := 3;
        ELSIF x =- 13612 THEN
            exp_f := 3;
        ELSIF x =- 13611 THEN
            exp_f := 3;
        ELSIF x =- 13610 THEN
            exp_f := 3;
        ELSIF x =- 13609 THEN
            exp_f := 3;
        ELSIF x =- 13608 THEN
            exp_f := 3;
        ELSIF x =- 13607 THEN
            exp_f := 3;
        ELSIF x =- 13606 THEN
            exp_f := 3;
        ELSIF x =- 13605 THEN
            exp_f := 3;
        ELSIF x =- 13604 THEN
            exp_f := 3;
        ELSIF x =- 13603 THEN
            exp_f := 3;
        ELSIF x =- 13602 THEN
            exp_f := 3;
        ELSIF x =- 13601 THEN
            exp_f := 3;
        ELSIF x =- 13600 THEN
            exp_f := 3;
        ELSIF x =- 13599 THEN
            exp_f := 3;
        ELSIF x =- 13598 THEN
            exp_f := 3;
        ELSIF x =- 13597 THEN
            exp_f := 3;
        ELSIF x =- 13596 THEN
            exp_f := 3;
        ELSIF x =- 13595 THEN
            exp_f := 3;
        ELSIF x =- 13594 THEN
            exp_f := 3;
        ELSIF x =- 13593 THEN
            exp_f := 3;
        ELSIF x =- 13592 THEN
            exp_f := 3;
        ELSIF x =- 13591 THEN
            exp_f := 3;
        ELSIF x =- 13590 THEN
            exp_f := 3;
        ELSIF x =- 13589 THEN
            exp_f := 3;
        ELSIF x =- 13588 THEN
            exp_f := 3;
        ELSIF x =- 13587 THEN
            exp_f := 3;
        ELSIF x =- 13586 THEN
            exp_f := 3;
        ELSIF x =- 13585 THEN
            exp_f := 3;
        ELSIF x =- 13584 THEN
            exp_f := 3;
        ELSIF x =- 13583 THEN
            exp_f := 3;
        ELSIF x =- 13582 THEN
            exp_f := 3;
        ELSIF x =- 13581 THEN
            exp_f := 3;
        ELSIF x =- 13580 THEN
            exp_f := 3;
        ELSIF x =- 13579 THEN
            exp_f := 3;
        ELSIF x =- 13578 THEN
            exp_f := 3;
        ELSIF x =- 13577 THEN
            exp_f := 3;
        ELSIF x =- 13576 THEN
            exp_f := 3;
        ELSIF x =- 13575 THEN
            exp_f := 3;
        ELSIF x =- 13574 THEN
            exp_f := 3;
        ELSIF x =- 13573 THEN
            exp_f := 3;
        ELSIF x =- 13572 THEN
            exp_f := 3;
        ELSIF x =- 13571 THEN
            exp_f := 3;
        ELSIF x =- 13570 THEN
            exp_f := 3;
        ELSIF x =- 13569 THEN
            exp_f := 3;
        ELSIF x =- 13568 THEN
            exp_f := 3;
        ELSIF x =- 13567 THEN
            exp_f := 3;
        ELSIF x =- 13566 THEN
            exp_f := 3;
        ELSIF x =- 13565 THEN
            exp_f := 3;
        ELSIF x =- 13564 THEN
            exp_f := 3;
        ELSIF x =- 13563 THEN
            exp_f := 3;
        ELSIF x =- 13562 THEN
            exp_f := 3;
        ELSIF x =- 13561 THEN
            exp_f := 3;
        ELSIF x =- 13560 THEN
            exp_f := 3;
        ELSIF x =- 13559 THEN
            exp_f := 3;
        ELSIF x =- 13558 THEN
            exp_f := 3;
        ELSIF x =- 13557 THEN
            exp_f := 3;
        ELSIF x =- 13556 THEN
            exp_f := 3;
        ELSIF x =- 13555 THEN
            exp_f := 3;
        ELSIF x =- 13554 THEN
            exp_f := 3;
        ELSIF x =- 13553 THEN
            exp_f := 3;
        ELSIF x =- 13552 THEN
            exp_f := 3;
        ELSIF x =- 13551 THEN
            exp_f := 3;
        ELSIF x =- 13550 THEN
            exp_f := 3;
        ELSIF x =- 13549 THEN
            exp_f := 3;
        ELSIF x =- 13548 THEN
            exp_f := 3;
        ELSIF x =- 13547 THEN
            exp_f := 3;
        ELSIF x =- 13546 THEN
            exp_f := 3;
        ELSIF x =- 13545 THEN
            exp_f := 3;
        ELSIF x =- 13544 THEN
            exp_f := 3;
        ELSIF x =- 13543 THEN
            exp_f := 3;
        ELSIF x =- 13542 THEN
            exp_f := 3;
        ELSIF x =- 13541 THEN
            exp_f := 3;
        ELSIF x =- 13540 THEN
            exp_f := 3;
        ELSIF x =- 13539 THEN
            exp_f := 3;
        ELSIF x =- 13538 THEN
            exp_f := 3;
        ELSIF x =- 13537 THEN
            exp_f := 3;
        ELSIF x =- 13536 THEN
            exp_f := 3;
        ELSIF x =- 13535 THEN
            exp_f := 3;
        ELSIF x =- 13534 THEN
            exp_f := 3;
        ELSIF x =- 13533 THEN
            exp_f := 3;
        ELSIF x =- 13532 THEN
            exp_f := 3;
        ELSIF x =- 13531 THEN
            exp_f := 3;
        ELSIF x =- 13530 THEN
            exp_f := 3;
        ELSIF x =- 13529 THEN
            exp_f := 3;
        ELSIF x =- 13528 THEN
            exp_f := 3;
        ELSIF x =- 13527 THEN
            exp_f := 3;
        ELSIF x =- 13526 THEN
            exp_f := 3;
        ELSIF x =- 13525 THEN
            exp_f := 3;
        ELSIF x =- 13524 THEN
            exp_f := 3;
        ELSIF x =- 13523 THEN
            exp_f := 3;
        ELSIF x =- 13522 THEN
            exp_f := 3;
        ELSIF x =- 13521 THEN
            exp_f := 3;
        ELSIF x =- 13520 THEN
            exp_f := 3;
        ELSIF x =- 13519 THEN
            exp_f := 3;
        ELSIF x =- 13518 THEN
            exp_f := 3;
        ELSIF x =- 13517 THEN
            exp_f := 3;
        ELSIF x =- 13516 THEN
            exp_f := 3;
        ELSIF x =- 13515 THEN
            exp_f := 3;
        ELSIF x =- 13514 THEN
            exp_f := 3;
        ELSIF x =- 13513 THEN
            exp_f := 3;
        ELSIF x =- 13512 THEN
            exp_f := 3;
        ELSIF x =- 13511 THEN
            exp_f := 3;
        ELSIF x =- 13510 THEN
            exp_f := 3;
        ELSIF x =- 13509 THEN
            exp_f := 3;
        ELSIF x =- 13508 THEN
            exp_f := 3;
        ELSIF x =- 13507 THEN
            exp_f := 3;
        ELSIF x =- 13506 THEN
            exp_f := 3;
        ELSIF x =- 13505 THEN
            exp_f := 3;
        ELSIF x =- 13504 THEN
            exp_f := 3;
        ELSIF x =- 13503 THEN
            exp_f := 3;
        ELSIF x =- 13502 THEN
            exp_f := 3;
        ELSIF x =- 13501 THEN
            exp_f := 3;
        ELSIF x =- 13500 THEN
            exp_f := 3;
        ELSIF x =- 13499 THEN
            exp_f := 3;
        ELSIF x =- 13498 THEN
            exp_f := 3;
        ELSIF x =- 13497 THEN
            exp_f := 3;
        ELSIF x =- 13496 THEN
            exp_f := 3;
        ELSIF x =- 13495 THEN
            exp_f := 3;
        ELSIF x =- 13494 THEN
            exp_f := 3;
        ELSIF x =- 13493 THEN
            exp_f := 3;
        ELSIF x =- 13492 THEN
            exp_f := 3;
        ELSIF x =- 13491 THEN
            exp_f := 3;
        ELSIF x =- 13490 THEN
            exp_f := 3;
        ELSIF x =- 13489 THEN
            exp_f := 3;
        ELSIF x =- 13488 THEN
            exp_f := 3;
        ELSIF x =- 13487 THEN
            exp_f := 3;
        ELSIF x =- 13486 THEN
            exp_f := 3;
        ELSIF x =- 13485 THEN
            exp_f := 3;
        ELSIF x =- 13484 THEN
            exp_f := 3;
        ELSIF x =- 13483 THEN
            exp_f := 3;
        ELSIF x =- 13482 THEN
            exp_f := 3;
        ELSIF x =- 13481 THEN
            exp_f := 3;
        ELSIF x =- 13480 THEN
            exp_f := 3;
        ELSIF x =- 13479 THEN
            exp_f := 3;
        ELSIF x =- 13478 THEN
            exp_f := 3;
        ELSIF x =- 13477 THEN
            exp_f := 3;
        ELSIF x =- 13476 THEN
            exp_f := 3;
        ELSIF x =- 13475 THEN
            exp_f := 3;
        ELSIF x =- 13474 THEN
            exp_f := 3;
        ELSIF x =- 13473 THEN
            exp_f := 3;
        ELSIF x =- 13472 THEN
            exp_f := 3;
        ELSIF x =- 13471 THEN
            exp_f := 3;
        ELSIF x =- 13470 THEN
            exp_f := 3;
        ELSIF x =- 13469 THEN
            exp_f := 3;
        ELSIF x =- 13468 THEN
            exp_f := 3;
        ELSIF x =- 13467 THEN
            exp_f := 3;
        ELSIF x =- 13466 THEN
            exp_f := 3;
        ELSIF x =- 13465 THEN
            exp_f := 3;
        ELSIF x =- 13464 THEN
            exp_f := 3;
        ELSIF x =- 13463 THEN
            exp_f := 3;
        ELSIF x =- 13462 THEN
            exp_f := 3;
        ELSIF x =- 13461 THEN
            exp_f := 3;
        ELSIF x =- 13460 THEN
            exp_f := 3;
        ELSIF x =- 13459 THEN
            exp_f := 3;
        ELSIF x =- 13458 THEN
            exp_f := 3;
        ELSIF x =- 13457 THEN
            exp_f := 3;
        ELSIF x =- 13456 THEN
            exp_f := 3;
        ELSIF x =- 13455 THEN
            exp_f := 3;
        ELSIF x =- 13454 THEN
            exp_f := 3;
        ELSIF x =- 13453 THEN
            exp_f := 3;
        ELSIF x =- 13452 THEN
            exp_f := 3;
        ELSIF x =- 13451 THEN
            exp_f := 3;
        ELSIF x =- 13450 THEN
            exp_f := 3;
        ELSIF x =- 13449 THEN
            exp_f := 3;
        ELSIF x =- 13448 THEN
            exp_f := 3;
        ELSIF x =- 13447 THEN
            exp_f := 3;
        ELSIF x =- 13446 THEN
            exp_f := 3;
        ELSIF x =- 13445 THEN
            exp_f := 3;
        ELSIF x =- 13444 THEN
            exp_f := 3;
        ELSIF x =- 13443 THEN
            exp_f := 3;
        ELSIF x =- 13442 THEN
            exp_f := 3;
        ELSIF x =- 13441 THEN
            exp_f := 3;
        ELSIF x =- 13440 THEN
            exp_f := 3;
        ELSIF x =- 13439 THEN
            exp_f := 3;
        ELSIF x =- 13438 THEN
            exp_f := 3;
        ELSIF x =- 13437 THEN
            exp_f := 3;
        ELSIF x =- 13436 THEN
            exp_f := 3;
        ELSIF x =- 13435 THEN
            exp_f := 3;
        ELSIF x =- 13434 THEN
            exp_f := 3;
        ELSIF x =- 13433 THEN
            exp_f := 3;
        ELSIF x =- 13432 THEN
            exp_f := 3;
        ELSIF x =- 13431 THEN
            exp_f := 3;
        ELSIF x =- 13430 THEN
            exp_f := 3;
        ELSIF x =- 13429 THEN
            exp_f := 3;
        ELSIF x =- 13428 THEN
            exp_f := 3;
        ELSIF x =- 13427 THEN
            exp_f := 3;
        ELSIF x =- 13426 THEN
            exp_f := 3;
        ELSIF x =- 13425 THEN
            exp_f := 3;
        ELSIF x =- 13424 THEN
            exp_f := 3;
        ELSIF x =- 13423 THEN
            exp_f := 3;
        ELSIF x =- 13422 THEN
            exp_f := 3;
        ELSIF x =- 13421 THEN
            exp_f := 3;
        ELSIF x =- 13420 THEN
            exp_f := 3;
        ELSIF x =- 13419 THEN
            exp_f := 3;
        ELSIF x =- 13418 THEN
            exp_f := 3;
        ELSIF x =- 13417 THEN
            exp_f := 3;
        ELSIF x =- 13416 THEN
            exp_f := 3;
        ELSIF x =- 13415 THEN
            exp_f := 3;
        ELSIF x =- 13414 THEN
            exp_f := 3;
        ELSIF x =- 13413 THEN
            exp_f := 3;
        ELSIF x =- 13412 THEN
            exp_f := 3;
        ELSIF x =- 13411 THEN
            exp_f := 3;
        ELSIF x =- 13410 THEN
            exp_f := 3;
        ELSIF x =- 13409 THEN
            exp_f := 3;
        ELSIF x =- 13408 THEN
            exp_f := 3;
        ELSIF x =- 13407 THEN
            exp_f := 3;
        ELSIF x =- 13406 THEN
            exp_f := 3;
        ELSIF x =- 13405 THEN
            exp_f := 3;
        ELSIF x =- 13404 THEN
            exp_f := 3;
        ELSIF x =- 13403 THEN
            exp_f := 3;
        ELSIF x =- 13402 THEN
            exp_f := 3;
        ELSIF x =- 13401 THEN
            exp_f := 3;
        ELSIF x =- 13400 THEN
            exp_f := 3;
        ELSIF x =- 13399 THEN
            exp_f := 3;
        ELSIF x =- 13398 THEN
            exp_f := 3;
        ELSIF x =- 13397 THEN
            exp_f := 3;
        ELSIF x =- 13396 THEN
            exp_f := 3;
        ELSIF x =- 13395 THEN
            exp_f := 3;
        ELSIF x =- 13394 THEN
            exp_f := 3;
        ELSIF x =- 13393 THEN
            exp_f := 3;
        ELSIF x =- 13392 THEN
            exp_f := 3;
        ELSIF x =- 13391 THEN
            exp_f := 3;
        ELSIF x =- 13390 THEN
            exp_f := 3;
        ELSIF x =- 13389 THEN
            exp_f := 3;
        ELSIF x =- 13388 THEN
            exp_f := 3;
        ELSIF x =- 13387 THEN
            exp_f := 3;
        ELSIF x =- 13386 THEN
            exp_f := 3;
        ELSIF x =- 13385 THEN
            exp_f := 3;
        ELSIF x =- 13384 THEN
            exp_f := 3;
        ELSIF x =- 13383 THEN
            exp_f := 3;
        ELSIF x =- 13382 THEN
            exp_f := 3;
        ELSIF x =- 13381 THEN
            exp_f := 3;
        ELSIF x =- 13380 THEN
            exp_f := 3;
        ELSIF x =- 13379 THEN
            exp_f := 3;
        ELSIF x =- 13378 THEN
            exp_f := 3;
        ELSIF x =- 13377 THEN
            exp_f := 3;
        ELSIF x =- 13376 THEN
            exp_f := 3;
        ELSIF x =- 13375 THEN
            exp_f := 3;
        ELSIF x =- 13374 THEN
            exp_f := 3;
        ELSIF x =- 13373 THEN
            exp_f := 3;
        ELSIF x =- 13372 THEN
            exp_f := 3;
        ELSIF x =- 13371 THEN
            exp_f := 3;
        ELSIF x =- 13370 THEN
            exp_f := 3;
        ELSIF x =- 13369 THEN
            exp_f := 3;
        ELSIF x =- 13368 THEN
            exp_f := 3;
        ELSIF x =- 13367 THEN
            exp_f := 3;
        ELSIF x =- 13366 THEN
            exp_f := 3;
        ELSIF x =- 13365 THEN
            exp_f := 3;
        ELSIF x =- 13364 THEN
            exp_f := 3;
        ELSIF x =- 13363 THEN
            exp_f := 3;
        ELSIF x =- 13362 THEN
            exp_f := 3;
        ELSIF x =- 13361 THEN
            exp_f := 3;
        ELSIF x =- 13360 THEN
            exp_f := 3;
        ELSIF x =- 13359 THEN
            exp_f := 3;
        ELSIF x =- 13358 THEN
            exp_f := 3;
        ELSIF x =- 13357 THEN
            exp_f := 3;
        ELSIF x =- 13356 THEN
            exp_f := 3;
        ELSIF x =- 13355 THEN
            exp_f := 3;
        ELSIF x =- 13354 THEN
            exp_f := 3;
        ELSIF x =- 13353 THEN
            exp_f := 3;
        ELSIF x =- 13352 THEN
            exp_f := 3;
        ELSIF x =- 13351 THEN
            exp_f := 3;
        ELSIF x =- 13350 THEN
            exp_f := 3;
        ELSIF x =- 13349 THEN
            exp_f := 3;
        ELSIF x =- 13348 THEN
            exp_f := 3;
        ELSIF x =- 13347 THEN
            exp_f := 3;
        ELSIF x =- 13346 THEN
            exp_f := 3;
        ELSIF x =- 13345 THEN
            exp_f := 3;
        ELSIF x =- 13344 THEN
            exp_f := 3;
        ELSIF x =- 13343 THEN
            exp_f := 3;
        ELSIF x =- 13342 THEN
            exp_f := 3;
        ELSIF x =- 13341 THEN
            exp_f := 3;
        ELSIF x =- 13340 THEN
            exp_f := 3;
        ELSIF x =- 13339 THEN
            exp_f := 3;
        ELSIF x =- 13338 THEN
            exp_f := 3;
        ELSIF x =- 13337 THEN
            exp_f := 3;
        ELSIF x =- 13336 THEN
            exp_f := 3;
        ELSIF x =- 13335 THEN
            exp_f := 3;
        ELSIF x =- 13334 THEN
            exp_f := 3;
        ELSIF x =- 13333 THEN
            exp_f := 3;
        ELSIF x =- 13332 THEN
            exp_f := 3;
        ELSIF x =- 13331 THEN
            exp_f := 3;
        ELSIF x =- 13330 THEN
            exp_f := 3;
        ELSIF x =- 13329 THEN
            exp_f := 3;
        ELSIF x =- 13328 THEN
            exp_f := 3;
        ELSIF x =- 13327 THEN
            exp_f := 3;
        ELSIF x =- 13326 THEN
            exp_f := 3;
        ELSIF x =- 13325 THEN
            exp_f := 3;
        ELSIF x =- 13324 THEN
            exp_f := 3;
        ELSIF x =- 13323 THEN
            exp_f := 3;
        ELSIF x =- 13322 THEN
            exp_f := 3;
        ELSIF x =- 13321 THEN
            exp_f := 3;
        ELSIF x =- 13320 THEN
            exp_f := 3;
        ELSIF x =- 13319 THEN
            exp_f := 3;
        ELSIF x =- 13318 THEN
            exp_f := 3;
        ELSIF x =- 13317 THEN
            exp_f := 3;
        ELSIF x =- 13316 THEN
            exp_f := 3;
        ELSIF x =- 13315 THEN
            exp_f := 3;
        ELSIF x =- 13314 THEN
            exp_f := 3;
        ELSIF x =- 13313 THEN
            exp_f := 3;
        ELSIF x =- 13312 THEN
            exp_f := 3;
        ELSIF x =- 13311 THEN
            exp_f := 3;
        ELSIF x =- 13310 THEN
            exp_f := 3;
        ELSIF x =- 13309 THEN
            exp_f := 3;
        ELSIF x =- 13308 THEN
            exp_f := 3;
        ELSIF x =- 13307 THEN
            exp_f := 3;
        ELSIF x =- 13306 THEN
            exp_f := 3;
        ELSIF x =- 13305 THEN
            exp_f := 3;
        ELSIF x =- 13304 THEN
            exp_f := 3;
        ELSIF x =- 13303 THEN
            exp_f := 3;
        ELSIF x =- 13302 THEN
            exp_f := 3;
        ELSIF x =- 13301 THEN
            exp_f := 3;
        ELSIF x =- 13300 THEN
            exp_f := 3;
        ELSIF x =- 13299 THEN
            exp_f := 3;
        ELSIF x =- 13298 THEN
            exp_f := 3;
        ELSIF x =- 13297 THEN
            exp_f := 3;
        ELSIF x =- 13296 THEN
            exp_f := 3;
        ELSIF x =- 13295 THEN
            exp_f := 3;
        ELSIF x =- 13294 THEN
            exp_f := 3;
        ELSIF x =- 13293 THEN
            exp_f := 3;
        ELSIF x =- 13292 THEN
            exp_f := 3;
        ELSIF x =- 13291 THEN
            exp_f := 3;
        ELSIF x =- 13290 THEN
            exp_f := 3;
        ELSIF x =- 13289 THEN
            exp_f := 3;
        ELSIF x =- 13288 THEN
            exp_f := 3;
        ELSIF x =- 13287 THEN
            exp_f := 3;
        ELSIF x =- 13286 THEN
            exp_f := 3;
        ELSIF x =- 13285 THEN
            exp_f := 3;
        ELSIF x =- 13284 THEN
            exp_f := 3;
        ELSIF x =- 13283 THEN
            exp_f := 3;
        ELSIF x =- 13282 THEN
            exp_f := 3;
        ELSIF x =- 13281 THEN
            exp_f := 3;
        ELSIF x =- 13280 THEN
            exp_f := 3;
        ELSIF x =- 13279 THEN
            exp_f := 3;
        ELSIF x =- 13278 THEN
            exp_f := 3;
        ELSIF x =- 13277 THEN
            exp_f := 3;
        ELSIF x =- 13276 THEN
            exp_f := 3;
        ELSIF x =- 13275 THEN
            exp_f := 3;
        ELSIF x =- 13274 THEN
            exp_f := 3;
        ELSIF x =- 13273 THEN
            exp_f := 3;
        ELSIF x =- 13272 THEN
            exp_f := 3;
        ELSIF x =- 13271 THEN
            exp_f := 3;
        ELSIF x =- 13270 THEN
            exp_f := 3;
        ELSIF x =- 13269 THEN
            exp_f := 3;
        ELSIF x =- 13268 THEN
            exp_f := 3;
        ELSIF x =- 13267 THEN
            exp_f := 3;
        ELSIF x =- 13266 THEN
            exp_f := 3;
        ELSIF x =- 13265 THEN
            exp_f := 3;
        ELSIF x =- 13264 THEN
            exp_f := 3;
        ELSIF x =- 13263 THEN
            exp_f := 3;
        ELSIF x =- 13262 THEN
            exp_f := 3;
        ELSIF x =- 13261 THEN
            exp_f := 3;
        ELSIF x =- 13260 THEN
            exp_f := 3;
        ELSIF x =- 13259 THEN
            exp_f := 3;
        ELSIF x =- 13258 THEN
            exp_f := 3;
        ELSIF x =- 13257 THEN
            exp_f := 3;
        ELSIF x =- 13256 THEN
            exp_f := 3;
        ELSIF x =- 13255 THEN
            exp_f := 3;
        ELSIF x =- 13254 THEN
            exp_f := 3;
        ELSIF x =- 13253 THEN
            exp_f := 3;
        ELSIF x =- 13252 THEN
            exp_f := 3;
        ELSIF x =- 13251 THEN
            exp_f := 3;
        ELSIF x =- 13250 THEN
            exp_f := 3;
        ELSIF x =- 13249 THEN
            exp_f := 3;
        ELSIF x =- 13248 THEN
            exp_f := 3;
        ELSIF x =- 13247 THEN
            exp_f := 3;
        ELSIF x =- 13246 THEN
            exp_f := 3;
        ELSIF x =- 13245 THEN
            exp_f := 3;
        ELSIF x =- 13244 THEN
            exp_f := 3;
        ELSIF x =- 13243 THEN
            exp_f := 3;
        ELSIF x =- 13242 THEN
            exp_f := 3;
        ELSIF x =- 13241 THEN
            exp_f := 3;
        ELSIF x =- 13240 THEN
            exp_f := 3;
        ELSIF x =- 13239 THEN
            exp_f := 3;
        ELSIF x =- 13238 THEN
            exp_f := 3;
        ELSIF x =- 13237 THEN
            exp_f := 3;
        ELSIF x =- 13236 THEN
            exp_f := 3;
        ELSIF x =- 13235 THEN
            exp_f := 3;
        ELSIF x =- 13234 THEN
            exp_f := 3;
        ELSIF x =- 13233 THEN
            exp_f := 3;
        ELSIF x =- 13232 THEN
            exp_f := 3;
        ELSIF x =- 13231 THEN
            exp_f := 3;
        ELSIF x =- 13230 THEN
            exp_f := 3;
        ELSIF x =- 13229 THEN
            exp_f := 3;
        ELSIF x =- 13228 THEN
            exp_f := 3;
        ELSIF x =- 13227 THEN
            exp_f := 3;
        ELSIF x =- 13226 THEN
            exp_f := 3;
        ELSIF x =- 13225 THEN
            exp_f := 3;
        ELSIF x =- 13224 THEN
            exp_f := 3;
        ELSIF x =- 13223 THEN
            exp_f := 3;
        ELSIF x =- 13222 THEN
            exp_f := 3;
        ELSIF x =- 13221 THEN
            exp_f := 3;
        ELSIF x =- 13220 THEN
            exp_f := 3;
        ELSIF x =- 13219 THEN
            exp_f := 3;
        ELSIF x =- 13218 THEN
            exp_f := 3;
        ELSIF x =- 13217 THEN
            exp_f := 3;
        ELSIF x =- 13216 THEN
            exp_f := 3;
        ELSIF x =- 13215 THEN
            exp_f := 3;
        ELSIF x =- 13214 THEN
            exp_f := 3;
        ELSIF x =- 13213 THEN
            exp_f := 3;
        ELSIF x =- 13212 THEN
            exp_f := 3;
        ELSIF x =- 13211 THEN
            exp_f := 3;
        ELSIF x =- 13210 THEN
            exp_f := 3;
        ELSIF x =- 13209 THEN
            exp_f := 3;
        ELSIF x =- 13208 THEN
            exp_f := 3;
        ELSIF x =- 13207 THEN
            exp_f := 3;
        ELSIF x =- 13206 THEN
            exp_f := 3;
        ELSIF x =- 13205 THEN
            exp_f := 3;
        ELSIF x =- 13204 THEN
            exp_f := 3;
        ELSIF x =- 13203 THEN
            exp_f := 3;
        ELSIF x =- 13202 THEN
            exp_f := 3;
        ELSIF x =- 13201 THEN
            exp_f := 3;
        ELSIF x =- 13200 THEN
            exp_f := 3;
        ELSIF x =- 13199 THEN
            exp_f := 3;
        ELSIF x =- 13198 THEN
            exp_f := 3;
        ELSIF x =- 13197 THEN
            exp_f := 3;
        ELSIF x =- 13196 THEN
            exp_f := 3;
        ELSIF x =- 13195 THEN
            exp_f := 3;
        ELSIF x =- 13194 THEN
            exp_f := 3;
        ELSIF x =- 13193 THEN
            exp_f := 3;
        ELSIF x =- 13192 THEN
            exp_f := 3;
        ELSIF x =- 13191 THEN
            exp_f := 3;
        ELSIF x =- 13190 THEN
            exp_f := 3;
        ELSIF x =- 13189 THEN
            exp_f := 3;
        ELSIF x =- 13188 THEN
            exp_f := 3;
        ELSIF x =- 13187 THEN
            exp_f := 3;
        ELSIF x =- 13186 THEN
            exp_f := 3;
        ELSIF x =- 13185 THEN
            exp_f := 3;
        ELSIF x =- 13184 THEN
            exp_f := 3;
        ELSIF x =- 13183 THEN
            exp_f := 3;
        ELSIF x =- 13182 THEN
            exp_f := 3;
        ELSIF x =- 13181 THEN
            exp_f := 3;
        ELSIF x =- 13180 THEN
            exp_f := 3;
        ELSIF x =- 13179 THEN
            exp_f := 3;
        ELSIF x =- 13178 THEN
            exp_f := 3;
        ELSIF x =- 13177 THEN
            exp_f := 3;
        ELSIF x =- 13176 THEN
            exp_f := 3;
        ELSIF x =- 13175 THEN
            exp_f := 3;
        ELSIF x =- 13174 THEN
            exp_f := 3;
        ELSIF x =- 13173 THEN
            exp_f := 3;
        ELSIF x =- 13172 THEN
            exp_f := 3;
        ELSIF x =- 13171 THEN
            exp_f := 3;
        ELSIF x =- 13170 THEN
            exp_f := 3;
        ELSIF x =- 13169 THEN
            exp_f := 3;
        ELSIF x =- 13168 THEN
            exp_f := 3;
        ELSIF x =- 13167 THEN
            exp_f := 3;
        ELSIF x =- 13166 THEN
            exp_f := 3;
        ELSIF x =- 13165 THEN
            exp_f := 3;
        ELSIF x =- 13164 THEN
            exp_f := 3;
        ELSIF x =- 13163 THEN
            exp_f := 3;
        ELSIF x =- 13162 THEN
            exp_f := 3;
        ELSIF x =- 13161 THEN
            exp_f := 3;
        ELSIF x =- 13160 THEN
            exp_f := 3;
        ELSIF x =- 13159 THEN
            exp_f := 3;
        ELSIF x =- 13158 THEN
            exp_f := 3;
        ELSIF x =- 13157 THEN
            exp_f := 3;
        ELSIF x =- 13156 THEN
            exp_f := 3;
        ELSIF x =- 13155 THEN
            exp_f := 3;
        ELSIF x =- 13154 THEN
            exp_f := 3;
        ELSIF x =- 13153 THEN
            exp_f := 3;
        ELSIF x =- 13152 THEN
            exp_f := 3;
        ELSIF x =- 13151 THEN
            exp_f := 3;
        ELSIF x =- 13150 THEN
            exp_f := 3;
        ELSIF x =- 13149 THEN
            exp_f := 3;
        ELSIF x =- 13148 THEN
            exp_f := 3;
        ELSIF x =- 13147 THEN
            exp_f := 3;
        ELSIF x =- 13146 THEN
            exp_f := 3;
        ELSIF x =- 13145 THEN
            exp_f := 3;
        ELSIF x =- 13144 THEN
            exp_f := 3;
        ELSIF x =- 13143 THEN
            exp_f := 3;
        ELSIF x =- 13142 THEN
            exp_f := 3;
        ELSIF x =- 13141 THEN
            exp_f := 3;
        ELSIF x =- 13140 THEN
            exp_f := 3;
        ELSIF x =- 13139 THEN
            exp_f := 3;
        ELSIF x =- 13138 THEN
            exp_f := 3;
        ELSIF x =- 13137 THEN
            exp_f := 3;
        ELSIF x =- 13136 THEN
            exp_f := 3;
        ELSIF x =- 13135 THEN
            exp_f := 3;
        ELSIF x =- 13134 THEN
            exp_f := 3;
        ELSIF x =- 13133 THEN
            exp_f := 3;
        ELSIF x =- 13132 THEN
            exp_f := 3;
        ELSIF x =- 13131 THEN
            exp_f := 3;
        ELSIF x =- 13130 THEN
            exp_f := 3;
        ELSIF x =- 13129 THEN
            exp_f := 3;
        ELSIF x =- 13128 THEN
            exp_f := 3;
        ELSIF x =- 13127 THEN
            exp_f := 3;
        ELSIF x =- 13126 THEN
            exp_f := 3;
        ELSIF x =- 13125 THEN
            exp_f := 3;
        ELSIF x =- 13124 THEN
            exp_f := 3;
        ELSIF x =- 13123 THEN
            exp_f := 3;
        ELSIF x =- 13122 THEN
            exp_f := 3;
        ELSIF x =- 13121 THEN
            exp_f := 3;
        ELSIF x =- 13120 THEN
            exp_f := 3;
        ELSIF x =- 13119 THEN
            exp_f := 3;
        ELSIF x =- 13118 THEN
            exp_f := 3;
        ELSIF x =- 13117 THEN
            exp_f := 3;
        ELSIF x =- 13116 THEN
            exp_f := 3;
        ELSIF x =- 13115 THEN
            exp_f := 3;
        ELSIF x =- 13114 THEN
            exp_f := 3;
        ELSIF x =- 13113 THEN
            exp_f := 3;
        ELSIF x =- 13112 THEN
            exp_f := 3;
        ELSIF x =- 13111 THEN
            exp_f := 3;
        ELSIF x =- 13110 THEN
            exp_f := 3;
        ELSIF x =- 13109 THEN
            exp_f := 3;
        ELSIF x =- 13108 THEN
            exp_f := 3;
        ELSIF x =- 13107 THEN
            exp_f := 3;
        ELSIF x =- 13106 THEN
            exp_f := 3;
        ELSIF x =- 13105 THEN
            exp_f := 3;
        ELSIF x =- 13104 THEN
            exp_f := 3;
        ELSIF x =- 13103 THEN
            exp_f := 3;
        ELSIF x =- 13102 THEN
            exp_f := 3;
        ELSIF x =- 13101 THEN
            exp_f := 3;
        ELSIF x =- 13100 THEN
            exp_f := 3;
        ELSIF x =- 13099 THEN
            exp_f := 3;
        ELSIF x =- 13098 THEN
            exp_f := 3;
        ELSIF x =- 13097 THEN
            exp_f := 3;
        ELSIF x =- 13096 THEN
            exp_f := 3;
        ELSIF x =- 13095 THEN
            exp_f := 3;
        ELSIF x =- 13094 THEN
            exp_f := 3;
        ELSIF x =- 13093 THEN
            exp_f := 3;
        ELSIF x =- 13092 THEN
            exp_f := 3;
        ELSIF x =- 13091 THEN
            exp_f := 3;
        ELSIF x =- 13090 THEN
            exp_f := 3;
        ELSIF x =- 13089 THEN
            exp_f := 3;
        ELSIF x =- 13088 THEN
            exp_f := 3;
        ELSIF x =- 13087 THEN
            exp_f := 3;
        ELSIF x =- 13086 THEN
            exp_f := 3;
        ELSIF x =- 13085 THEN
            exp_f := 3;
        ELSIF x =- 13084 THEN
            exp_f := 3;
        ELSIF x =- 13083 THEN
            exp_f := 3;
        ELSIF x =- 13082 THEN
            exp_f := 3;
        ELSIF x =- 13081 THEN
            exp_f := 3;
        ELSIF x =- 13080 THEN
            exp_f := 3;
        ELSIF x =- 13079 THEN
            exp_f := 3;
        ELSIF x =- 13078 THEN
            exp_f := 3;
        ELSIF x =- 13077 THEN
            exp_f := 3;
        ELSIF x =- 13076 THEN
            exp_f := 3;
        ELSIF x =- 13075 THEN
            exp_f := 3;
        ELSIF x =- 13074 THEN
            exp_f := 3;
        ELSIF x =- 13073 THEN
            exp_f := 3;
        ELSIF x =- 13072 THEN
            exp_f := 3;
        ELSIF x =- 13071 THEN
            exp_f := 3;
        ELSIF x =- 13070 THEN
            exp_f := 3;
        ELSIF x =- 13069 THEN
            exp_f := 3;
        ELSIF x =- 13068 THEN
            exp_f := 3;
        ELSIF x =- 13067 THEN
            exp_f := 3;
        ELSIF x =- 13066 THEN
            exp_f := 3;
        ELSIF x =- 13065 THEN
            exp_f := 3;
        ELSIF x =- 13064 THEN
            exp_f := 3;
        ELSIF x =- 13063 THEN
            exp_f := 3;
        ELSIF x =- 13062 THEN
            exp_f := 3;
        ELSIF x =- 13061 THEN
            exp_f := 3;
        ELSIF x =- 13060 THEN
            exp_f := 3;
        ELSIF x =- 13059 THEN
            exp_f := 3;
        ELSIF x =- 13058 THEN
            exp_f := 3;
        ELSIF x =- 13057 THEN
            exp_f := 3;
        ELSIF x =- 13056 THEN
            exp_f := 3;
        ELSIF x =- 13055 THEN
            exp_f := 3;
        ELSIF x =- 13054 THEN
            exp_f := 3;
        ELSIF x =- 13053 THEN
            exp_f := 3;
        ELSIF x =- 13052 THEN
            exp_f := 3;
        ELSIF x =- 13051 THEN
            exp_f := 3;
        ELSIF x =- 13050 THEN
            exp_f := 3;
        ELSIF x =- 13049 THEN
            exp_f := 3;
        ELSIF x =- 13048 THEN
            exp_f := 3;
        ELSIF x =- 13047 THEN
            exp_f := 3;
        ELSIF x =- 13046 THEN
            exp_f := 3;
        ELSIF x =- 13045 THEN
            exp_f := 3;
        ELSIF x =- 13044 THEN
            exp_f := 3;
        ELSIF x =- 13043 THEN
            exp_f := 3;
        ELSIF x =- 13042 THEN
            exp_f := 3;
        ELSIF x =- 13041 THEN
            exp_f := 3;
        ELSIF x =- 13040 THEN
            exp_f := 3;
        ELSIF x =- 13039 THEN
            exp_f := 3;
        ELSIF x =- 13038 THEN
            exp_f := 3;
        ELSIF x =- 13037 THEN
            exp_f := 3;
        ELSIF x =- 13036 THEN
            exp_f := 3;
        ELSIF x =- 13035 THEN
            exp_f := 3;
        ELSIF x =- 13034 THEN
            exp_f := 3;
        ELSIF x =- 13033 THEN
            exp_f := 3;
        ELSIF x =- 13032 THEN
            exp_f := 3;
        ELSIF x =- 13031 THEN
            exp_f := 3;
        ELSIF x =- 13030 THEN
            exp_f := 3;
        ELSIF x =- 13029 THEN
            exp_f := 3;
        ELSIF x =- 13028 THEN
            exp_f := 3;
        ELSIF x =- 13027 THEN
            exp_f := 3;
        ELSIF x =- 13026 THEN
            exp_f := 3;
        ELSIF x =- 13025 THEN
            exp_f := 3;
        ELSIF x =- 13024 THEN
            exp_f := 3;
        ELSIF x =- 13023 THEN
            exp_f := 3;
        ELSIF x =- 13022 THEN
            exp_f := 3;
        ELSIF x =- 13021 THEN
            exp_f := 3;
        ELSIF x =- 13020 THEN
            exp_f := 3;
        ELSIF x =- 13019 THEN
            exp_f := 3;
        ELSIF x =- 13018 THEN
            exp_f := 3;
        ELSIF x =- 13017 THEN
            exp_f := 3;
        ELSIF x =- 13016 THEN
            exp_f := 3;
        ELSIF x =- 13015 THEN
            exp_f := 3;
        ELSIF x =- 13014 THEN
            exp_f := 3;
        ELSIF x =- 13013 THEN
            exp_f := 3;
        ELSIF x =- 13012 THEN
            exp_f := 3;
        ELSIF x =- 13011 THEN
            exp_f := 3;
        ELSIF x =- 13010 THEN
            exp_f := 3;
        ELSIF x =- 13009 THEN
            exp_f := 3;
        ELSIF x =- 13008 THEN
            exp_f := 3;
        ELSIF x =- 13007 THEN
            exp_f := 3;
        ELSIF x =- 13006 THEN
            exp_f := 3;
        ELSIF x =- 13005 THEN
            exp_f := 3;
        ELSIF x =- 13004 THEN
            exp_f := 3;
        ELSIF x =- 13003 THEN
            exp_f := 3;
        ELSIF x =- 13002 THEN
            exp_f := 3;
        ELSIF x =- 13001 THEN
            exp_f := 3;
        ELSIF x =- 13000 THEN
            exp_f := 3;
        ELSIF x =- 12999 THEN
            exp_f := 3;
        ELSIF x =- 12998 THEN
            exp_f := 3;
        ELSIF x =- 12997 THEN
            exp_f := 3;
        ELSIF x =- 12996 THEN
            exp_f := 3;
        ELSIF x =- 12995 THEN
            exp_f := 3;
        ELSIF x =- 12994 THEN
            exp_f := 3;
        ELSIF x =- 12993 THEN
            exp_f := 3;
        ELSIF x =- 12992 THEN
            exp_f := 3;
        ELSIF x =- 12991 THEN
            exp_f := 3;
        ELSIF x =- 12990 THEN
            exp_f := 3;
        ELSIF x =- 12989 THEN
            exp_f := 3;
        ELSIF x =- 12988 THEN
            exp_f := 3;
        ELSIF x =- 12987 THEN
            exp_f := 3;
        ELSIF x =- 12986 THEN
            exp_f := 3;
        ELSIF x =- 12985 THEN
            exp_f := 3;
        ELSIF x =- 12984 THEN
            exp_f := 3;
        ELSIF x =- 12983 THEN
            exp_f := 3;
        ELSIF x =- 12982 THEN
            exp_f := 3;
        ELSIF x =- 12981 THEN
            exp_f := 3;
        ELSIF x =- 12980 THEN
            exp_f := 3;
        ELSIF x =- 12979 THEN
            exp_f := 3;
        ELSIF x =- 12978 THEN
            exp_f := 3;
        ELSIF x =- 12977 THEN
            exp_f := 3;
        ELSIF x =- 12976 THEN
            exp_f := 3;
        ELSIF x =- 12975 THEN
            exp_f := 3;
        ELSIF x =- 12974 THEN
            exp_f := 3;
        ELSIF x =- 12973 THEN
            exp_f := 3;
        ELSIF x =- 12972 THEN
            exp_f := 3;
        ELSIF x =- 12971 THEN
            exp_f := 3;
        ELSIF x =- 12970 THEN
            exp_f := 3;
        ELSIF x =- 12969 THEN
            exp_f := 3;
        ELSIF x =- 12968 THEN
            exp_f := 3;
        ELSIF x =- 12967 THEN
            exp_f := 3;
        ELSIF x =- 12966 THEN
            exp_f := 3;
        ELSIF x =- 12965 THEN
            exp_f := 3;
        ELSIF x =- 12964 THEN
            exp_f := 3;
        ELSIF x =- 12963 THEN
            exp_f := 3;
        ELSIF x =- 12962 THEN
            exp_f := 3;
        ELSIF x =- 12961 THEN
            exp_f := 3;
        ELSIF x =- 12960 THEN
            exp_f := 3;
        ELSIF x =- 12959 THEN
            exp_f := 3;
        ELSIF x =- 12958 THEN
            exp_f := 3;
        ELSIF x =- 12957 THEN
            exp_f := 3;
        ELSIF x =- 12956 THEN
            exp_f := 3;
        ELSIF x =- 12955 THEN
            exp_f := 3;
        ELSIF x =- 12954 THEN
            exp_f := 3;
        ELSIF x =- 12953 THEN
            exp_f := 3;
        ELSIF x =- 12952 THEN
            exp_f := 3;
        ELSIF x =- 12951 THEN
            exp_f := 3;
        ELSIF x =- 12950 THEN
            exp_f := 3;
        ELSIF x =- 12949 THEN
            exp_f := 3;
        ELSIF x =- 12948 THEN
            exp_f := 3;
        ELSIF x =- 12947 THEN
            exp_f := 3;
        ELSIF x =- 12946 THEN
            exp_f := 3;
        ELSIF x =- 12945 THEN
            exp_f := 3;
        ELSIF x =- 12944 THEN
            exp_f := 3;
        ELSIF x =- 12943 THEN
            exp_f := 3;
        ELSIF x =- 12942 THEN
            exp_f := 3;
        ELSIF x =- 12941 THEN
            exp_f := 3;
        ELSIF x =- 12940 THEN
            exp_f := 3;
        ELSIF x =- 12939 THEN
            exp_f := 3;
        ELSIF x =- 12938 THEN
            exp_f := 3;
        ELSIF x =- 12937 THEN
            exp_f := 3;
        ELSIF x =- 12936 THEN
            exp_f := 3;
        ELSIF x =- 12935 THEN
            exp_f := 3;
        ELSIF x =- 12934 THEN
            exp_f := 3;
        ELSIF x =- 12933 THEN
            exp_f := 3;
        ELSIF x =- 12932 THEN
            exp_f := 3;
        ELSIF x =- 12931 THEN
            exp_f := 3;
        ELSIF x =- 12930 THEN
            exp_f := 3;
        ELSIF x =- 12929 THEN
            exp_f := 3;
        ELSIF x =- 12928 THEN
            exp_f := 3;
        ELSIF x =- 12927 THEN
            exp_f := 3;
        ELSIF x =- 12926 THEN
            exp_f := 3;
        ELSIF x =- 12925 THEN
            exp_f := 3;
        ELSIF x =- 12924 THEN
            exp_f := 3;
        ELSIF x =- 12923 THEN
            exp_f := 3;
        ELSIF x =- 12922 THEN
            exp_f := 3;
        ELSIF x =- 12921 THEN
            exp_f := 3;
        ELSIF x =- 12920 THEN
            exp_f := 3;
        ELSIF x =- 12919 THEN
            exp_f := 3;
        ELSIF x =- 12918 THEN
            exp_f := 3;
        ELSIF x =- 12917 THEN
            exp_f := 3;
        ELSIF x =- 12916 THEN
            exp_f := 3;
        ELSIF x =- 12915 THEN
            exp_f := 3;
        ELSIF x =- 12914 THEN
            exp_f := 3;
        ELSIF x =- 12913 THEN
            exp_f := 3;
        ELSIF x =- 12912 THEN
            exp_f := 3;
        ELSIF x =- 12911 THEN
            exp_f := 3;
        ELSIF x =- 12910 THEN
            exp_f := 3;
        ELSIF x =- 12909 THEN
            exp_f := 3;
        ELSIF x =- 12908 THEN
            exp_f := 3;
        ELSIF x =- 12907 THEN
            exp_f := 3;
        ELSIF x =- 12906 THEN
            exp_f := 3;
        ELSIF x =- 12905 THEN
            exp_f := 3;
        ELSIF x =- 12904 THEN
            exp_f := 3;
        ELSIF x =- 12903 THEN
            exp_f := 3;
        ELSIF x =- 12902 THEN
            exp_f := 3;
        ELSIF x =- 12901 THEN
            exp_f := 3;
        ELSIF x =- 12900 THEN
            exp_f := 3;
        ELSIF x =- 12899 THEN
            exp_f := 3;
        ELSIF x =- 12898 THEN
            exp_f := 3;
        ELSIF x =- 12897 THEN
            exp_f := 3;
        ELSIF x =- 12896 THEN
            exp_f := 3;
        ELSIF x =- 12895 THEN
            exp_f := 3;
        ELSIF x =- 12894 THEN
            exp_f := 3;
        ELSIF x =- 12893 THEN
            exp_f := 3;
        ELSIF x =- 12892 THEN
            exp_f := 3;
        ELSIF x =- 12891 THEN
            exp_f := 3;
        ELSIF x =- 12890 THEN
            exp_f := 3;
        ELSIF x =- 12889 THEN
            exp_f := 3;
        ELSIF x =- 12888 THEN
            exp_f := 3;
        ELSIF x =- 12887 THEN
            exp_f := 3;
        ELSIF x =- 12886 THEN
            exp_f := 3;
        ELSIF x =- 12885 THEN
            exp_f := 3;
        ELSIF x =- 12884 THEN
            exp_f := 3;
        ELSIF x =- 12883 THEN
            exp_f := 3;
        ELSIF x =- 12882 THEN
            exp_f := 3;
        ELSIF x =- 12881 THEN
            exp_f := 3;
        ELSIF x =- 12880 THEN
            exp_f := 3;
        ELSIF x =- 12879 THEN
            exp_f := 3;
        ELSIF x =- 12878 THEN
            exp_f := 3;
        ELSIF x =- 12877 THEN
            exp_f := 3;
        ELSIF x =- 12876 THEN
            exp_f := 3;
        ELSIF x =- 12875 THEN
            exp_f := 3;
        ELSIF x =- 12874 THEN
            exp_f := 3;
        ELSIF x =- 12873 THEN
            exp_f := 3;
        ELSIF x =- 12872 THEN
            exp_f := 3;
        ELSIF x =- 12871 THEN
            exp_f := 3;
        ELSIF x =- 12870 THEN
            exp_f := 3;
        ELSIF x =- 12869 THEN
            exp_f := 3;
        ELSIF x =- 12868 THEN
            exp_f := 3;
        ELSIF x =- 12867 THEN
            exp_f := 3;
        ELSIF x =- 12866 THEN
            exp_f := 3;
        ELSIF x =- 12865 THEN
            exp_f := 3;
        ELSIF x =- 12864 THEN
            exp_f := 3;
        ELSIF x =- 12863 THEN
            exp_f := 3;
        ELSIF x =- 12862 THEN
            exp_f := 3;
        ELSIF x =- 12861 THEN
            exp_f := 3;
        ELSIF x =- 12860 THEN
            exp_f := 3;
        ELSIF x =- 12859 THEN
            exp_f := 3;
        ELSIF x =- 12858 THEN
            exp_f := 3;
        ELSIF x =- 12857 THEN
            exp_f := 3;
        ELSIF x =- 12856 THEN
            exp_f := 3;
        ELSIF x =- 12855 THEN
            exp_f := 3;
        ELSIF x =- 12854 THEN
            exp_f := 3;
        ELSIF x =- 12853 THEN
            exp_f := 3;
        ELSIF x =- 12852 THEN
            exp_f := 3;
        ELSIF x =- 12851 THEN
            exp_f := 3;
        ELSIF x =- 12850 THEN
            exp_f := 3;
        ELSIF x =- 12849 THEN
            exp_f := 3;
        ELSIF x =- 12848 THEN
            exp_f := 3;
        ELSIF x =- 12847 THEN
            exp_f := 3;
        ELSIF x =- 12846 THEN
            exp_f := 3;
        ELSIF x =- 12845 THEN
            exp_f := 3;
        ELSIF x =- 12844 THEN
            exp_f := 3;
        ELSIF x =- 12843 THEN
            exp_f := 3;
        ELSIF x =- 12842 THEN
            exp_f := 3;
        ELSIF x =- 12841 THEN
            exp_f := 3;
        ELSIF x =- 12840 THEN
            exp_f := 3;
        ELSIF x =- 12839 THEN
            exp_f := 3;
        ELSIF x =- 12838 THEN
            exp_f := 3;
        ELSIF x =- 12837 THEN
            exp_f := 3;
        ELSIF x =- 12836 THEN
            exp_f := 3;
        ELSIF x =- 12835 THEN
            exp_f := 3;
        ELSIF x =- 12834 THEN
            exp_f := 3;
        ELSIF x =- 12833 THEN
            exp_f := 3;
        ELSIF x =- 12832 THEN
            exp_f := 3;
        ELSIF x =- 12831 THEN
            exp_f := 3;
        ELSIF x =- 12830 THEN
            exp_f := 3;
        ELSIF x =- 12829 THEN
            exp_f := 3;
        ELSIF x =- 12828 THEN
            exp_f := 3;
        ELSIF x =- 12827 THEN
            exp_f := 3;
        ELSIF x =- 12826 THEN
            exp_f := 3;
        ELSIF x =- 12825 THEN
            exp_f := 3;
        ELSIF x =- 12824 THEN
            exp_f := 3;
        ELSIF x =- 12823 THEN
            exp_f := 3;
        ELSIF x =- 12822 THEN
            exp_f := 3;
        ELSIF x =- 12821 THEN
            exp_f := 3;
        ELSIF x =- 12820 THEN
            exp_f := 3;
        ELSIF x =- 12819 THEN
            exp_f := 3;
        ELSIF x =- 12818 THEN
            exp_f := 3;
        ELSIF x =- 12817 THEN
            exp_f := 3;
        ELSIF x =- 12816 THEN
            exp_f := 3;
        ELSIF x =- 12815 THEN
            exp_f := 3;
        ELSIF x =- 12814 THEN
            exp_f := 3;
        ELSIF x =- 12813 THEN
            exp_f := 3;
        ELSIF x =- 12812 THEN
            exp_f := 3;
        ELSIF x =- 12811 THEN
            exp_f := 3;
        ELSIF x =- 12810 THEN
            exp_f := 3;
        ELSIF x =- 12809 THEN
            exp_f := 3;
        ELSIF x =- 12808 THEN
            exp_f := 3;
        ELSIF x =- 12807 THEN
            exp_f := 3;
        ELSIF x =- 12806 THEN
            exp_f := 3;
        ELSIF x =- 12805 THEN
            exp_f := 3;
        ELSIF x =- 12804 THEN
            exp_f := 3;
        ELSIF x =- 12803 THEN
            exp_f := 3;
        ELSIF x =- 12802 THEN
            exp_f := 3;
        ELSIF x =- 12801 THEN
            exp_f := 3;
        ELSIF x =- 12800 THEN
            exp_f := 3;
        ELSIF x =- 12799 THEN
            exp_f := 4;
        ELSIF x =- 12798 THEN
            exp_f := 4;
        ELSIF x =- 12797 THEN
            exp_f := 4;
        ELSIF x =- 12796 THEN
            exp_f := 4;
        ELSIF x =- 12795 THEN
            exp_f := 4;
        ELSIF x =- 12794 THEN
            exp_f := 4;
        ELSIF x =- 12793 THEN
            exp_f := 4;
        ELSIF x =- 12792 THEN
            exp_f := 4;
        ELSIF x =- 12791 THEN
            exp_f := 4;
        ELSIF x =- 12790 THEN
            exp_f := 4;
        ELSIF x =- 12789 THEN
            exp_f := 4;
        ELSIF x =- 12788 THEN
            exp_f := 4;
        ELSIF x =- 12787 THEN
            exp_f := 4;
        ELSIF x =- 12786 THEN
            exp_f := 4;
        ELSIF x =- 12785 THEN
            exp_f := 4;
        ELSIF x =- 12784 THEN
            exp_f := 4;
        ELSIF x =- 12783 THEN
            exp_f := 4;
        ELSIF x =- 12782 THEN
            exp_f := 4;
        ELSIF x =- 12781 THEN
            exp_f := 4;
        ELSIF x =- 12780 THEN
            exp_f := 4;
        ELSIF x =- 12779 THEN
            exp_f := 4;
        ELSIF x =- 12778 THEN
            exp_f := 4;
        ELSIF x =- 12777 THEN
            exp_f := 4;
        ELSIF x =- 12776 THEN
            exp_f := 4;
        ELSIF x =- 12775 THEN
            exp_f := 4;
        ELSIF x =- 12774 THEN
            exp_f := 4;
        ELSIF x =- 12773 THEN
            exp_f := 4;
        ELSIF x =- 12772 THEN
            exp_f := 4;
        ELSIF x =- 12771 THEN
            exp_f := 4;
        ELSIF x =- 12770 THEN
            exp_f := 4;
        ELSIF x =- 12769 THEN
            exp_f := 4;
        ELSIF x =- 12768 THEN
            exp_f := 4;
        ELSIF x =- 12767 THEN
            exp_f := 4;
        ELSIF x =- 12766 THEN
            exp_f := 4;
        ELSIF x =- 12765 THEN
            exp_f := 4;
        ELSIF x =- 12764 THEN
            exp_f := 4;
        ELSIF x =- 12763 THEN
            exp_f := 4;
        ELSIF x =- 12762 THEN
            exp_f := 4;
        ELSIF x =- 12761 THEN
            exp_f := 4;
        ELSIF x =- 12760 THEN
            exp_f := 4;
        ELSIF x =- 12759 THEN
            exp_f := 4;
        ELSIF x =- 12758 THEN
            exp_f := 4;
        ELSIF x =- 12757 THEN
            exp_f := 4;
        ELSIF x =- 12756 THEN
            exp_f := 4;
        ELSIF x =- 12755 THEN
            exp_f := 4;
        ELSIF x =- 12754 THEN
            exp_f := 4;
        ELSIF x =- 12753 THEN
            exp_f := 4;
        ELSIF x =- 12752 THEN
            exp_f := 4;
        ELSIF x =- 12751 THEN
            exp_f := 4;
        ELSIF x =- 12750 THEN
            exp_f := 4;
        ELSIF x =- 12749 THEN
            exp_f := 4;
        ELSIF x =- 12748 THEN
            exp_f := 4;
        ELSIF x =- 12747 THEN
            exp_f := 4;
        ELSIF x =- 12746 THEN
            exp_f := 4;
        ELSIF x =- 12745 THEN
            exp_f := 4;
        ELSIF x =- 12744 THEN
            exp_f := 4;
        ELSIF x =- 12743 THEN
            exp_f := 4;
        ELSIF x =- 12742 THEN
            exp_f := 4;
        ELSIF x =- 12741 THEN
            exp_f := 4;
        ELSIF x =- 12740 THEN
            exp_f := 4;
        ELSIF x =- 12739 THEN
            exp_f := 4;
        ELSIF x =- 12738 THEN
            exp_f := 4;
        ELSIF x =- 12737 THEN
            exp_f := 4;
        ELSIF x =- 12736 THEN
            exp_f := 4;
        ELSIF x =- 12735 THEN
            exp_f := 4;
        ELSIF x =- 12734 THEN
            exp_f := 4;
        ELSIF x =- 12733 THEN
            exp_f := 4;
        ELSIF x =- 12732 THEN
            exp_f := 4;
        ELSIF x =- 12731 THEN
            exp_f := 4;
        ELSIF x =- 12730 THEN
            exp_f := 4;
        ELSIF x =- 12729 THEN
            exp_f := 4;
        ELSIF x =- 12728 THEN
            exp_f := 4;
        ELSIF x =- 12727 THEN
            exp_f := 4;
        ELSIF x =- 12726 THEN
            exp_f := 4;
        ELSIF x =- 12725 THEN
            exp_f := 4;
        ELSIF x =- 12724 THEN
            exp_f := 4;
        ELSIF x =- 12723 THEN
            exp_f := 4;
        ELSIF x =- 12722 THEN
            exp_f := 4;
        ELSIF x =- 12721 THEN
            exp_f := 4;
        ELSIF x =- 12720 THEN
            exp_f := 4;
        ELSIF x =- 12719 THEN
            exp_f := 4;
        ELSIF x =- 12718 THEN
            exp_f := 4;
        ELSIF x =- 12717 THEN
            exp_f := 4;
        ELSIF x =- 12716 THEN
            exp_f := 4;
        ELSIF x =- 12715 THEN
            exp_f := 4;
        ELSIF x =- 12714 THEN
            exp_f := 4;
        ELSIF x =- 12713 THEN
            exp_f := 4;
        ELSIF x =- 12712 THEN
            exp_f := 4;
        ELSIF x =- 12711 THEN
            exp_f := 4;
        ELSIF x =- 12710 THEN
            exp_f := 4;
        ELSIF x =- 12709 THEN
            exp_f := 4;
        ELSIF x =- 12708 THEN
            exp_f := 4;
        ELSIF x =- 12707 THEN
            exp_f := 4;
        ELSIF x =- 12706 THEN
            exp_f := 4;
        ELSIF x =- 12705 THEN
            exp_f := 4;
        ELSIF x =- 12704 THEN
            exp_f := 4;
        ELSIF x =- 12703 THEN
            exp_f := 4;
        ELSIF x =- 12702 THEN
            exp_f := 4;
        ELSIF x =- 12701 THEN
            exp_f := 4;
        ELSIF x =- 12700 THEN
            exp_f := 4;
        ELSIF x =- 12699 THEN
            exp_f := 4;
        ELSIF x =- 12698 THEN
            exp_f := 4;
        ELSIF x =- 12697 THEN
            exp_f := 4;
        ELSIF x =- 12696 THEN
            exp_f := 4;
        ELSIF x =- 12695 THEN
            exp_f := 4;
        ELSIF x =- 12694 THEN
            exp_f := 4;
        ELSIF x =- 12693 THEN
            exp_f := 4;
        ELSIF x =- 12692 THEN
            exp_f := 4;
        ELSIF x =- 12691 THEN
            exp_f := 4;
        ELSIF x =- 12690 THEN
            exp_f := 4;
        ELSIF x =- 12689 THEN
            exp_f := 4;
        ELSIF x =- 12688 THEN
            exp_f := 4;
        ELSIF x =- 12687 THEN
            exp_f := 4;
        ELSIF x =- 12686 THEN
            exp_f := 4;
        ELSIF x =- 12685 THEN
            exp_f := 4;
        ELSIF x =- 12684 THEN
            exp_f := 4;
        ELSIF x =- 12683 THEN
            exp_f := 4;
        ELSIF x =- 12682 THEN
            exp_f := 4;
        ELSIF x =- 12681 THEN
            exp_f := 4;
        ELSIF x =- 12680 THEN
            exp_f := 4;
        ELSIF x =- 12679 THEN
            exp_f := 4;
        ELSIF x =- 12678 THEN
            exp_f := 4;
        ELSIF x =- 12677 THEN
            exp_f := 4;
        ELSIF x =- 12676 THEN
            exp_f := 4;
        ELSIF x =- 12675 THEN
            exp_f := 4;
        ELSIF x =- 12674 THEN
            exp_f := 4;
        ELSIF x =- 12673 THEN
            exp_f := 4;
        ELSIF x =- 12672 THEN
            exp_f := 4;
        ELSIF x =- 12671 THEN
            exp_f := 4;
        ELSIF x =- 12670 THEN
            exp_f := 4;
        ELSIF x =- 12669 THEN
            exp_f := 4;
        ELSIF x =- 12668 THEN
            exp_f := 4;
        ELSIF x =- 12667 THEN
            exp_f := 4;
        ELSIF x =- 12666 THEN
            exp_f := 4;
        ELSIF x =- 12665 THEN
            exp_f := 4;
        ELSIF x =- 12664 THEN
            exp_f := 4;
        ELSIF x =- 12663 THEN
            exp_f := 4;
        ELSIF x =- 12662 THEN
            exp_f := 4;
        ELSIF x =- 12661 THEN
            exp_f := 4;
        ELSIF x =- 12660 THEN
            exp_f := 4;
        ELSIF x =- 12659 THEN
            exp_f := 4;
        ELSIF x =- 12658 THEN
            exp_f := 4;
        ELSIF x =- 12657 THEN
            exp_f := 4;
        ELSIF x =- 12656 THEN
            exp_f := 4;
        ELSIF x =- 12655 THEN
            exp_f := 4;
        ELSIF x =- 12654 THEN
            exp_f := 4;
        ELSIF x =- 12653 THEN
            exp_f := 4;
        ELSIF x =- 12652 THEN
            exp_f := 4;
        ELSIF x =- 12651 THEN
            exp_f := 4;
        ELSIF x =- 12650 THEN
            exp_f := 4;
        ELSIF x =- 12649 THEN
            exp_f := 4;
        ELSIF x =- 12648 THEN
            exp_f := 4;
        ELSIF x =- 12647 THEN
            exp_f := 4;
        ELSIF x =- 12646 THEN
            exp_f := 4;
        ELSIF x =- 12645 THEN
            exp_f := 4;
        ELSIF x =- 12644 THEN
            exp_f := 4;
        ELSIF x =- 12643 THEN
            exp_f := 4;
        ELSIF x =- 12642 THEN
            exp_f := 4;
        ELSIF x =- 12641 THEN
            exp_f := 4;
        ELSIF x =- 12640 THEN
            exp_f := 4;
        ELSIF x =- 12639 THEN
            exp_f := 4;
        ELSIF x =- 12638 THEN
            exp_f := 4;
        ELSIF x =- 12637 THEN
            exp_f := 4;
        ELSIF x =- 12636 THEN
            exp_f := 4;
        ELSIF x =- 12635 THEN
            exp_f := 4;
        ELSIF x =- 12634 THEN
            exp_f := 4;
        ELSIF x =- 12633 THEN
            exp_f := 4;
        ELSIF x =- 12632 THEN
            exp_f := 4;
        ELSIF x =- 12631 THEN
            exp_f := 4;
        ELSIF x =- 12630 THEN
            exp_f := 4;
        ELSIF x =- 12629 THEN
            exp_f := 4;
        ELSIF x =- 12628 THEN
            exp_f := 4;
        ELSIF x =- 12627 THEN
            exp_f := 4;
        ELSIF x =- 12626 THEN
            exp_f := 4;
        ELSIF x =- 12625 THEN
            exp_f := 4;
        ELSIF x =- 12624 THEN
            exp_f := 4;
        ELSIF x =- 12623 THEN
            exp_f := 4;
        ELSIF x =- 12622 THEN
            exp_f := 4;
        ELSIF x =- 12621 THEN
            exp_f := 4;
        ELSIF x =- 12620 THEN
            exp_f := 4;
        ELSIF x =- 12619 THEN
            exp_f := 4;
        ELSIF x =- 12618 THEN
            exp_f := 4;
        ELSIF x =- 12617 THEN
            exp_f := 4;
        ELSIF x =- 12616 THEN
            exp_f := 4;
        ELSIF x =- 12615 THEN
            exp_f := 4;
        ELSIF x =- 12614 THEN
            exp_f := 4;
        ELSIF x =- 12613 THEN
            exp_f := 4;
        ELSIF x =- 12612 THEN
            exp_f := 4;
        ELSIF x =- 12611 THEN
            exp_f := 4;
        ELSIF x =- 12610 THEN
            exp_f := 4;
        ELSIF x =- 12609 THEN
            exp_f := 4;
        ELSIF x =- 12608 THEN
            exp_f := 4;
        ELSIF x =- 12607 THEN
            exp_f := 4;
        ELSIF x =- 12606 THEN
            exp_f := 4;
        ELSIF x =- 12605 THEN
            exp_f := 4;
        ELSIF x =- 12604 THEN
            exp_f := 4;
        ELSIF x =- 12603 THEN
            exp_f := 4;
        ELSIF x =- 12602 THEN
            exp_f := 4;
        ELSIF x =- 12601 THEN
            exp_f := 4;
        ELSIF x =- 12600 THEN
            exp_f := 4;
        ELSIF x =- 12599 THEN
            exp_f := 4;
        ELSIF x =- 12598 THEN
            exp_f := 4;
        ELSIF x =- 12597 THEN
            exp_f := 4;
        ELSIF x =- 12596 THEN
            exp_f := 4;
        ELSIF x =- 12595 THEN
            exp_f := 4;
        ELSIF x =- 12594 THEN
            exp_f := 4;
        ELSIF x =- 12593 THEN
            exp_f := 4;
        ELSIF x =- 12592 THEN
            exp_f := 4;
        ELSIF x =- 12591 THEN
            exp_f := 4;
        ELSIF x =- 12590 THEN
            exp_f := 4;
        ELSIF x =- 12589 THEN
            exp_f := 4;
        ELSIF x =- 12588 THEN
            exp_f := 4;
        ELSIF x =- 12587 THEN
            exp_f := 4;
        ELSIF x =- 12586 THEN
            exp_f := 4;
        ELSIF x =- 12585 THEN
            exp_f := 4;
        ELSIF x =- 12584 THEN
            exp_f := 4;
        ELSIF x =- 12583 THEN
            exp_f := 4;
        ELSIF x =- 12582 THEN
            exp_f := 4;
        ELSIF x =- 12581 THEN
            exp_f := 4;
        ELSIF x =- 12580 THEN
            exp_f := 4;
        ELSIF x =- 12579 THEN
            exp_f := 4;
        ELSIF x =- 12578 THEN
            exp_f := 4;
        ELSIF x =- 12577 THEN
            exp_f := 4;
        ELSIF x =- 12576 THEN
            exp_f := 4;
        ELSIF x =- 12575 THEN
            exp_f := 4;
        ELSIF x =- 12574 THEN
            exp_f := 4;
        ELSIF x =- 12573 THEN
            exp_f := 4;
        ELSIF x =- 12572 THEN
            exp_f := 4;
        ELSIF x =- 12571 THEN
            exp_f := 4;
        ELSIF x =- 12570 THEN
            exp_f := 4;
        ELSIF x =- 12569 THEN
            exp_f := 4;
        ELSIF x =- 12568 THEN
            exp_f := 4;
        ELSIF x =- 12567 THEN
            exp_f := 4;
        ELSIF x =- 12566 THEN
            exp_f := 4;
        ELSIF x =- 12565 THEN
            exp_f := 4;
        ELSIF x =- 12564 THEN
            exp_f := 4;
        ELSIF x =- 12563 THEN
            exp_f := 4;
        ELSIF x =- 12562 THEN
            exp_f := 4;
        ELSIF x =- 12561 THEN
            exp_f := 4;
        ELSIF x =- 12560 THEN
            exp_f := 4;
        ELSIF x =- 12559 THEN
            exp_f := 4;
        ELSIF x =- 12558 THEN
            exp_f := 4;
        ELSIF x =- 12557 THEN
            exp_f := 4;
        ELSIF x =- 12556 THEN
            exp_f := 4;
        ELSIF x =- 12555 THEN
            exp_f := 4;
        ELSIF x =- 12554 THEN
            exp_f := 4;
        ELSIF x =- 12553 THEN
            exp_f := 4;
        ELSIF x =- 12552 THEN
            exp_f := 4;
        ELSIF x =- 12551 THEN
            exp_f := 4;
        ELSIF x =- 12550 THEN
            exp_f := 4;
        ELSIF x =- 12549 THEN
            exp_f := 4;
        ELSIF x =- 12548 THEN
            exp_f := 4;
        ELSIF x =- 12547 THEN
            exp_f := 4;
        ELSIF x =- 12546 THEN
            exp_f := 4;
        ELSIF x =- 12545 THEN
            exp_f := 4;
        ELSIF x =- 12544 THEN
            exp_f := 4;
        ELSIF x =- 12543 THEN
            exp_f := 4;
        ELSIF x =- 12542 THEN
            exp_f := 4;
        ELSIF x =- 12541 THEN
            exp_f := 4;
        ELSIF x =- 12540 THEN
            exp_f := 4;
        ELSIF x =- 12539 THEN
            exp_f := 4;
        ELSIF x =- 12538 THEN
            exp_f := 4;
        ELSIF x =- 12537 THEN
            exp_f := 4;
        ELSIF x =- 12536 THEN
            exp_f := 4;
        ELSIF x =- 12535 THEN
            exp_f := 4;
        ELSIF x =- 12534 THEN
            exp_f := 4;
        ELSIF x =- 12533 THEN
            exp_f := 4;
        ELSIF x =- 12532 THEN
            exp_f := 4;
        ELSIF x =- 12531 THEN
            exp_f := 4;
        ELSIF x =- 12530 THEN
            exp_f := 4;
        ELSIF x =- 12529 THEN
            exp_f := 4;
        ELSIF x =- 12528 THEN
            exp_f := 4;
        ELSIF x =- 12527 THEN
            exp_f := 4;
        ELSIF x =- 12526 THEN
            exp_f := 4;
        ELSIF x =- 12525 THEN
            exp_f := 4;
        ELSIF x =- 12524 THEN
            exp_f := 4;
        ELSIF x =- 12523 THEN
            exp_f := 4;
        ELSIF x =- 12522 THEN
            exp_f := 4;
        ELSIF x =- 12521 THEN
            exp_f := 4;
        ELSIF x =- 12520 THEN
            exp_f := 4;
        ELSIF x =- 12519 THEN
            exp_f := 4;
        ELSIF x =- 12518 THEN
            exp_f := 4;
        ELSIF x =- 12517 THEN
            exp_f := 4;
        ELSIF x =- 12516 THEN
            exp_f := 4;
        ELSIF x =- 12515 THEN
            exp_f := 4;
        ELSIF x =- 12514 THEN
            exp_f := 4;
        ELSIF x =- 12513 THEN
            exp_f := 4;
        ELSIF x =- 12512 THEN
            exp_f := 4;
        ELSIF x =- 12511 THEN
            exp_f := 4;
        ELSIF x =- 12510 THEN
            exp_f := 4;
        ELSIF x =- 12509 THEN
            exp_f := 4;
        ELSIF x =- 12508 THEN
            exp_f := 4;
        ELSIF x =- 12507 THEN
            exp_f := 4;
        ELSIF x =- 12506 THEN
            exp_f := 4;
        ELSIF x =- 12505 THEN
            exp_f := 4;
        ELSIF x =- 12504 THEN
            exp_f := 4;
        ELSIF x =- 12503 THEN
            exp_f := 4;
        ELSIF x =- 12502 THEN
            exp_f := 4;
        ELSIF x =- 12501 THEN
            exp_f := 4;
        ELSIF x =- 12500 THEN
            exp_f := 4;
        ELSIF x =- 12499 THEN
            exp_f := 4;
        ELSIF x =- 12498 THEN
            exp_f := 4;
        ELSIF x =- 12497 THEN
            exp_f := 4;
        ELSIF x =- 12496 THEN
            exp_f := 4;
        ELSIF x =- 12495 THEN
            exp_f := 4;
        ELSIF x =- 12494 THEN
            exp_f := 4;
        ELSIF x =- 12493 THEN
            exp_f := 4;
        ELSIF x =- 12492 THEN
            exp_f := 4;
        ELSIF x =- 12491 THEN
            exp_f := 4;
        ELSIF x =- 12490 THEN
            exp_f := 4;
        ELSIF x =- 12489 THEN
            exp_f := 4;
        ELSIF x =- 12488 THEN
            exp_f := 4;
        ELSIF x =- 12487 THEN
            exp_f := 4;
        ELSIF x =- 12486 THEN
            exp_f := 4;
        ELSIF x =- 12485 THEN
            exp_f := 4;
        ELSIF x =- 12484 THEN
            exp_f := 4;
        ELSIF x =- 12483 THEN
            exp_f := 4;
        ELSIF x =- 12482 THEN
            exp_f := 4;
        ELSIF x =- 12481 THEN
            exp_f := 4;
        ELSIF x =- 12480 THEN
            exp_f := 4;
        ELSIF x =- 12479 THEN
            exp_f := 4;
        ELSIF x =- 12478 THEN
            exp_f := 4;
        ELSIF x =- 12477 THEN
            exp_f := 4;
        ELSIF x =- 12476 THEN
            exp_f := 4;
        ELSIF x =- 12475 THEN
            exp_f := 4;
        ELSIF x =- 12474 THEN
            exp_f := 4;
        ELSIF x =- 12473 THEN
            exp_f := 4;
        ELSIF x =- 12472 THEN
            exp_f := 4;
        ELSIF x =- 12471 THEN
            exp_f := 4;
        ELSIF x =- 12470 THEN
            exp_f := 4;
        ELSIF x =- 12469 THEN
            exp_f := 4;
        ELSIF x =- 12468 THEN
            exp_f := 4;
        ELSIF x =- 12467 THEN
            exp_f := 4;
        ELSIF x =- 12466 THEN
            exp_f := 4;
        ELSIF x =- 12465 THEN
            exp_f := 4;
        ELSIF x =- 12464 THEN
            exp_f := 4;
        ELSIF x =- 12463 THEN
            exp_f := 4;
        ELSIF x =- 12462 THEN
            exp_f := 4;
        ELSIF x =- 12461 THEN
            exp_f := 4;
        ELSIF x =- 12460 THEN
            exp_f := 4;
        ELSIF x =- 12459 THEN
            exp_f := 4;
        ELSIF x =- 12458 THEN
            exp_f := 4;
        ELSIF x =- 12457 THEN
            exp_f := 4;
        ELSIF x =- 12456 THEN
            exp_f := 4;
        ELSIF x =- 12455 THEN
            exp_f := 4;
        ELSIF x =- 12454 THEN
            exp_f := 4;
        ELSIF x =- 12453 THEN
            exp_f := 4;
        ELSIF x =- 12452 THEN
            exp_f := 4;
        ELSIF x =- 12451 THEN
            exp_f := 4;
        ELSIF x =- 12450 THEN
            exp_f := 4;
        ELSIF x =- 12449 THEN
            exp_f := 4;
        ELSIF x =- 12448 THEN
            exp_f := 4;
        ELSIF x =- 12447 THEN
            exp_f := 4;
        ELSIF x =- 12446 THEN
            exp_f := 4;
        ELSIF x =- 12445 THEN
            exp_f := 4;
        ELSIF x =- 12444 THEN
            exp_f := 4;
        ELSIF x =- 12443 THEN
            exp_f := 4;
        ELSIF x =- 12442 THEN
            exp_f := 4;
        ELSIF x =- 12441 THEN
            exp_f := 4;
        ELSIF x =- 12440 THEN
            exp_f := 4;
        ELSIF x =- 12439 THEN
            exp_f := 4;
        ELSIF x =- 12438 THEN
            exp_f := 4;
        ELSIF x =- 12437 THEN
            exp_f := 4;
        ELSIF x =- 12436 THEN
            exp_f := 4;
        ELSIF x =- 12435 THEN
            exp_f := 4;
        ELSIF x =- 12434 THEN
            exp_f := 4;
        ELSIF x =- 12433 THEN
            exp_f := 4;
        ELSIF x =- 12432 THEN
            exp_f := 4;
        ELSIF x =- 12431 THEN
            exp_f := 4;
        ELSIF x =- 12430 THEN
            exp_f := 4;
        ELSIF x =- 12429 THEN
            exp_f := 4;
        ELSIF x =- 12428 THEN
            exp_f := 4;
        ELSIF x =- 12427 THEN
            exp_f := 4;
        ELSIF x =- 12426 THEN
            exp_f := 4;
        ELSIF x =- 12425 THEN
            exp_f := 4;
        ELSIF x =- 12424 THEN
            exp_f := 4;
        ELSIF x =- 12423 THEN
            exp_f := 4;
        ELSIF x =- 12422 THEN
            exp_f := 4;
        ELSIF x =- 12421 THEN
            exp_f := 4;
        ELSIF x =- 12420 THEN
            exp_f := 4;
        ELSIF x =- 12419 THEN
            exp_f := 4;
        ELSIF x =- 12418 THEN
            exp_f := 4;
        ELSIF x =- 12417 THEN
            exp_f := 4;
        ELSIF x =- 12416 THEN
            exp_f := 4;
        ELSIF x =- 12415 THEN
            exp_f := 4;
        ELSIF x =- 12414 THEN
            exp_f := 4;
        ELSIF x =- 12413 THEN
            exp_f := 4;
        ELSIF x =- 12412 THEN
            exp_f := 4;
        ELSIF x =- 12411 THEN
            exp_f := 4;
        ELSIF x =- 12410 THEN
            exp_f := 4;
        ELSIF x =- 12409 THEN
            exp_f := 4;
        ELSIF x =- 12408 THEN
            exp_f := 4;
        ELSIF x =- 12407 THEN
            exp_f := 4;
        ELSIF x =- 12406 THEN
            exp_f := 4;
        ELSIF x =- 12405 THEN
            exp_f := 4;
        ELSIF x =- 12404 THEN
            exp_f := 4;
        ELSIF x =- 12403 THEN
            exp_f := 4;
        ELSIF x =- 12402 THEN
            exp_f := 4;
        ELSIF x =- 12401 THEN
            exp_f := 4;
        ELSIF x =- 12400 THEN
            exp_f := 4;
        ELSIF x =- 12399 THEN
            exp_f := 4;
        ELSIF x =- 12398 THEN
            exp_f := 4;
        ELSIF x =- 12397 THEN
            exp_f := 4;
        ELSIF x =- 12396 THEN
            exp_f := 4;
        ELSIF x =- 12395 THEN
            exp_f := 4;
        ELSIF x =- 12394 THEN
            exp_f := 4;
        ELSIF x =- 12393 THEN
            exp_f := 4;
        ELSIF x =- 12392 THEN
            exp_f := 4;
        ELSIF x =- 12391 THEN
            exp_f := 4;
        ELSIF x =- 12390 THEN
            exp_f := 4;
        ELSIF x =- 12389 THEN
            exp_f := 4;
        ELSIF x =- 12388 THEN
            exp_f := 4;
        ELSIF x =- 12387 THEN
            exp_f := 4;
        ELSIF x =- 12386 THEN
            exp_f := 4;
        ELSIF x =- 12385 THEN
            exp_f := 4;
        ELSIF x =- 12384 THEN
            exp_f := 4;
        ELSIF x =- 12383 THEN
            exp_f := 4;
        ELSIF x =- 12382 THEN
            exp_f := 4;
        ELSIF x =- 12381 THEN
            exp_f := 4;
        ELSIF x =- 12380 THEN
            exp_f := 4;
        ELSIF x =- 12379 THEN
            exp_f := 4;
        ELSIF x =- 12378 THEN
            exp_f := 4;
        ELSIF x =- 12377 THEN
            exp_f := 4;
        ELSIF x =- 12376 THEN
            exp_f := 4;
        ELSIF x =- 12375 THEN
            exp_f := 4;
        ELSIF x =- 12374 THEN
            exp_f := 4;
        ELSIF x =- 12373 THEN
            exp_f := 4;
        ELSIF x =- 12372 THEN
            exp_f := 4;
        ELSIF x =- 12371 THEN
            exp_f := 4;
        ELSIF x =- 12370 THEN
            exp_f := 4;
        ELSIF x =- 12369 THEN
            exp_f := 4;
        ELSIF x =- 12368 THEN
            exp_f := 4;
        ELSIF x =- 12367 THEN
            exp_f := 4;
        ELSIF x =- 12366 THEN
            exp_f := 4;
        ELSIF x =- 12365 THEN
            exp_f := 4;
        ELSIF x =- 12364 THEN
            exp_f := 4;
        ELSIF x =- 12363 THEN
            exp_f := 4;
        ELSIF x =- 12362 THEN
            exp_f := 4;
        ELSIF x =- 12361 THEN
            exp_f := 4;
        ELSIF x =- 12360 THEN
            exp_f := 4;
        ELSIF x =- 12359 THEN
            exp_f := 4;
        ELSIF x =- 12358 THEN
            exp_f := 4;
        ELSIF x =- 12357 THEN
            exp_f := 4;
        ELSIF x =- 12356 THEN
            exp_f := 4;
        ELSIF x =- 12355 THEN
            exp_f := 4;
        ELSIF x =- 12354 THEN
            exp_f := 4;
        ELSIF x =- 12353 THEN
            exp_f := 4;
        ELSIF x =- 12352 THEN
            exp_f := 4;
        ELSIF x =- 12351 THEN
            exp_f := 4;
        ELSIF x =- 12350 THEN
            exp_f := 4;
        ELSIF x =- 12349 THEN
            exp_f := 4;
        ELSIF x =- 12348 THEN
            exp_f := 4;
        ELSIF x =- 12347 THEN
            exp_f := 4;
        ELSIF x =- 12346 THEN
            exp_f := 4;
        ELSIF x =- 12345 THEN
            exp_f := 4;
        ELSIF x =- 12344 THEN
            exp_f := 4;
        ELSIF x =- 12343 THEN
            exp_f := 4;
        ELSIF x =- 12342 THEN
            exp_f := 4;
        ELSIF x =- 12341 THEN
            exp_f := 4;
        ELSIF x =- 12340 THEN
            exp_f := 4;
        ELSIF x =- 12339 THEN
            exp_f := 4;
        ELSIF x =- 12338 THEN
            exp_f := 4;
        ELSIF x =- 12337 THEN
            exp_f := 4;
        ELSIF x =- 12336 THEN
            exp_f := 4;
        ELSIF x =- 12335 THEN
            exp_f := 4;
        ELSIF x =- 12334 THEN
            exp_f := 4;
        ELSIF x =- 12333 THEN
            exp_f := 4;
        ELSIF x =- 12332 THEN
            exp_f := 4;
        ELSIF x =- 12331 THEN
            exp_f := 4;
        ELSIF x =- 12330 THEN
            exp_f := 4;
        ELSIF x =- 12329 THEN
            exp_f := 4;
        ELSIF x =- 12328 THEN
            exp_f := 4;
        ELSIF x =- 12327 THEN
            exp_f := 4;
        ELSIF x =- 12326 THEN
            exp_f := 4;
        ELSIF x =- 12325 THEN
            exp_f := 4;
        ELSIF x =- 12324 THEN
            exp_f := 4;
        ELSIF x =- 12323 THEN
            exp_f := 4;
        ELSIF x =- 12322 THEN
            exp_f := 4;
        ELSIF x =- 12321 THEN
            exp_f := 4;
        ELSIF x =- 12320 THEN
            exp_f := 4;
        ELSIF x =- 12319 THEN
            exp_f := 4;
        ELSIF x =- 12318 THEN
            exp_f := 4;
        ELSIF x =- 12317 THEN
            exp_f := 4;
        ELSIF x =- 12316 THEN
            exp_f := 4;
        ELSIF x =- 12315 THEN
            exp_f := 4;
        ELSIF x =- 12314 THEN
            exp_f := 4;
        ELSIF x =- 12313 THEN
            exp_f := 4;
        ELSIF x =- 12312 THEN
            exp_f := 4;
        ELSIF x =- 12311 THEN
            exp_f := 4;
        ELSIF x =- 12310 THEN
            exp_f := 4;
        ELSIF x =- 12309 THEN
            exp_f := 4;
        ELSIF x =- 12308 THEN
            exp_f := 4;
        ELSIF x =- 12307 THEN
            exp_f := 4;
        ELSIF x =- 12306 THEN
            exp_f := 4;
        ELSIF x =- 12305 THEN
            exp_f := 4;
        ELSIF x =- 12304 THEN
            exp_f := 4;
        ELSIF x =- 12303 THEN
            exp_f := 4;
        ELSIF x =- 12302 THEN
            exp_f := 4;
        ELSIF x =- 12301 THEN
            exp_f := 4;
        ELSIF x =- 12300 THEN
            exp_f := 4;
        ELSIF x =- 12299 THEN
            exp_f := 4;
        ELSIF x =- 12298 THEN
            exp_f := 4;
        ELSIF x =- 12297 THEN
            exp_f := 4;
        ELSIF x =- 12296 THEN
            exp_f := 4;
        ELSIF x =- 12295 THEN
            exp_f := 4;
        ELSIF x =- 12294 THEN
            exp_f := 4;
        ELSIF x =- 12293 THEN
            exp_f := 4;
        ELSIF x =- 12292 THEN
            exp_f := 4;
        ELSIF x =- 12291 THEN
            exp_f := 4;
        ELSIF x =- 12290 THEN
            exp_f := 4;
        ELSIF x =- 12289 THEN
            exp_f := 4;
        ELSIF x =- 12288 THEN
            exp_f := 4;
        ELSIF x =- 12287 THEN
            exp_f := 6;
        ELSIF x =- 12286 THEN
            exp_f := 6;
        ELSIF x =- 12285 THEN
            exp_f := 6;
        ELSIF x =- 12284 THEN
            exp_f := 6;
        ELSIF x =- 12283 THEN
            exp_f := 6;
        ELSIF x =- 12282 THEN
            exp_f := 6;
        ELSIF x =- 12281 THEN
            exp_f := 6;
        ELSIF x =- 12280 THEN
            exp_f := 6;
        ELSIF x =- 12279 THEN
            exp_f := 6;
        ELSIF x =- 12278 THEN
            exp_f := 6;
        ELSIF x =- 12277 THEN
            exp_f := 6;
        ELSIF x =- 12276 THEN
            exp_f := 6;
        ELSIF x =- 12275 THEN
            exp_f := 6;
        ELSIF x =- 12274 THEN
            exp_f := 6;
        ELSIF x =- 12273 THEN
            exp_f := 6;
        ELSIF x =- 12272 THEN
            exp_f := 6;
        ELSIF x =- 12271 THEN
            exp_f := 6;
        ELSIF x =- 12270 THEN
            exp_f := 6;
        ELSIF x =- 12269 THEN
            exp_f := 6;
        ELSIF x =- 12268 THEN
            exp_f := 6;
        ELSIF x =- 12267 THEN
            exp_f := 6;
        ELSIF x =- 12266 THEN
            exp_f := 6;
        ELSIF x =- 12265 THEN
            exp_f := 6;
        ELSIF x =- 12264 THEN
            exp_f := 6;
        ELSIF x =- 12263 THEN
            exp_f := 6;
        ELSIF x =- 12262 THEN
            exp_f := 6;
        ELSIF x =- 12261 THEN
            exp_f := 6;
        ELSIF x =- 12260 THEN
            exp_f := 6;
        ELSIF x =- 12259 THEN
            exp_f := 6;
        ELSIF x =- 12258 THEN
            exp_f := 6;
        ELSIF x =- 12257 THEN
            exp_f := 6;
        ELSIF x =- 12256 THEN
            exp_f := 6;
        ELSIF x =- 12255 THEN
            exp_f := 6;
        ELSIF x =- 12254 THEN
            exp_f := 6;
        ELSIF x =- 12253 THEN
            exp_f := 6;
        ELSIF x =- 12252 THEN
            exp_f := 6;
        ELSIF x =- 12251 THEN
            exp_f := 6;
        ELSIF x =- 12250 THEN
            exp_f := 6;
        ELSIF x =- 12249 THEN
            exp_f := 6;
        ELSIF x =- 12248 THEN
            exp_f := 6;
        ELSIF x =- 12247 THEN
            exp_f := 6;
        ELSIF x =- 12246 THEN
            exp_f := 6;
        ELSIF x =- 12245 THEN
            exp_f := 6;
        ELSIF x =- 12244 THEN
            exp_f := 6;
        ELSIF x =- 12243 THEN
            exp_f := 6;
        ELSIF x =- 12242 THEN
            exp_f := 6;
        ELSIF x =- 12241 THEN
            exp_f := 6;
        ELSIF x =- 12240 THEN
            exp_f := 6;
        ELSIF x =- 12239 THEN
            exp_f := 6;
        ELSIF x =- 12238 THEN
            exp_f := 6;
        ELSIF x =- 12237 THEN
            exp_f := 6;
        ELSIF x =- 12236 THEN
            exp_f := 6;
        ELSIF x =- 12235 THEN
            exp_f := 6;
        ELSIF x =- 12234 THEN
            exp_f := 6;
        ELSIF x =- 12233 THEN
            exp_f := 6;
        ELSIF x =- 12232 THEN
            exp_f := 6;
        ELSIF x =- 12231 THEN
            exp_f := 6;
        ELSIF x =- 12230 THEN
            exp_f := 6;
        ELSIF x =- 12229 THEN
            exp_f := 6;
        ELSIF x =- 12228 THEN
            exp_f := 6;
        ELSIF x =- 12227 THEN
            exp_f := 6;
        ELSIF x =- 12226 THEN
            exp_f := 6;
        ELSIF x =- 12225 THEN
            exp_f := 6;
        ELSIF x =- 12224 THEN
            exp_f := 6;
        ELSIF x =- 12223 THEN
            exp_f := 6;
        ELSIF x =- 12222 THEN
            exp_f := 6;
        ELSIF x =- 12221 THEN
            exp_f := 6;
        ELSIF x =- 12220 THEN
            exp_f := 6;
        ELSIF x =- 12219 THEN
            exp_f := 6;
        ELSIF x =- 12218 THEN
            exp_f := 6;
        ELSIF x =- 12217 THEN
            exp_f := 6;
        ELSIF x =- 12216 THEN
            exp_f := 6;
        ELSIF x =- 12215 THEN
            exp_f := 6;
        ELSIF x =- 12214 THEN
            exp_f := 6;
        ELSIF x =- 12213 THEN
            exp_f := 6;
        ELSIF x =- 12212 THEN
            exp_f := 6;
        ELSIF x =- 12211 THEN
            exp_f := 6;
        ELSIF x =- 12210 THEN
            exp_f := 6;
        ELSIF x =- 12209 THEN
            exp_f := 6;
        ELSIF x =- 12208 THEN
            exp_f := 6;
        ELSIF x =- 12207 THEN
            exp_f := 6;
        ELSIF x =- 12206 THEN
            exp_f := 6;
        ELSIF x =- 12205 THEN
            exp_f := 6;
        ELSIF x =- 12204 THEN
            exp_f := 6;
        ELSIF x =- 12203 THEN
            exp_f := 6;
        ELSIF x =- 12202 THEN
            exp_f := 6;
        ELSIF x =- 12201 THEN
            exp_f := 6;
        ELSIF x =- 12200 THEN
            exp_f := 6;
        ELSIF x =- 12199 THEN
            exp_f := 6;
        ELSIF x =- 12198 THEN
            exp_f := 6;
        ELSIF x =- 12197 THEN
            exp_f := 6;
        ELSIF x =- 12196 THEN
            exp_f := 6;
        ELSIF x =- 12195 THEN
            exp_f := 6;
        ELSIF x =- 12194 THEN
            exp_f := 6;
        ELSIF x =- 12193 THEN
            exp_f := 6;
        ELSIF x =- 12192 THEN
            exp_f := 6;
        ELSIF x =- 12191 THEN
            exp_f := 6;
        ELSIF x =- 12190 THEN
            exp_f := 6;
        ELSIF x =- 12189 THEN
            exp_f := 6;
        ELSIF x =- 12188 THEN
            exp_f := 6;
        ELSIF x =- 12187 THEN
            exp_f := 6;
        ELSIF x =- 12186 THEN
            exp_f := 6;
        ELSIF x =- 12185 THEN
            exp_f := 6;
        ELSIF x =- 12184 THEN
            exp_f := 6;
        ELSIF x =- 12183 THEN
            exp_f := 6;
        ELSIF x =- 12182 THEN
            exp_f := 6;
        ELSIF x =- 12181 THEN
            exp_f := 6;
        ELSIF x =- 12180 THEN
            exp_f := 6;
        ELSIF x =- 12179 THEN
            exp_f := 6;
        ELSIF x =- 12178 THEN
            exp_f := 6;
        ELSIF x =- 12177 THEN
            exp_f := 6;
        ELSIF x =- 12176 THEN
            exp_f := 6;
        ELSIF x =- 12175 THEN
            exp_f := 6;
        ELSIF x =- 12174 THEN
            exp_f := 6;
        ELSIF x =- 12173 THEN
            exp_f := 6;
        ELSIF x =- 12172 THEN
            exp_f := 6;
        ELSIF x =- 12171 THEN
            exp_f := 6;
        ELSIF x =- 12170 THEN
            exp_f := 6;
        ELSIF x =- 12169 THEN
            exp_f := 6;
        ELSIF x =- 12168 THEN
            exp_f := 6;
        ELSIF x =- 12167 THEN
            exp_f := 6;
        ELSIF x =- 12166 THEN
            exp_f := 6;
        ELSIF x =- 12165 THEN
            exp_f := 6;
        ELSIF x =- 12164 THEN
            exp_f := 6;
        ELSIF x =- 12163 THEN
            exp_f := 6;
        ELSIF x =- 12162 THEN
            exp_f := 6;
        ELSIF x =- 12161 THEN
            exp_f := 6;
        ELSIF x =- 12160 THEN
            exp_f := 6;
        ELSIF x =- 12159 THEN
            exp_f := 6;
        ELSIF x =- 12158 THEN
            exp_f := 6;
        ELSIF x =- 12157 THEN
            exp_f := 6;
        ELSIF x =- 12156 THEN
            exp_f := 6;
        ELSIF x =- 12155 THEN
            exp_f := 6;
        ELSIF x =- 12154 THEN
            exp_f := 6;
        ELSIF x =- 12153 THEN
            exp_f := 6;
        ELSIF x =- 12152 THEN
            exp_f := 6;
        ELSIF x =- 12151 THEN
            exp_f := 6;
        ELSIF x =- 12150 THEN
            exp_f := 6;
        ELSIF x =- 12149 THEN
            exp_f := 6;
        ELSIF x =- 12148 THEN
            exp_f := 6;
        ELSIF x =- 12147 THEN
            exp_f := 6;
        ELSIF x =- 12146 THEN
            exp_f := 6;
        ELSIF x =- 12145 THEN
            exp_f := 6;
        ELSIF x =- 12144 THEN
            exp_f := 6;
        ELSIF x =- 12143 THEN
            exp_f := 6;
        ELSIF x =- 12142 THEN
            exp_f := 6;
        ELSIF x =- 12141 THEN
            exp_f := 6;
        ELSIF x =- 12140 THEN
            exp_f := 6;
        ELSIF x =- 12139 THEN
            exp_f := 6;
        ELSIF x =- 12138 THEN
            exp_f := 6;
        ELSIF x =- 12137 THEN
            exp_f := 6;
        ELSIF x =- 12136 THEN
            exp_f := 6;
        ELSIF x =- 12135 THEN
            exp_f := 6;
        ELSIF x =- 12134 THEN
            exp_f := 6;
        ELSIF x =- 12133 THEN
            exp_f := 6;
        ELSIF x =- 12132 THEN
            exp_f := 6;
        ELSIF x =- 12131 THEN
            exp_f := 6;
        ELSIF x =- 12130 THEN
            exp_f := 6;
        ELSIF x =- 12129 THEN
            exp_f := 6;
        ELSIF x =- 12128 THEN
            exp_f := 6;
        ELSIF x =- 12127 THEN
            exp_f := 6;
        ELSIF x =- 12126 THEN
            exp_f := 6;
        ELSIF x =- 12125 THEN
            exp_f := 6;
        ELSIF x =- 12124 THEN
            exp_f := 6;
        ELSIF x =- 12123 THEN
            exp_f := 6;
        ELSIF x =- 12122 THEN
            exp_f := 6;
        ELSIF x =- 12121 THEN
            exp_f := 6;
        ELSIF x =- 12120 THEN
            exp_f := 6;
        ELSIF x =- 12119 THEN
            exp_f := 6;
        ELSIF x =- 12118 THEN
            exp_f := 6;
        ELSIF x =- 12117 THEN
            exp_f := 6;
        ELSIF x =- 12116 THEN
            exp_f := 6;
        ELSIF x =- 12115 THEN
            exp_f := 6;
        ELSIF x =- 12114 THEN
            exp_f := 6;
        ELSIF x =- 12113 THEN
            exp_f := 6;
        ELSIF x =- 12112 THEN
            exp_f := 6;
        ELSIF x =- 12111 THEN
            exp_f := 6;
        ELSIF x =- 12110 THEN
            exp_f := 6;
        ELSIF x =- 12109 THEN
            exp_f := 6;
        ELSIF x =- 12108 THEN
            exp_f := 6;
        ELSIF x =- 12107 THEN
            exp_f := 6;
        ELSIF x =- 12106 THEN
            exp_f := 6;
        ELSIF x =- 12105 THEN
            exp_f := 6;
        ELSIF x =- 12104 THEN
            exp_f := 6;
        ELSIF x =- 12103 THEN
            exp_f := 6;
        ELSIF x =- 12102 THEN
            exp_f := 6;
        ELSIF x =- 12101 THEN
            exp_f := 6;
        ELSIF x =- 12100 THEN
            exp_f := 6;
        ELSIF x =- 12099 THEN
            exp_f := 6;
        ELSIF x =- 12098 THEN
            exp_f := 6;
        ELSIF x =- 12097 THEN
            exp_f := 6;
        ELSIF x =- 12096 THEN
            exp_f := 6;
        ELSIF x =- 12095 THEN
            exp_f := 6;
        ELSIF x =- 12094 THEN
            exp_f := 6;
        ELSIF x =- 12093 THEN
            exp_f := 6;
        ELSIF x =- 12092 THEN
            exp_f := 6;
        ELSIF x =- 12091 THEN
            exp_f := 6;
        ELSIF x =- 12090 THEN
            exp_f := 6;
        ELSIF x =- 12089 THEN
            exp_f := 6;
        ELSIF x =- 12088 THEN
            exp_f := 6;
        ELSIF x =- 12087 THEN
            exp_f := 6;
        ELSIF x =- 12086 THEN
            exp_f := 6;
        ELSIF x =- 12085 THEN
            exp_f := 6;
        ELSIF x =- 12084 THEN
            exp_f := 6;
        ELSIF x =- 12083 THEN
            exp_f := 6;
        ELSIF x =- 12082 THEN
            exp_f := 6;
        ELSIF x =- 12081 THEN
            exp_f := 6;
        ELSIF x =- 12080 THEN
            exp_f := 6;
        ELSIF x =- 12079 THEN
            exp_f := 6;
        ELSIF x =- 12078 THEN
            exp_f := 6;
        ELSIF x =- 12077 THEN
            exp_f := 6;
        ELSIF x =- 12076 THEN
            exp_f := 6;
        ELSIF x =- 12075 THEN
            exp_f := 6;
        ELSIF x =- 12074 THEN
            exp_f := 6;
        ELSIF x =- 12073 THEN
            exp_f := 6;
        ELSIF x =- 12072 THEN
            exp_f := 6;
        ELSIF x =- 12071 THEN
            exp_f := 6;
        ELSIF x =- 12070 THEN
            exp_f := 6;
        ELSIF x =- 12069 THEN
            exp_f := 6;
        ELSIF x =- 12068 THEN
            exp_f := 6;
        ELSIF x =- 12067 THEN
            exp_f := 6;
        ELSIF x =- 12066 THEN
            exp_f := 6;
        ELSIF x =- 12065 THEN
            exp_f := 6;
        ELSIF x =- 12064 THEN
            exp_f := 6;
        ELSIF x =- 12063 THEN
            exp_f := 6;
        ELSIF x =- 12062 THEN
            exp_f := 6;
        ELSIF x =- 12061 THEN
            exp_f := 6;
        ELSIF x =- 12060 THEN
            exp_f := 6;
        ELSIF x =- 12059 THEN
            exp_f := 6;
        ELSIF x =- 12058 THEN
            exp_f := 6;
        ELSIF x =- 12057 THEN
            exp_f := 6;
        ELSIF x =- 12056 THEN
            exp_f := 6;
        ELSIF x =- 12055 THEN
            exp_f := 6;
        ELSIF x =- 12054 THEN
            exp_f := 6;
        ELSIF x =- 12053 THEN
            exp_f := 6;
        ELSIF x =- 12052 THEN
            exp_f := 6;
        ELSIF x =- 12051 THEN
            exp_f := 6;
        ELSIF x =- 12050 THEN
            exp_f := 6;
        ELSIF x =- 12049 THEN
            exp_f := 6;
        ELSIF x =- 12048 THEN
            exp_f := 6;
        ELSIF x =- 12047 THEN
            exp_f := 6;
        ELSIF x =- 12046 THEN
            exp_f := 6;
        ELSIF x =- 12045 THEN
            exp_f := 6;
        ELSIF x =- 12044 THEN
            exp_f := 6;
        ELSIF x =- 12043 THEN
            exp_f := 6;
        ELSIF x =- 12042 THEN
            exp_f := 6;
        ELSIF x =- 12041 THEN
            exp_f := 6;
        ELSIF x =- 12040 THEN
            exp_f := 6;
        ELSIF x =- 12039 THEN
            exp_f := 6;
        ELSIF x =- 12038 THEN
            exp_f := 6;
        ELSIF x =- 12037 THEN
            exp_f := 6;
        ELSIF x =- 12036 THEN
            exp_f := 6;
        ELSIF x =- 12035 THEN
            exp_f := 6;
        ELSIF x =- 12034 THEN
            exp_f := 6;
        ELSIF x =- 12033 THEN
            exp_f := 6;
        ELSIF x =- 12032 THEN
            exp_f := 6;
        ELSIF x =- 12031 THEN
            exp_f := 6;
        ELSIF x =- 12030 THEN
            exp_f := 6;
        ELSIF x =- 12029 THEN
            exp_f := 6;
        ELSIF x =- 12028 THEN
            exp_f := 6;
        ELSIF x =- 12027 THEN
            exp_f := 6;
        ELSIF x =- 12026 THEN
            exp_f := 6;
        ELSIF x =- 12025 THEN
            exp_f := 6;
        ELSIF x =- 12024 THEN
            exp_f := 6;
        ELSIF x =- 12023 THEN
            exp_f := 6;
        ELSIF x =- 12022 THEN
            exp_f := 6;
        ELSIF x =- 12021 THEN
            exp_f := 6;
        ELSIF x =- 12020 THEN
            exp_f := 6;
        ELSIF x =- 12019 THEN
            exp_f := 6;
        ELSIF x =- 12018 THEN
            exp_f := 6;
        ELSIF x =- 12017 THEN
            exp_f := 6;
        ELSIF x =- 12016 THEN
            exp_f := 6;
        ELSIF x =- 12015 THEN
            exp_f := 6;
        ELSIF x =- 12014 THEN
            exp_f := 6;
        ELSIF x =- 12013 THEN
            exp_f := 6;
        ELSIF x =- 12012 THEN
            exp_f := 6;
        ELSIF x =- 12011 THEN
            exp_f := 6;
        ELSIF x =- 12010 THEN
            exp_f := 6;
        ELSIF x =- 12009 THEN
            exp_f := 6;
        ELSIF x =- 12008 THEN
            exp_f := 6;
        ELSIF x =- 12007 THEN
            exp_f := 6;
        ELSIF x =- 12006 THEN
            exp_f := 6;
        ELSIF x =- 12005 THEN
            exp_f := 6;
        ELSIF x =- 12004 THEN
            exp_f := 6;
        ELSIF x =- 12003 THEN
            exp_f := 6;
        ELSIF x =- 12002 THEN
            exp_f := 6;
        ELSIF x =- 12001 THEN
            exp_f := 6;
        ELSIF x =- 12000 THEN
            exp_f := 6;
        ELSIF x =- 11999 THEN
            exp_f := 6;
        ELSIF x =- 11998 THEN
            exp_f := 6;
        ELSIF x =- 11997 THEN
            exp_f := 6;
        ELSIF x =- 11996 THEN
            exp_f := 6;
        ELSIF x =- 11995 THEN
            exp_f := 6;
        ELSIF x =- 11994 THEN
            exp_f := 6;
        ELSIF x =- 11993 THEN
            exp_f := 6;
        ELSIF x =- 11992 THEN
            exp_f := 6;
        ELSIF x =- 11991 THEN
            exp_f := 6;
        ELSIF x =- 11990 THEN
            exp_f := 6;
        ELSIF x =- 11989 THEN
            exp_f := 6;
        ELSIF x =- 11988 THEN
            exp_f := 6;
        ELSIF x =- 11987 THEN
            exp_f := 6;
        ELSIF x =- 11986 THEN
            exp_f := 6;
        ELSIF x =- 11985 THEN
            exp_f := 6;
        ELSIF x =- 11984 THEN
            exp_f := 6;
        ELSIF x =- 11983 THEN
            exp_f := 6;
        ELSIF x =- 11982 THEN
            exp_f := 6;
        ELSIF x =- 11981 THEN
            exp_f := 6;
        ELSIF x =- 11980 THEN
            exp_f := 6;
        ELSIF x =- 11979 THEN
            exp_f := 6;
        ELSIF x =- 11978 THEN
            exp_f := 6;
        ELSIF x =- 11977 THEN
            exp_f := 6;
        ELSIF x =- 11976 THEN
            exp_f := 6;
        ELSIF x =- 11975 THEN
            exp_f := 6;
        ELSIF x =- 11974 THEN
            exp_f := 6;
        ELSIF x =- 11973 THEN
            exp_f := 6;
        ELSIF x =- 11972 THEN
            exp_f := 6;
        ELSIF x =- 11971 THEN
            exp_f := 6;
        ELSIF x =- 11970 THEN
            exp_f := 6;
        ELSIF x =- 11969 THEN
            exp_f := 6;
        ELSIF x =- 11968 THEN
            exp_f := 6;
        ELSIF x =- 11967 THEN
            exp_f := 6;
        ELSIF x =- 11966 THEN
            exp_f := 6;
        ELSIF x =- 11965 THEN
            exp_f := 6;
        ELSIF x =- 11964 THEN
            exp_f := 6;
        ELSIF x =- 11963 THEN
            exp_f := 6;
        ELSIF x =- 11962 THEN
            exp_f := 6;
        ELSIF x =- 11961 THEN
            exp_f := 6;
        ELSIF x =- 11960 THEN
            exp_f := 6;
        ELSIF x =- 11959 THEN
            exp_f := 6;
        ELSIF x =- 11958 THEN
            exp_f := 6;
        ELSIF x =- 11957 THEN
            exp_f := 6;
        ELSIF x =- 11956 THEN
            exp_f := 6;
        ELSIF x =- 11955 THEN
            exp_f := 6;
        ELSIF x =- 11954 THEN
            exp_f := 6;
        ELSIF x =- 11953 THEN
            exp_f := 6;
        ELSIF x =- 11952 THEN
            exp_f := 6;
        ELSIF x =- 11951 THEN
            exp_f := 6;
        ELSIF x =- 11950 THEN
            exp_f := 6;
        ELSIF x =- 11949 THEN
            exp_f := 6;
        ELSIF x =- 11948 THEN
            exp_f := 6;
        ELSIF x =- 11947 THEN
            exp_f := 6;
        ELSIF x =- 11946 THEN
            exp_f := 6;
        ELSIF x =- 11945 THEN
            exp_f := 6;
        ELSIF x =- 11944 THEN
            exp_f := 6;
        ELSIF x =- 11943 THEN
            exp_f := 6;
        ELSIF x =- 11942 THEN
            exp_f := 6;
        ELSIF x =- 11941 THEN
            exp_f := 6;
        ELSIF x =- 11940 THEN
            exp_f := 6;
        ELSIF x =- 11939 THEN
            exp_f := 6;
        ELSIF x =- 11938 THEN
            exp_f := 6;
        ELSIF x =- 11937 THEN
            exp_f := 6;
        ELSIF x =- 11936 THEN
            exp_f := 6;
        ELSIF x =- 11935 THEN
            exp_f := 6;
        ELSIF x =- 11934 THEN
            exp_f := 6;
        ELSIF x =- 11933 THEN
            exp_f := 6;
        ELSIF x =- 11932 THEN
            exp_f := 6;
        ELSIF x =- 11931 THEN
            exp_f := 6;
        ELSIF x =- 11930 THEN
            exp_f := 6;
        ELSIF x =- 11929 THEN
            exp_f := 6;
        ELSIF x =- 11928 THEN
            exp_f := 6;
        ELSIF x =- 11927 THEN
            exp_f := 6;
        ELSIF x =- 11926 THEN
            exp_f := 6;
        ELSIF x =- 11925 THEN
            exp_f := 6;
        ELSIF x =- 11924 THEN
            exp_f := 6;
        ELSIF x =- 11923 THEN
            exp_f := 6;
        ELSIF x =- 11922 THEN
            exp_f := 6;
        ELSIF x =- 11921 THEN
            exp_f := 6;
        ELSIF x =- 11920 THEN
            exp_f := 6;
        ELSIF x =- 11919 THEN
            exp_f := 6;
        ELSIF x =- 11918 THEN
            exp_f := 6;
        ELSIF x =- 11917 THEN
            exp_f := 6;
        ELSIF x =- 11916 THEN
            exp_f := 6;
        ELSIF x =- 11915 THEN
            exp_f := 6;
        ELSIF x =- 11914 THEN
            exp_f := 6;
        ELSIF x =- 11913 THEN
            exp_f := 6;
        ELSIF x =- 11912 THEN
            exp_f := 6;
        ELSIF x =- 11911 THEN
            exp_f := 6;
        ELSIF x =- 11910 THEN
            exp_f := 6;
        ELSIF x =- 11909 THEN
            exp_f := 6;
        ELSIF x =- 11908 THEN
            exp_f := 6;
        ELSIF x =- 11907 THEN
            exp_f := 6;
        ELSIF x =- 11906 THEN
            exp_f := 6;
        ELSIF x =- 11905 THEN
            exp_f := 6;
        ELSIF x =- 11904 THEN
            exp_f := 6;
        ELSIF x =- 11903 THEN
            exp_f := 6;
        ELSIF x =- 11902 THEN
            exp_f := 6;
        ELSIF x =- 11901 THEN
            exp_f := 6;
        ELSIF x =- 11900 THEN
            exp_f := 6;
        ELSIF x =- 11899 THEN
            exp_f := 6;
        ELSIF x =- 11898 THEN
            exp_f := 6;
        ELSIF x =- 11897 THEN
            exp_f := 6;
        ELSIF x =- 11896 THEN
            exp_f := 6;
        ELSIF x =- 11895 THEN
            exp_f := 6;
        ELSIF x =- 11894 THEN
            exp_f := 6;
        ELSIF x =- 11893 THEN
            exp_f := 6;
        ELSIF x =- 11892 THEN
            exp_f := 6;
        ELSIF x =- 11891 THEN
            exp_f := 6;
        ELSIF x =- 11890 THEN
            exp_f := 6;
        ELSIF x =- 11889 THEN
            exp_f := 6;
        ELSIF x =- 11888 THEN
            exp_f := 6;
        ELSIF x =- 11887 THEN
            exp_f := 6;
        ELSIF x =- 11886 THEN
            exp_f := 6;
        ELSIF x =- 11885 THEN
            exp_f := 6;
        ELSIF x =- 11884 THEN
            exp_f := 6;
        ELSIF x =- 11883 THEN
            exp_f := 6;
        ELSIF x =- 11882 THEN
            exp_f := 6;
        ELSIF x =- 11881 THEN
            exp_f := 6;
        ELSIF x =- 11880 THEN
            exp_f := 6;
        ELSIF x =- 11879 THEN
            exp_f := 6;
        ELSIF x =- 11878 THEN
            exp_f := 6;
        ELSIF x =- 11877 THEN
            exp_f := 6;
        ELSIF x =- 11876 THEN
            exp_f := 6;
        ELSIF x =- 11875 THEN
            exp_f := 6;
        ELSIF x =- 11874 THEN
            exp_f := 6;
        ELSIF x =- 11873 THEN
            exp_f := 6;
        ELSIF x =- 11872 THEN
            exp_f := 6;
        ELSIF x =- 11871 THEN
            exp_f := 6;
        ELSIF x =- 11870 THEN
            exp_f := 6;
        ELSIF x =- 11869 THEN
            exp_f := 6;
        ELSIF x =- 11868 THEN
            exp_f := 6;
        ELSIF x =- 11867 THEN
            exp_f := 6;
        ELSIF x =- 11866 THEN
            exp_f := 6;
        ELSIF x =- 11865 THEN
            exp_f := 6;
        ELSIF x =- 11864 THEN
            exp_f := 6;
        ELSIF x =- 11863 THEN
            exp_f := 6;
        ELSIF x =- 11862 THEN
            exp_f := 6;
        ELSIF x =- 11861 THEN
            exp_f := 6;
        ELSIF x =- 11860 THEN
            exp_f := 6;
        ELSIF x =- 11859 THEN
            exp_f := 6;
        ELSIF x =- 11858 THEN
            exp_f := 6;
        ELSIF x =- 11857 THEN
            exp_f := 6;
        ELSIF x =- 11856 THEN
            exp_f := 6;
        ELSIF x =- 11855 THEN
            exp_f := 6;
        ELSIF x =- 11854 THEN
            exp_f := 6;
        ELSIF x =- 11853 THEN
            exp_f := 6;
        ELSIF x =- 11852 THEN
            exp_f := 6;
        ELSIF x =- 11851 THEN
            exp_f := 6;
        ELSIF x =- 11850 THEN
            exp_f := 6;
        ELSIF x =- 11849 THEN
            exp_f := 6;
        ELSIF x =- 11848 THEN
            exp_f := 6;
        ELSIF x =- 11847 THEN
            exp_f := 6;
        ELSIF x =- 11846 THEN
            exp_f := 6;
        ELSIF x =- 11845 THEN
            exp_f := 6;
        ELSIF x =- 11844 THEN
            exp_f := 6;
        ELSIF x =- 11843 THEN
            exp_f := 6;
        ELSIF x =- 11842 THEN
            exp_f := 6;
        ELSIF x =- 11841 THEN
            exp_f := 6;
        ELSIF x =- 11840 THEN
            exp_f := 6;
        ELSIF x =- 11839 THEN
            exp_f := 6;
        ELSIF x =- 11838 THEN
            exp_f := 6;
        ELSIF x =- 11837 THEN
            exp_f := 6;
        ELSIF x =- 11836 THEN
            exp_f := 6;
        ELSIF x =- 11835 THEN
            exp_f := 6;
        ELSIF x =- 11834 THEN
            exp_f := 6;
        ELSIF x =- 11833 THEN
            exp_f := 6;
        ELSIF x =- 11832 THEN
            exp_f := 6;
        ELSIF x =- 11831 THEN
            exp_f := 6;
        ELSIF x =- 11830 THEN
            exp_f := 6;
        ELSIF x =- 11829 THEN
            exp_f := 6;
        ELSIF x =- 11828 THEN
            exp_f := 6;
        ELSIF x =- 11827 THEN
            exp_f := 6;
        ELSIF x =- 11826 THEN
            exp_f := 6;
        ELSIF x =- 11825 THEN
            exp_f := 6;
        ELSIF x =- 11824 THEN
            exp_f := 6;
        ELSIF x =- 11823 THEN
            exp_f := 6;
        ELSIF x =- 11822 THEN
            exp_f := 6;
        ELSIF x =- 11821 THEN
            exp_f := 6;
        ELSIF x =- 11820 THEN
            exp_f := 6;
        ELSIF x =- 11819 THEN
            exp_f := 6;
        ELSIF x =- 11818 THEN
            exp_f := 6;
        ELSIF x =- 11817 THEN
            exp_f := 6;
        ELSIF x =- 11816 THEN
            exp_f := 6;
        ELSIF x =- 11815 THEN
            exp_f := 6;
        ELSIF x =- 11814 THEN
            exp_f := 6;
        ELSIF x =- 11813 THEN
            exp_f := 6;
        ELSIF x =- 11812 THEN
            exp_f := 6;
        ELSIF x =- 11811 THEN
            exp_f := 6;
        ELSIF x =- 11810 THEN
            exp_f := 6;
        ELSIF x =- 11809 THEN
            exp_f := 6;
        ELSIF x =- 11808 THEN
            exp_f := 6;
        ELSIF x =- 11807 THEN
            exp_f := 6;
        ELSIF x =- 11806 THEN
            exp_f := 6;
        ELSIF x =- 11805 THEN
            exp_f := 6;
        ELSIF x =- 11804 THEN
            exp_f := 6;
        ELSIF x =- 11803 THEN
            exp_f := 6;
        ELSIF x =- 11802 THEN
            exp_f := 6;
        ELSIF x =- 11801 THEN
            exp_f := 6;
        ELSIF x =- 11800 THEN
            exp_f := 6;
        ELSIF x =- 11799 THEN
            exp_f := 6;
        ELSIF x =- 11798 THEN
            exp_f := 6;
        ELSIF x =- 11797 THEN
            exp_f := 6;
        ELSIF x =- 11796 THEN
            exp_f := 6;
        ELSIF x =- 11795 THEN
            exp_f := 6;
        ELSIF x =- 11794 THEN
            exp_f := 6;
        ELSIF x =- 11793 THEN
            exp_f := 6;
        ELSIF x =- 11792 THEN
            exp_f := 6;
        ELSIF x =- 11791 THEN
            exp_f := 6;
        ELSIF x =- 11790 THEN
            exp_f := 6;
        ELSIF x =- 11789 THEN
            exp_f := 6;
        ELSIF x =- 11788 THEN
            exp_f := 6;
        ELSIF x =- 11787 THEN
            exp_f := 6;
        ELSIF x =- 11786 THEN
            exp_f := 6;
        ELSIF x =- 11785 THEN
            exp_f := 6;
        ELSIF x =- 11784 THEN
            exp_f := 6;
        ELSIF x =- 11783 THEN
            exp_f := 6;
        ELSIF x =- 11782 THEN
            exp_f := 6;
        ELSIF x =- 11781 THEN
            exp_f := 6;
        ELSIF x =- 11780 THEN
            exp_f := 6;
        ELSIF x =- 11779 THEN
            exp_f := 6;
        ELSIF x =- 11778 THEN
            exp_f := 6;
        ELSIF x =- 11777 THEN
            exp_f := 6;
        ELSIF x =- 11776 THEN
            exp_f := 6;
        ELSIF x =- 11775 THEN
            exp_f := 7;
        ELSIF x =- 11774 THEN
            exp_f := 7;
        ELSIF x =- 11773 THEN
            exp_f := 7;
        ELSIF x =- 11772 THEN
            exp_f := 7;
        ELSIF x =- 11771 THEN
            exp_f := 7;
        ELSIF x =- 11770 THEN
            exp_f := 7;
        ELSIF x =- 11769 THEN
            exp_f := 7;
        ELSIF x =- 11768 THEN
            exp_f := 7;
        ELSIF x =- 11767 THEN
            exp_f := 7;
        ELSIF x =- 11766 THEN
            exp_f := 7;
        ELSIF x =- 11765 THEN
            exp_f := 7;
        ELSIF x =- 11764 THEN
            exp_f := 7;
        ELSIF x =- 11763 THEN
            exp_f := 7;
        ELSIF x =- 11762 THEN
            exp_f := 7;
        ELSIF x =- 11761 THEN
            exp_f := 7;
        ELSIF x =- 11760 THEN
            exp_f := 7;
        ELSIF x =- 11759 THEN
            exp_f := 7;
        ELSIF x =- 11758 THEN
            exp_f := 7;
        ELSIF x =- 11757 THEN
            exp_f := 7;
        ELSIF x =- 11756 THEN
            exp_f := 7;
        ELSIF x =- 11755 THEN
            exp_f := 7;
        ELSIF x =- 11754 THEN
            exp_f := 7;
        ELSIF x =- 11753 THEN
            exp_f := 7;
        ELSIF x =- 11752 THEN
            exp_f := 7;
        ELSIF x =- 11751 THEN
            exp_f := 7;
        ELSIF x =- 11750 THEN
            exp_f := 7;
        ELSIF x =- 11749 THEN
            exp_f := 7;
        ELSIF x =- 11748 THEN
            exp_f := 7;
        ELSIF x =- 11747 THEN
            exp_f := 7;
        ELSIF x =- 11746 THEN
            exp_f := 7;
        ELSIF x =- 11745 THEN
            exp_f := 7;
        ELSIF x =- 11744 THEN
            exp_f := 7;
        ELSIF x =- 11743 THEN
            exp_f := 7;
        ELSIF x =- 11742 THEN
            exp_f := 7;
        ELSIF x =- 11741 THEN
            exp_f := 7;
        ELSIF x =- 11740 THEN
            exp_f := 7;
        ELSIF x =- 11739 THEN
            exp_f := 7;
        ELSIF x =- 11738 THEN
            exp_f := 7;
        ELSIF x =- 11737 THEN
            exp_f := 7;
        ELSIF x =- 11736 THEN
            exp_f := 7;
        ELSIF x =- 11735 THEN
            exp_f := 7;
        ELSIF x =- 11734 THEN
            exp_f := 7;
        ELSIF x =- 11733 THEN
            exp_f := 7;
        ELSIF x =- 11732 THEN
            exp_f := 7;
        ELSIF x =- 11731 THEN
            exp_f := 7;
        ELSIF x =- 11730 THEN
            exp_f := 7;
        ELSIF x =- 11729 THEN
            exp_f := 7;
        ELSIF x =- 11728 THEN
            exp_f := 7;
        ELSIF x =- 11727 THEN
            exp_f := 7;
        ELSIF x =- 11726 THEN
            exp_f := 7;
        ELSIF x =- 11725 THEN
            exp_f := 7;
        ELSIF x =- 11724 THEN
            exp_f := 7;
        ELSIF x =- 11723 THEN
            exp_f := 7;
        ELSIF x =- 11722 THEN
            exp_f := 7;
        ELSIF x =- 11721 THEN
            exp_f := 7;
        ELSIF x =- 11720 THEN
            exp_f := 7;
        ELSIF x =- 11719 THEN
            exp_f := 7;
        ELSIF x =- 11718 THEN
            exp_f := 7;
        ELSIF x =- 11717 THEN
            exp_f := 7;
        ELSIF x =- 11716 THEN
            exp_f := 7;
        ELSIF x =- 11715 THEN
            exp_f := 7;
        ELSIF x =- 11714 THEN
            exp_f := 7;
        ELSIF x =- 11713 THEN
            exp_f := 7;
        ELSIF x =- 11712 THEN
            exp_f := 7;
        ELSIF x =- 11711 THEN
            exp_f := 7;
        ELSIF x =- 11710 THEN
            exp_f := 7;
        ELSIF x =- 11709 THEN
            exp_f := 7;
        ELSIF x =- 11708 THEN
            exp_f := 7;
        ELSIF x =- 11707 THEN
            exp_f := 7;
        ELSIF x =- 11706 THEN
            exp_f := 7;
        ELSIF x =- 11705 THEN
            exp_f := 7;
        ELSIF x =- 11704 THEN
            exp_f := 7;
        ELSIF x =- 11703 THEN
            exp_f := 7;
        ELSIF x =- 11702 THEN
            exp_f := 7;
        ELSIF x =- 11701 THEN
            exp_f := 7;
        ELSIF x =- 11700 THEN
            exp_f := 7;
        ELSIF x =- 11699 THEN
            exp_f := 7;
        ELSIF x =- 11698 THEN
            exp_f := 7;
        ELSIF x =- 11697 THEN
            exp_f := 7;
        ELSIF x =- 11696 THEN
            exp_f := 7;
        ELSIF x =- 11695 THEN
            exp_f := 7;
        ELSIF x =- 11694 THEN
            exp_f := 7;
        ELSIF x =- 11693 THEN
            exp_f := 7;
        ELSIF x =- 11692 THEN
            exp_f := 7;
        ELSIF x =- 11691 THEN
            exp_f := 7;
        ELSIF x =- 11690 THEN
            exp_f := 7;
        ELSIF x =- 11689 THEN
            exp_f := 7;
        ELSIF x =- 11688 THEN
            exp_f := 7;
        ELSIF x =- 11687 THEN
            exp_f := 7;
        ELSIF x =- 11686 THEN
            exp_f := 7;
        ELSIF x =- 11685 THEN
            exp_f := 7;
        ELSIF x =- 11684 THEN
            exp_f := 7;
        ELSIF x =- 11683 THEN
            exp_f := 7;
        ELSIF x =- 11682 THEN
            exp_f := 7;
        ELSIF x =- 11681 THEN
            exp_f := 7;
        ELSIF x =- 11680 THEN
            exp_f := 7;
        ELSIF x =- 11679 THEN
            exp_f := 7;
        ELSIF x =- 11678 THEN
            exp_f := 7;
        ELSIF x =- 11677 THEN
            exp_f := 7;
        ELSIF x =- 11676 THEN
            exp_f := 7;
        ELSIF x =- 11675 THEN
            exp_f := 7;
        ELSIF x =- 11674 THEN
            exp_f := 7;
        ELSIF x =- 11673 THEN
            exp_f := 7;
        ELSIF x =- 11672 THEN
            exp_f := 7;
        ELSIF x =- 11671 THEN
            exp_f := 7;
        ELSIF x =- 11670 THEN
            exp_f := 7;
        ELSIF x =- 11669 THEN
            exp_f := 7;
        ELSIF x =- 11668 THEN
            exp_f := 7;
        ELSIF x =- 11667 THEN
            exp_f := 7;
        ELSIF x =- 11666 THEN
            exp_f := 7;
        ELSIF x =- 11665 THEN
            exp_f := 7;
        ELSIF x =- 11664 THEN
            exp_f := 7;
        ELSIF x =- 11663 THEN
            exp_f := 7;
        ELSIF x =- 11662 THEN
            exp_f := 7;
        ELSIF x =- 11661 THEN
            exp_f := 7;
        ELSIF x =- 11660 THEN
            exp_f := 7;
        ELSIF x =- 11659 THEN
            exp_f := 7;
        ELSIF x =- 11658 THEN
            exp_f := 7;
        ELSIF x =- 11657 THEN
            exp_f := 7;
        ELSIF x =- 11656 THEN
            exp_f := 7;
        ELSIF x =- 11655 THEN
            exp_f := 7;
        ELSIF x =- 11654 THEN
            exp_f := 7;
        ELSIF x =- 11653 THEN
            exp_f := 7;
        ELSIF x =- 11652 THEN
            exp_f := 7;
        ELSIF x =- 11651 THEN
            exp_f := 7;
        ELSIF x =- 11650 THEN
            exp_f := 7;
        ELSIF x =- 11649 THEN
            exp_f := 7;
        ELSIF x =- 11648 THEN
            exp_f := 7;
        ELSIF x =- 11647 THEN
            exp_f := 7;
        ELSIF x =- 11646 THEN
            exp_f := 7;
        ELSIF x =- 11645 THEN
            exp_f := 7;
        ELSIF x =- 11644 THEN
            exp_f := 7;
        ELSIF x =- 11643 THEN
            exp_f := 7;
        ELSIF x =- 11642 THEN
            exp_f := 7;
        ELSIF x =- 11641 THEN
            exp_f := 7;
        ELSIF x =- 11640 THEN
            exp_f := 7;
        ELSIF x =- 11639 THEN
            exp_f := 7;
        ELSIF x =- 11638 THEN
            exp_f := 7;
        ELSIF x =- 11637 THEN
            exp_f := 7;
        ELSIF x =- 11636 THEN
            exp_f := 7;
        ELSIF x =- 11635 THEN
            exp_f := 7;
        ELSIF x =- 11634 THEN
            exp_f := 7;
        ELSIF x =- 11633 THEN
            exp_f := 7;
        ELSIF x =- 11632 THEN
            exp_f := 7;
        ELSIF x =- 11631 THEN
            exp_f := 7;
        ELSIF x =- 11630 THEN
            exp_f := 7;
        ELSIF x =- 11629 THEN
            exp_f := 7;
        ELSIF x =- 11628 THEN
            exp_f := 7;
        ELSIF x =- 11627 THEN
            exp_f := 7;
        ELSIF x =- 11626 THEN
            exp_f := 7;
        ELSIF x =- 11625 THEN
            exp_f := 7;
        ELSIF x =- 11624 THEN
            exp_f := 7;
        ELSIF x =- 11623 THEN
            exp_f := 7;
        ELSIF x =- 11622 THEN
            exp_f := 7;
        ELSIF x =- 11621 THEN
            exp_f := 7;
        ELSIF x =- 11620 THEN
            exp_f := 7;
        ELSIF x =- 11619 THEN
            exp_f := 7;
        ELSIF x =- 11618 THEN
            exp_f := 7;
        ELSIF x =- 11617 THEN
            exp_f := 7;
        ELSIF x =- 11616 THEN
            exp_f := 7;
        ELSIF x =- 11615 THEN
            exp_f := 7;
        ELSIF x =- 11614 THEN
            exp_f := 7;
        ELSIF x =- 11613 THEN
            exp_f := 7;
        ELSIF x =- 11612 THEN
            exp_f := 7;
        ELSIF x =- 11611 THEN
            exp_f := 7;
        ELSIF x =- 11610 THEN
            exp_f := 7;
        ELSIF x =- 11609 THEN
            exp_f := 7;
        ELSIF x =- 11608 THEN
            exp_f := 7;
        ELSIF x =- 11607 THEN
            exp_f := 7;
        ELSIF x =- 11606 THEN
            exp_f := 7;
        ELSIF x =- 11605 THEN
            exp_f := 8;
        ELSIF x =- 11604 THEN
            exp_f := 8;
        ELSIF x =- 11603 THEN
            exp_f := 8;
        ELSIF x =- 11602 THEN
            exp_f := 8;
        ELSIF x =- 11601 THEN
            exp_f := 8;
        ELSIF x =- 11600 THEN
            exp_f := 8;
        ELSIF x =- 11599 THEN
            exp_f := 8;
        ELSIF x =- 11598 THEN
            exp_f := 8;
        ELSIF x =- 11597 THEN
            exp_f := 8;
        ELSIF x =- 11596 THEN
            exp_f := 8;
        ELSIF x =- 11595 THEN
            exp_f := 8;
        ELSIF x =- 11594 THEN
            exp_f := 8;
        ELSIF x =- 11593 THEN
            exp_f := 8;
        ELSIF x =- 11592 THEN
            exp_f := 8;
        ELSIF x =- 11591 THEN
            exp_f := 8;
        ELSIF x =- 11590 THEN
            exp_f := 8;
        ELSIF x =- 11589 THEN
            exp_f := 8;
        ELSIF x =- 11588 THEN
            exp_f := 8;
        ELSIF x =- 11587 THEN
            exp_f := 8;
        ELSIF x =- 11586 THEN
            exp_f := 8;
        ELSIF x =- 11585 THEN
            exp_f := 8;
        ELSIF x =- 11584 THEN
            exp_f := 8;
        ELSIF x =- 11583 THEN
            exp_f := 8;
        ELSIF x =- 11582 THEN
            exp_f := 8;
        ELSIF x =- 11581 THEN
            exp_f := 8;
        ELSIF x =- 11580 THEN
            exp_f := 8;
        ELSIF x =- 11579 THEN
            exp_f := 8;
        ELSIF x =- 11578 THEN
            exp_f := 8;
        ELSIF x =- 11577 THEN
            exp_f := 8;
        ELSIF x =- 11576 THEN
            exp_f := 8;
        ELSIF x =- 11575 THEN
            exp_f := 8;
        ELSIF x =- 11574 THEN
            exp_f := 8;
        ELSIF x =- 11573 THEN
            exp_f := 8;
        ELSIF x =- 11572 THEN
            exp_f := 8;
        ELSIF x =- 11571 THEN
            exp_f := 8;
        ELSIF x =- 11570 THEN
            exp_f := 8;
        ELSIF x =- 11569 THEN
            exp_f := 8;
        ELSIF x =- 11568 THEN
            exp_f := 8;
        ELSIF x =- 11567 THEN
            exp_f := 8;
        ELSIF x =- 11566 THEN
            exp_f := 8;
        ELSIF x =- 11565 THEN
            exp_f := 8;
        ELSIF x =- 11564 THEN
            exp_f := 8;
        ELSIF x =- 11563 THEN
            exp_f := 8;
        ELSIF x =- 11562 THEN
            exp_f := 8;
        ELSIF x =- 11561 THEN
            exp_f := 8;
        ELSIF x =- 11560 THEN
            exp_f := 8;
        ELSIF x =- 11559 THEN
            exp_f := 8;
        ELSIF x =- 11558 THEN
            exp_f := 8;
        ELSIF x =- 11557 THEN
            exp_f := 8;
        ELSIF x =- 11556 THEN
            exp_f := 8;
        ELSIF x =- 11555 THEN
            exp_f := 8;
        ELSIF x =- 11554 THEN
            exp_f := 8;
        ELSIF x =- 11553 THEN
            exp_f := 8;
        ELSIF x =- 11552 THEN
            exp_f := 8;
        ELSIF x =- 11551 THEN
            exp_f := 8;
        ELSIF x =- 11550 THEN
            exp_f := 8;
        ELSIF x =- 11549 THEN
            exp_f := 8;
        ELSIF x =- 11548 THEN
            exp_f := 8;
        ELSIF x =- 11547 THEN
            exp_f := 8;
        ELSIF x =- 11546 THEN
            exp_f := 8;
        ELSIF x =- 11545 THEN
            exp_f := 8;
        ELSIF x =- 11544 THEN
            exp_f := 8;
        ELSIF x =- 11543 THEN
            exp_f := 8;
        ELSIF x =- 11542 THEN
            exp_f := 8;
        ELSIF x =- 11541 THEN
            exp_f := 8;
        ELSIF x =- 11540 THEN
            exp_f := 8;
        ELSIF x =- 11539 THEN
            exp_f := 8;
        ELSIF x =- 11538 THEN
            exp_f := 8;
        ELSIF x =- 11537 THEN
            exp_f := 8;
        ELSIF x =- 11536 THEN
            exp_f := 8;
        ELSIF x =- 11535 THEN
            exp_f := 8;
        ELSIF x =- 11534 THEN
            exp_f := 8;
        ELSIF x =- 11533 THEN
            exp_f := 8;
        ELSIF x =- 11532 THEN
            exp_f := 8;
        ELSIF x =- 11531 THEN
            exp_f := 8;
        ELSIF x =- 11530 THEN
            exp_f := 8;
        ELSIF x =- 11529 THEN
            exp_f := 8;
        ELSIF x =- 11528 THEN
            exp_f := 8;
        ELSIF x =- 11527 THEN
            exp_f := 8;
        ELSIF x =- 11526 THEN
            exp_f := 8;
        ELSIF x =- 11525 THEN
            exp_f := 8;
        ELSIF x =- 11524 THEN
            exp_f := 8;
        ELSIF x =- 11523 THEN
            exp_f := 8;
        ELSIF x =- 11522 THEN
            exp_f := 8;
        ELSIF x =- 11521 THEN
            exp_f := 8;
        ELSIF x =- 11520 THEN
            exp_f := 8;
        ELSIF x =- 11519 THEN
            exp_f := 8;
        ELSIF x =- 11518 THEN
            exp_f := 8;
        ELSIF x =- 11517 THEN
            exp_f := 8;
        ELSIF x =- 11516 THEN
            exp_f := 8;
        ELSIF x =- 11515 THEN
            exp_f := 8;
        ELSIF x =- 11514 THEN
            exp_f := 8;
        ELSIF x =- 11513 THEN
            exp_f := 8;
        ELSIF x =- 11512 THEN
            exp_f := 8;
        ELSIF x =- 11511 THEN
            exp_f := 8;
        ELSIF x =- 11510 THEN
            exp_f := 8;
        ELSIF x =- 11509 THEN
            exp_f := 8;
        ELSIF x =- 11508 THEN
            exp_f := 8;
        ELSIF x =- 11507 THEN
            exp_f := 8;
        ELSIF x =- 11506 THEN
            exp_f := 8;
        ELSIF x =- 11505 THEN
            exp_f := 8;
        ELSIF x =- 11504 THEN
            exp_f := 8;
        ELSIF x =- 11503 THEN
            exp_f := 8;
        ELSIF x =- 11502 THEN
            exp_f := 8;
        ELSIF x =- 11501 THEN
            exp_f := 8;
        ELSIF x =- 11500 THEN
            exp_f := 8;
        ELSIF x =- 11499 THEN
            exp_f := 8;
        ELSIF x =- 11498 THEN
            exp_f := 8;
        ELSIF x =- 11497 THEN
            exp_f := 8;
        ELSIF x =- 11496 THEN
            exp_f := 8;
        ELSIF x =- 11495 THEN
            exp_f := 8;
        ELSIF x =- 11494 THEN
            exp_f := 8;
        ELSIF x =- 11493 THEN
            exp_f := 8;
        ELSIF x =- 11492 THEN
            exp_f := 8;
        ELSIF x =- 11491 THEN
            exp_f := 8;
        ELSIF x =- 11490 THEN
            exp_f := 8;
        ELSIF x =- 11489 THEN
            exp_f := 8;
        ELSIF x =- 11488 THEN
            exp_f := 8;
        ELSIF x =- 11487 THEN
            exp_f := 8;
        ELSIF x =- 11486 THEN
            exp_f := 8;
        ELSIF x =- 11485 THEN
            exp_f := 8;
        ELSIF x =- 11484 THEN
            exp_f := 8;
        ELSIF x =- 11483 THEN
            exp_f := 8;
        ELSIF x =- 11482 THEN
            exp_f := 8;
        ELSIF x =- 11481 THEN
            exp_f := 8;
        ELSIF x =- 11480 THEN
            exp_f := 8;
        ELSIF x =- 11479 THEN
            exp_f := 8;
        ELSIF x =- 11478 THEN
            exp_f := 8;
        ELSIF x =- 11477 THEN
            exp_f := 8;
        ELSIF x =- 11476 THEN
            exp_f := 8;
        ELSIF x =- 11475 THEN
            exp_f := 8;
        ELSIF x =- 11474 THEN
            exp_f := 8;
        ELSIF x =- 11473 THEN
            exp_f := 8;
        ELSIF x =- 11472 THEN
            exp_f := 8;
        ELSIF x =- 11471 THEN
            exp_f := 8;
        ELSIF x =- 11470 THEN
            exp_f := 8;
        ELSIF x =- 11469 THEN
            exp_f := 8;
        ELSIF x =- 11468 THEN
            exp_f := 8;
        ELSIF x =- 11467 THEN
            exp_f := 8;
        ELSIF x =- 11466 THEN
            exp_f := 8;
        ELSIF x =- 11465 THEN
            exp_f := 8;
        ELSIF x =- 11464 THEN
            exp_f := 8;
        ELSIF x =- 11463 THEN
            exp_f := 8;
        ELSIF x =- 11462 THEN
            exp_f := 8;
        ELSIF x =- 11461 THEN
            exp_f := 8;
        ELSIF x =- 11460 THEN
            exp_f := 8;
        ELSIF x =- 11459 THEN
            exp_f := 8;
        ELSIF x =- 11458 THEN
            exp_f := 8;
        ELSIF x =- 11457 THEN
            exp_f := 8;
        ELSIF x =- 11456 THEN
            exp_f := 8;
        ELSIF x =- 11455 THEN
            exp_f := 8;
        ELSIF x =- 11454 THEN
            exp_f := 8;
        ELSIF x =- 11453 THEN
            exp_f := 8;
        ELSIF x =- 11452 THEN
            exp_f := 8;
        ELSIF x =- 11451 THEN
            exp_f := 8;
        ELSIF x =- 11450 THEN
            exp_f := 8;
        ELSIF x =- 11449 THEN
            exp_f := 8;
        ELSIF x =- 11448 THEN
            exp_f := 8;
        ELSIF x =- 11447 THEN
            exp_f := 8;
        ELSIF x =- 11446 THEN
            exp_f := 8;
        ELSIF x =- 11445 THEN
            exp_f := 8;
        ELSIF x =- 11444 THEN
            exp_f := 8;
        ELSIF x =- 11443 THEN
            exp_f := 8;
        ELSIF x =- 11442 THEN
            exp_f := 8;
        ELSIF x =- 11441 THEN
            exp_f := 8;
        ELSIF x =- 11440 THEN
            exp_f := 8;
        ELSIF x =- 11439 THEN
            exp_f := 8;
        ELSIF x =- 11438 THEN
            exp_f := 8;
        ELSIF x =- 11437 THEN
            exp_f := 8;
        ELSIF x =- 11436 THEN
            exp_f := 8;
        ELSIF x =- 11435 THEN
            exp_f := 8;
        ELSIF x =- 11434 THEN
            exp_f := 8;
        ELSIF x =- 11433 THEN
            exp_f := 8;
        ELSIF x =- 11432 THEN
            exp_f := 8;
        ELSIF x =- 11431 THEN
            exp_f := 8;
        ELSIF x =- 11430 THEN
            exp_f := 8;
        ELSIF x =- 11429 THEN
            exp_f := 8;
        ELSIF x =- 11428 THEN
            exp_f := 8;
        ELSIF x =- 11427 THEN
            exp_f := 8;
        ELSIF x =- 11426 THEN
            exp_f := 8;
        ELSIF x =- 11425 THEN
            exp_f := 8;
        ELSIF x =- 11424 THEN
            exp_f := 8;
        ELSIF x =- 11423 THEN
            exp_f := 8;
        ELSIF x =- 11422 THEN
            exp_f := 8;
        ELSIF x =- 11421 THEN
            exp_f := 8;
        ELSIF x =- 11420 THEN
            exp_f := 8;
        ELSIF x =- 11419 THEN
            exp_f := 8;
        ELSIF x =- 11418 THEN
            exp_f := 8;
        ELSIF x =- 11417 THEN
            exp_f := 8;
        ELSIF x =- 11416 THEN
            exp_f := 8;
        ELSIF x =- 11415 THEN
            exp_f := 8;
        ELSIF x =- 11414 THEN
            exp_f := 8;
        ELSIF x =- 11413 THEN
            exp_f := 8;
        ELSIF x =- 11412 THEN
            exp_f := 8;
        ELSIF x =- 11411 THEN
            exp_f := 8;
        ELSIF x =- 11410 THEN
            exp_f := 8;
        ELSIF x =- 11409 THEN
            exp_f := 8;
        ELSIF x =- 11408 THEN
            exp_f := 8;
        ELSIF x =- 11407 THEN
            exp_f := 8;
        ELSIF x =- 11406 THEN
            exp_f := 8;
        ELSIF x =- 11405 THEN
            exp_f := 8;
        ELSIF x =- 11404 THEN
            exp_f := 8;
        ELSIF x =- 11403 THEN
            exp_f := 8;
        ELSIF x =- 11402 THEN
            exp_f := 8;
        ELSIF x =- 11401 THEN
            exp_f := 8;
        ELSIF x =- 11400 THEN
            exp_f := 8;
        ELSIF x =- 11399 THEN
            exp_f := 8;
        ELSIF x =- 11398 THEN
            exp_f := 8;
        ELSIF x =- 11397 THEN
            exp_f := 8;
        ELSIF x =- 11396 THEN
            exp_f := 8;
        ELSIF x =- 11395 THEN
            exp_f := 8;
        ELSIF x =- 11394 THEN
            exp_f := 8;
        ELSIF x =- 11393 THEN
            exp_f := 8;
        ELSIF x =- 11392 THEN
            exp_f := 8;
        ELSIF x =- 11391 THEN
            exp_f := 8;
        ELSIF x =- 11390 THEN
            exp_f := 8;
        ELSIF x =- 11389 THEN
            exp_f := 8;
        ELSIF x =- 11388 THEN
            exp_f := 8;
        ELSIF x =- 11387 THEN
            exp_f := 8;
        ELSIF x =- 11386 THEN
            exp_f := 8;
        ELSIF x =- 11385 THEN
            exp_f := 8;
        ELSIF x =- 11384 THEN
            exp_f := 8;
        ELSIF x =- 11383 THEN
            exp_f := 8;
        ELSIF x =- 11382 THEN
            exp_f := 8;
        ELSIF x =- 11381 THEN
            exp_f := 8;
        ELSIF x =- 11380 THEN
            exp_f := 8;
        ELSIF x =- 11379 THEN
            exp_f := 8;
        ELSIF x =- 11378 THEN
            exp_f := 8;
        ELSIF x =- 11377 THEN
            exp_f := 9;
        ELSIF x =- 11376 THEN
            exp_f := 9;
        ELSIF x =- 11375 THEN
            exp_f := 9;
        ELSIF x =- 11374 THEN
            exp_f := 9;
        ELSIF x =- 11373 THEN
            exp_f := 9;
        ELSIF x =- 11372 THEN
            exp_f := 9;
        ELSIF x =- 11371 THEN
            exp_f := 9;
        ELSIF x =- 11370 THEN
            exp_f := 9;
        ELSIF x =- 11369 THEN
            exp_f := 9;
        ELSIF x =- 11368 THEN
            exp_f := 9;
        ELSIF x =- 11367 THEN
            exp_f := 9;
        ELSIF x =- 11366 THEN
            exp_f := 9;
        ELSIF x =- 11365 THEN
            exp_f := 9;
        ELSIF x =- 11364 THEN
            exp_f := 9;
        ELSIF x =- 11363 THEN
            exp_f := 9;
        ELSIF x =- 11362 THEN
            exp_f := 9;
        ELSIF x =- 11361 THEN
            exp_f := 9;
        ELSIF x =- 11360 THEN
            exp_f := 9;
        ELSIF x =- 11359 THEN
            exp_f := 9;
        ELSIF x =- 11358 THEN
            exp_f := 9;
        ELSIF x =- 11357 THEN
            exp_f := 9;
        ELSIF x =- 11356 THEN
            exp_f := 9;
        ELSIF x =- 11355 THEN
            exp_f := 9;
        ELSIF x =- 11354 THEN
            exp_f := 9;
        ELSIF x =- 11353 THEN
            exp_f := 9;
        ELSIF x =- 11352 THEN
            exp_f := 9;
        ELSIF x =- 11351 THEN
            exp_f := 9;
        ELSIF x =- 11350 THEN
            exp_f := 9;
        ELSIF x =- 11349 THEN
            exp_f := 9;
        ELSIF x =- 11348 THEN
            exp_f := 9;
        ELSIF x =- 11347 THEN
            exp_f := 9;
        ELSIF x =- 11346 THEN
            exp_f := 9;
        ELSIF x =- 11345 THEN
            exp_f := 9;
        ELSIF x =- 11344 THEN
            exp_f := 9;
        ELSIF x =- 11343 THEN
            exp_f := 9;
        ELSIF x =- 11342 THEN
            exp_f := 9;
        ELSIF x =- 11341 THEN
            exp_f := 9;
        ELSIF x =- 11340 THEN
            exp_f := 9;
        ELSIF x =- 11339 THEN
            exp_f := 9;
        ELSIF x =- 11338 THEN
            exp_f := 9;
        ELSIF x =- 11337 THEN
            exp_f := 9;
        ELSIF x =- 11336 THEN
            exp_f := 9;
        ELSIF x =- 11335 THEN
            exp_f := 9;
        ELSIF x =- 11334 THEN
            exp_f := 9;
        ELSIF x =- 11333 THEN
            exp_f := 9;
        ELSIF x =- 11332 THEN
            exp_f := 9;
        ELSIF x =- 11331 THEN
            exp_f := 9;
        ELSIF x =- 11330 THEN
            exp_f := 9;
        ELSIF x =- 11329 THEN
            exp_f := 9;
        ELSIF x =- 11328 THEN
            exp_f := 9;
        ELSIF x =- 11327 THEN
            exp_f := 9;
        ELSIF x =- 11326 THEN
            exp_f := 9;
        ELSIF x =- 11325 THEN
            exp_f := 9;
        ELSIF x =- 11324 THEN
            exp_f := 9;
        ELSIF x =- 11323 THEN
            exp_f := 9;
        ELSIF x =- 11322 THEN
            exp_f := 9;
        ELSIF x =- 11321 THEN
            exp_f := 9;
        ELSIF x =- 11320 THEN
            exp_f := 9;
        ELSIF x =- 11319 THEN
            exp_f := 9;
        ELSIF x =- 11318 THEN
            exp_f := 9;
        ELSIF x =- 11317 THEN
            exp_f := 9;
        ELSIF x =- 11316 THEN
            exp_f := 9;
        ELSIF x =- 11315 THEN
            exp_f := 9;
        ELSIF x =- 11314 THEN
            exp_f := 9;
        ELSIF x =- 11313 THEN
            exp_f := 9;
        ELSIF x =- 11312 THEN
            exp_f := 9;
        ELSIF x =- 11311 THEN
            exp_f := 9;
        ELSIF x =- 11310 THEN
            exp_f := 9;
        ELSIF x =- 11309 THEN
            exp_f := 9;
        ELSIF x =- 11308 THEN
            exp_f := 9;
        ELSIF x =- 11307 THEN
            exp_f := 9;
        ELSIF x =- 11306 THEN
            exp_f := 9;
        ELSIF x =- 11305 THEN
            exp_f := 9;
        ELSIF x =- 11304 THEN
            exp_f := 9;
        ELSIF x =- 11303 THEN
            exp_f := 9;
        ELSIF x =- 11302 THEN
            exp_f := 9;
        ELSIF x =- 11301 THEN
            exp_f := 9;
        ELSIF x =- 11300 THEN
            exp_f := 9;
        ELSIF x =- 11299 THEN
            exp_f := 9;
        ELSIF x =- 11298 THEN
            exp_f := 9;
        ELSIF x =- 11297 THEN
            exp_f := 9;
        ELSIF x =- 11296 THEN
            exp_f := 9;
        ELSIF x =- 11295 THEN
            exp_f := 9;
        ELSIF x =- 11294 THEN
            exp_f := 9;
        ELSIF x =- 11293 THEN
            exp_f := 9;
        ELSIF x =- 11292 THEN
            exp_f := 9;
        ELSIF x =- 11291 THEN
            exp_f := 9;
        ELSIF x =- 11290 THEN
            exp_f := 9;
        ELSIF x =- 11289 THEN
            exp_f := 9;
        ELSIF x =- 11288 THEN
            exp_f := 9;
        ELSIF x =- 11287 THEN
            exp_f := 9;
        ELSIF x =- 11286 THEN
            exp_f := 9;
        ELSIF x =- 11285 THEN
            exp_f := 9;
        ELSIF x =- 11284 THEN
            exp_f := 9;
        ELSIF x =- 11283 THEN
            exp_f := 9;
        ELSIF x =- 11282 THEN
            exp_f := 9;
        ELSIF x =- 11281 THEN
            exp_f := 9;
        ELSIF x =- 11280 THEN
            exp_f := 9;
        ELSIF x =- 11279 THEN
            exp_f := 9;
        ELSIF x =- 11278 THEN
            exp_f := 9;
        ELSIF x =- 11277 THEN
            exp_f := 9;
        ELSIF x =- 11276 THEN
            exp_f := 9;
        ELSIF x =- 11275 THEN
            exp_f := 9;
        ELSIF x =- 11274 THEN
            exp_f := 9;
        ELSIF x =- 11273 THEN
            exp_f := 9;
        ELSIF x =- 11272 THEN
            exp_f := 9;
        ELSIF x =- 11271 THEN
            exp_f := 9;
        ELSIF x =- 11270 THEN
            exp_f := 9;
        ELSIF x =- 11269 THEN
            exp_f := 9;
        ELSIF x =- 11268 THEN
            exp_f := 9;
        ELSIF x =- 11267 THEN
            exp_f := 9;
        ELSIF x =- 11266 THEN
            exp_f := 9;
        ELSIF x =- 11265 THEN
            exp_f := 9;
        ELSIF x =- 11264 THEN
            exp_f := 9;
        ELSIF x =- 11263 THEN
            exp_f := 9;
        ELSIF x =- 11262 THEN
            exp_f := 9;
        ELSIF x =- 11261 THEN
            exp_f := 9;
        ELSIF x =- 11260 THEN
            exp_f := 9;
        ELSIF x =- 11259 THEN
            exp_f := 9;
        ELSIF x =- 11258 THEN
            exp_f := 9;
        ELSIF x =- 11257 THEN
            exp_f := 9;
        ELSIF x =- 11256 THEN
            exp_f := 9;
        ELSIF x =- 11255 THEN
            exp_f := 9;
        ELSIF x =- 11254 THEN
            exp_f := 9;
        ELSIF x =- 11253 THEN
            exp_f := 9;
        ELSIF x =- 11252 THEN
            exp_f := 9;
        ELSIF x =- 11251 THEN
            exp_f := 9;
        ELSIF x =- 11250 THEN
            exp_f := 9;
        ELSIF x =- 11249 THEN
            exp_f := 9;
        ELSIF x =- 11248 THEN
            exp_f := 9;
        ELSIF x =- 11247 THEN
            exp_f := 9;
        ELSIF x =- 11246 THEN
            exp_f := 9;
        ELSIF x =- 11245 THEN
            exp_f := 9;
        ELSIF x =- 11244 THEN
            exp_f := 9;
        ELSIF x =- 11243 THEN
            exp_f := 9;
        ELSIF x =- 11242 THEN
            exp_f := 9;
        ELSIF x =- 11241 THEN
            exp_f := 9;
        ELSIF x =- 11240 THEN
            exp_f := 9;
        ELSIF x =- 11239 THEN
            exp_f := 9;
        ELSIF x =- 11238 THEN
            exp_f := 9;
        ELSIF x =- 11237 THEN
            exp_f := 9;
        ELSIF x =- 11236 THEN
            exp_f := 9;
        ELSIF x =- 11235 THEN
            exp_f := 9;
        ELSIF x =- 11234 THEN
            exp_f := 9;
        ELSIF x =- 11233 THEN
            exp_f := 9;
        ELSIF x =- 11232 THEN
            exp_f := 9;
        ELSIF x =- 11231 THEN
            exp_f := 9;
        ELSIF x =- 11230 THEN
            exp_f := 9;
        ELSIF x =- 11229 THEN
            exp_f := 9;
        ELSIF x =- 11228 THEN
            exp_f := 9;
        ELSIF x =- 11227 THEN
            exp_f := 9;
        ELSIF x =- 11226 THEN
            exp_f := 9;
        ELSIF x =- 11225 THEN
            exp_f := 9;
        ELSIF x =- 11224 THEN
            exp_f := 9;
        ELSIF x =- 11223 THEN
            exp_f := 9;
        ELSIF x =- 11222 THEN
            exp_f := 9;
        ELSIF x =- 11221 THEN
            exp_f := 9;
        ELSIF x =- 11220 THEN
            exp_f := 9;
        ELSIF x =- 11219 THEN
            exp_f := 9;
        ELSIF x =- 11218 THEN
            exp_f := 9;
        ELSIF x =- 11217 THEN
            exp_f := 9;
        ELSIF x =- 11216 THEN
            exp_f := 9;
        ELSIF x =- 11215 THEN
            exp_f := 9;
        ELSIF x =- 11214 THEN
            exp_f := 9;
        ELSIF x =- 11213 THEN
            exp_f := 9;
        ELSIF x =- 11212 THEN
            exp_f := 9;
        ELSIF x =- 11211 THEN
            exp_f := 9;
        ELSIF x =- 11210 THEN
            exp_f := 9;
        ELSIF x =- 11209 THEN
            exp_f := 9;
        ELSIF x =- 11208 THEN
            exp_f := 9;
        ELSIF x =- 11207 THEN
            exp_f := 9;
        ELSIF x =- 11206 THEN
            exp_f := 9;
        ELSIF x =- 11205 THEN
            exp_f := 9;
        ELSIF x =- 11204 THEN
            exp_f := 9;
        ELSIF x =- 11203 THEN
            exp_f := 9;
        ELSIF x =- 11202 THEN
            exp_f := 9;
        ELSIF x =- 11201 THEN
            exp_f := 9;
        ELSIF x =- 11200 THEN
            exp_f := 9;
        ELSIF x =- 11199 THEN
            exp_f := 9;
        ELSIF x =- 11198 THEN
            exp_f := 9;
        ELSIF x =- 11197 THEN
            exp_f := 9;
        ELSIF x =- 11196 THEN
            exp_f := 9;
        ELSIF x =- 11195 THEN
            exp_f := 9;
        ELSIF x =- 11194 THEN
            exp_f := 9;
        ELSIF x =- 11193 THEN
            exp_f := 9;
        ELSIF x =- 11192 THEN
            exp_f := 9;
        ELSIF x =- 11191 THEN
            exp_f := 9;
        ELSIF x =- 11190 THEN
            exp_f := 9;
        ELSIF x =- 11189 THEN
            exp_f := 9;
        ELSIF x =- 11188 THEN
            exp_f := 9;
        ELSIF x =- 11187 THEN
            exp_f := 9;
        ELSIF x =- 11186 THEN
            exp_f := 9;
        ELSIF x =- 11185 THEN
            exp_f := 9;
        ELSIF x =- 11184 THEN
            exp_f := 9;
        ELSIF x =- 11183 THEN
            exp_f := 9;
        ELSIF x =- 11182 THEN
            exp_f := 9;
        ELSIF x =- 11181 THEN
            exp_f := 9;
        ELSIF x =- 11180 THEN
            exp_f := 9;
        ELSIF x =- 11179 THEN
            exp_f := 9;
        ELSIF x =- 11178 THEN
            exp_f := 9;
        ELSIF x =- 11177 THEN
            exp_f := 9;
        ELSIF x =- 11176 THEN
            exp_f := 9;
        ELSIF x =- 11175 THEN
            exp_f := 9;
        ELSIF x =- 11174 THEN
            exp_f := 9;
        ELSIF x =- 11173 THEN
            exp_f := 9;
        ELSIF x =- 11172 THEN
            exp_f := 9;
        ELSIF x =- 11171 THEN
            exp_f := 9;
        ELSIF x =- 11170 THEN
            exp_f := 9;
        ELSIF x =- 11169 THEN
            exp_f := 9;
        ELSIF x =- 11168 THEN
            exp_f := 9;
        ELSIF x =- 11167 THEN
            exp_f := 9;
        ELSIF x =- 11166 THEN
            exp_f := 9;
        ELSIF x =- 11165 THEN
            exp_f := 9;
        ELSIF x =- 11164 THEN
            exp_f := 9;
        ELSIF x =- 11163 THEN
            exp_f := 9;
        ELSIF x =- 11162 THEN
            exp_f := 9;
        ELSIF x =- 11161 THEN
            exp_f := 9;
        ELSIF x =- 11160 THEN
            exp_f := 9;
        ELSIF x =- 11159 THEN
            exp_f := 9;
        ELSIF x =- 11158 THEN
            exp_f := 9;
        ELSIF x =- 11157 THEN
            exp_f := 9;
        ELSIF x =- 11156 THEN
            exp_f := 9;
        ELSIF x =- 11155 THEN
            exp_f := 9;
        ELSIF x =- 11154 THEN
            exp_f := 9;
        ELSIF x =- 11153 THEN
            exp_f := 9;
        ELSIF x =- 11152 THEN
            exp_f := 9;
        ELSIF x =- 11151 THEN
            exp_f := 9;
        ELSIF x =- 11150 THEN
            exp_f := 9;
        ELSIF x =- 11149 THEN
            exp_f := 9;
        ELSIF x =- 11148 THEN
            exp_f := 9;
        ELSIF x =- 11147 THEN
            exp_f := 9;
        ELSIF x =- 11146 THEN
            exp_f := 9;
        ELSIF x =- 11145 THEN
            exp_f := 9;
        ELSIF x =- 11144 THEN
            exp_f := 9;
        ELSIF x =- 11143 THEN
            exp_f := 9;
        ELSIF x =- 11142 THEN
            exp_f := 9;
        ELSIF x =- 11141 THEN
            exp_f := 9;
        ELSIF x =- 11140 THEN
            exp_f := 9;
        ELSIF x =- 11139 THEN
            exp_f := 9;
        ELSIF x =- 11138 THEN
            exp_f := 9;
        ELSIF x =- 11137 THEN
            exp_f := 9;
        ELSIF x =- 11136 THEN
            exp_f := 9;
        ELSIF x =- 11135 THEN
            exp_f := 9;
        ELSIF x =- 11134 THEN
            exp_f := 9;
        ELSIF x =- 11133 THEN
            exp_f := 9;
        ELSIF x =- 11132 THEN
            exp_f := 9;
        ELSIF x =- 11131 THEN
            exp_f := 9;
        ELSIF x =- 11130 THEN
            exp_f := 9;
        ELSIF x =- 11129 THEN
            exp_f := 9;
        ELSIF x =- 11128 THEN
            exp_f := 9;
        ELSIF x =- 11127 THEN
            exp_f := 9;
        ELSIF x =- 11126 THEN
            exp_f := 9;
        ELSIF x =- 11125 THEN
            exp_f := 9;
        ELSIF x =- 11124 THEN
            exp_f := 9;
        ELSIF x =- 11123 THEN
            exp_f := 9;
        ELSIF x =- 11122 THEN
            exp_f := 9;
        ELSIF x =- 11121 THEN
            exp_f := 9;
        ELSIF x =- 11120 THEN
            exp_f := 9;
        ELSIF x =- 11119 THEN
            exp_f := 9;
        ELSIF x =- 11118 THEN
            exp_f := 9;
        ELSIF x =- 11117 THEN
            exp_f := 9;
        ELSIF x =- 11116 THEN
            exp_f := 9;
        ELSIF x =- 11115 THEN
            exp_f := 9;
        ELSIF x =- 11114 THEN
            exp_f := 9;
        ELSIF x =- 11113 THEN
            exp_f := 9;
        ELSIF x =- 11112 THEN
            exp_f := 9;
        ELSIF x =- 11111 THEN
            exp_f := 9;
        ELSIF x =- 11110 THEN
            exp_f := 9;
        ELSIF x =- 11109 THEN
            exp_f := 9;
        ELSIF x =- 11108 THEN
            exp_f := 9;
        ELSIF x =- 11107 THEN
            exp_f := 9;
        ELSIF x =- 11106 THEN
            exp_f := 9;
        ELSIF x =- 11105 THEN
            exp_f := 9;
        ELSIF x =- 11104 THEN
            exp_f := 9;
        ELSIF x =- 11103 THEN
            exp_f := 9;
        ELSIF x =- 11102 THEN
            exp_f := 9;
        ELSIF x =- 11101 THEN
            exp_f := 9;
        ELSIF x =- 11100 THEN
            exp_f := 9;
        ELSIF x =- 11099 THEN
            exp_f := 9;
        ELSIF x =- 11098 THEN
            exp_f := 9;
        ELSIF x =- 11097 THEN
            exp_f := 9;
        ELSIF x =- 11096 THEN
            exp_f := 9;
        ELSIF x =- 11095 THEN
            exp_f := 9;
        ELSIF x =- 11094 THEN
            exp_f := 9;
        ELSIF x =- 11093 THEN
            exp_f := 10;
        ELSIF x =- 11092 THEN
            exp_f := 10;
        ELSIF x =- 11091 THEN
            exp_f := 10;
        ELSIF x =- 11090 THEN
            exp_f := 10;
        ELSIF x =- 11089 THEN
            exp_f := 10;
        ELSIF x =- 11088 THEN
            exp_f := 10;
        ELSIF x =- 11087 THEN
            exp_f := 10;
        ELSIF x =- 11086 THEN
            exp_f := 10;
        ELSIF x =- 11085 THEN
            exp_f := 10;
        ELSIF x =- 11084 THEN
            exp_f := 10;
        ELSIF x =- 11083 THEN
            exp_f := 10;
        ELSIF x =- 11082 THEN
            exp_f := 10;
        ELSIF x =- 11081 THEN
            exp_f := 10;
        ELSIF x =- 11080 THEN
            exp_f := 10;
        ELSIF x =- 11079 THEN
            exp_f := 10;
        ELSIF x =- 11078 THEN
            exp_f := 10;
        ELSIF x =- 11077 THEN
            exp_f := 10;
        ELSIF x =- 11076 THEN
            exp_f := 10;
        ELSIF x =- 11075 THEN
            exp_f := 10;
        ELSIF x =- 11074 THEN
            exp_f := 10;
        ELSIF x =- 11073 THEN
            exp_f := 10;
        ELSIF x =- 11072 THEN
            exp_f := 10;
        ELSIF x =- 11071 THEN
            exp_f := 10;
        ELSIF x =- 11070 THEN
            exp_f := 10;
        ELSIF x =- 11069 THEN
            exp_f := 10;
        ELSIF x =- 11068 THEN
            exp_f := 10;
        ELSIF x =- 11067 THEN
            exp_f := 10;
        ELSIF x =- 11066 THEN
            exp_f := 10;
        ELSIF x =- 11065 THEN
            exp_f := 10;
        ELSIF x =- 11064 THEN
            exp_f := 10;
        ELSIF x =- 11063 THEN
            exp_f := 10;
        ELSIF x =- 11062 THEN
            exp_f := 10;
        ELSIF x =- 11061 THEN
            exp_f := 10;
        ELSIF x =- 11060 THEN
            exp_f := 10;
        ELSIF x =- 11059 THEN
            exp_f := 10;
        ELSIF x =- 11058 THEN
            exp_f := 10;
        ELSIF x =- 11057 THEN
            exp_f := 10;
        ELSIF x =- 11056 THEN
            exp_f := 10;
        ELSIF x =- 11055 THEN
            exp_f := 10;
        ELSIF x =- 11054 THEN
            exp_f := 10;
        ELSIF x =- 11053 THEN
            exp_f := 10;
        ELSIF x =- 11052 THEN
            exp_f := 10;
        ELSIF x =- 11051 THEN
            exp_f := 10;
        ELSIF x =- 11050 THEN
            exp_f := 10;
        ELSIF x =- 11049 THEN
            exp_f := 10;
        ELSIF x =- 11048 THEN
            exp_f := 10;
        ELSIF x =- 11047 THEN
            exp_f := 10;
        ELSIF x =- 11046 THEN
            exp_f := 10;
        ELSIF x =- 11045 THEN
            exp_f := 10;
        ELSIF x =- 11044 THEN
            exp_f := 10;
        ELSIF x =- 11043 THEN
            exp_f := 10;
        ELSIF x =- 11042 THEN
            exp_f := 10;
        ELSIF x =- 11041 THEN
            exp_f := 10;
        ELSIF x =- 11040 THEN
            exp_f := 10;
        ELSIF x =- 11039 THEN
            exp_f := 10;
        ELSIF x =- 11038 THEN
            exp_f := 10;
        ELSIF x =- 11037 THEN
            exp_f := 10;
        ELSIF x =- 11036 THEN
            exp_f := 10;
        ELSIF x =- 11035 THEN
            exp_f := 10;
        ELSIF x =- 11034 THEN
            exp_f := 10;
        ELSIF x =- 11033 THEN
            exp_f := 10;
        ELSIF x =- 11032 THEN
            exp_f := 10;
        ELSIF x =- 11031 THEN
            exp_f := 10;
        ELSIF x =- 11030 THEN
            exp_f := 10;
        ELSIF x =- 11029 THEN
            exp_f := 10;
        ELSIF x =- 11028 THEN
            exp_f := 10;
        ELSIF x =- 11027 THEN
            exp_f := 10;
        ELSIF x =- 11026 THEN
            exp_f := 10;
        ELSIF x =- 11025 THEN
            exp_f := 10;
        ELSIF x =- 11024 THEN
            exp_f := 10;
        ELSIF x =- 11023 THEN
            exp_f := 10;
        ELSIF x =- 11022 THEN
            exp_f := 10;
        ELSIF x =- 11021 THEN
            exp_f := 10;
        ELSIF x =- 11020 THEN
            exp_f := 10;
        ELSIF x =- 11019 THEN
            exp_f := 10;
        ELSIF x =- 11018 THEN
            exp_f := 10;
        ELSIF x =- 11017 THEN
            exp_f := 10;
        ELSIF x =- 11016 THEN
            exp_f := 10;
        ELSIF x =- 11015 THEN
            exp_f := 10;
        ELSIF x =- 11014 THEN
            exp_f := 10;
        ELSIF x =- 11013 THEN
            exp_f := 10;
        ELSIF x =- 11012 THEN
            exp_f := 10;
        ELSIF x =- 11011 THEN
            exp_f := 10;
        ELSIF x =- 11010 THEN
            exp_f := 10;
        ELSIF x =- 11009 THEN
            exp_f := 10;
        ELSIF x =- 11008 THEN
            exp_f := 10;
        ELSIF x =- 11007 THEN
            exp_f := 10;
        ELSIF x =- 11006 THEN
            exp_f := 10;
        ELSIF x =- 11005 THEN
            exp_f := 10;
        ELSIF x =- 11004 THEN
            exp_f := 10;
        ELSIF x =- 11003 THEN
            exp_f := 10;
        ELSIF x =- 11002 THEN
            exp_f := 10;
        ELSIF x =- 11001 THEN
            exp_f := 10;
        ELSIF x =- 11000 THEN
            exp_f := 10;
        ELSIF x =- 10999 THEN
            exp_f := 10;
        ELSIF x =- 10998 THEN
            exp_f := 10;
        ELSIF x =- 10997 THEN
            exp_f := 10;
        ELSIF x =- 10996 THEN
            exp_f := 10;
        ELSIF x =- 10995 THEN
            exp_f := 10;
        ELSIF x =- 10994 THEN
            exp_f := 10;
        ELSIF x =- 10993 THEN
            exp_f := 10;
        ELSIF x =- 10992 THEN
            exp_f := 10;
        ELSIF x =- 10991 THEN
            exp_f := 10;
        ELSIF x =- 10990 THEN
            exp_f := 10;
        ELSIF x =- 10989 THEN
            exp_f := 10;
        ELSIF x =- 10988 THEN
            exp_f := 10;
        ELSIF x =- 10987 THEN
            exp_f := 10;
        ELSIF x =- 10986 THEN
            exp_f := 10;
        ELSIF x =- 10985 THEN
            exp_f := 10;
        ELSIF x =- 10984 THEN
            exp_f := 10;
        ELSIF x =- 10983 THEN
            exp_f := 10;
        ELSIF x =- 10982 THEN
            exp_f := 10;
        ELSIF x =- 10981 THEN
            exp_f := 10;
        ELSIF x =- 10980 THEN
            exp_f := 10;
        ELSIF x =- 10979 THEN
            exp_f := 10;
        ELSIF x =- 10978 THEN
            exp_f := 10;
        ELSIF x =- 10977 THEN
            exp_f := 10;
        ELSIF x =- 10976 THEN
            exp_f := 10;
        ELSIF x =- 10975 THEN
            exp_f := 10;
        ELSIF x =- 10974 THEN
            exp_f := 10;
        ELSIF x =- 10973 THEN
            exp_f := 10;
        ELSIF x =- 10972 THEN
            exp_f := 10;
        ELSIF x =- 10971 THEN
            exp_f := 10;
        ELSIF x =- 10970 THEN
            exp_f := 10;
        ELSIF x =- 10969 THEN
            exp_f := 10;
        ELSIF x =- 10968 THEN
            exp_f := 10;
        ELSIF x =- 10967 THEN
            exp_f := 10;
        ELSIF x =- 10966 THEN
            exp_f := 10;
        ELSIF x =- 10965 THEN
            exp_f := 10;
        ELSIF x =- 10964 THEN
            exp_f := 10;
        ELSIF x =- 10963 THEN
            exp_f := 10;
        ELSIF x =- 10962 THEN
            exp_f := 10;
        ELSIF x =- 10961 THEN
            exp_f := 10;
        ELSIF x =- 10960 THEN
            exp_f := 10;
        ELSIF x =- 10959 THEN
            exp_f := 10;
        ELSIF x =- 10958 THEN
            exp_f := 10;
        ELSIF x =- 10957 THEN
            exp_f := 10;
        ELSIF x =- 10956 THEN
            exp_f := 10;
        ELSIF x =- 10955 THEN
            exp_f := 10;
        ELSIF x =- 10954 THEN
            exp_f := 10;
        ELSIF x =- 10953 THEN
            exp_f := 10;
        ELSIF x =- 10952 THEN
            exp_f := 10;
        ELSIF x =- 10951 THEN
            exp_f := 10;
        ELSIF x =- 10950 THEN
            exp_f := 10;
        ELSIF x =- 10949 THEN
            exp_f := 10;
        ELSIF x =- 10948 THEN
            exp_f := 10;
        ELSIF x =- 10947 THEN
            exp_f := 10;
        ELSIF x =- 10946 THEN
            exp_f := 10;
        ELSIF x =- 10945 THEN
            exp_f := 10;
        ELSIF x =- 10944 THEN
            exp_f := 10;
        ELSIF x =- 10943 THEN
            exp_f := 10;
        ELSIF x =- 10942 THEN
            exp_f := 10;
        ELSIF x =- 10941 THEN
            exp_f := 10;
        ELSIF x =- 10940 THEN
            exp_f := 10;
        ELSIF x =- 10939 THEN
            exp_f := 10;
        ELSIF x =- 10938 THEN
            exp_f := 10;
        ELSIF x =- 10937 THEN
            exp_f := 10;
        ELSIF x =- 10936 THEN
            exp_f := 10;
        ELSIF x =- 10935 THEN
            exp_f := 10;
        ELSIF x =- 10934 THEN
            exp_f := 10;
        ELSIF x =- 10933 THEN
            exp_f := 10;
        ELSIF x =- 10932 THEN
            exp_f := 10;
        ELSIF x =- 10931 THEN
            exp_f := 10;
        ELSIF x =- 10930 THEN
            exp_f := 10;
        ELSIF x =- 10929 THEN
            exp_f := 10;
        ELSIF x =- 10928 THEN
            exp_f := 10;
        ELSIF x =- 10927 THEN
            exp_f := 10;
        ELSIF x =- 10926 THEN
            exp_f := 10;
        ELSIF x =- 10925 THEN
            exp_f := 10;
        ELSIF x =- 10924 THEN
            exp_f := 10;
        ELSIF x =- 10923 THEN
            exp_f := 10;
        ELSIF x =- 10922 THEN
            exp_f := 11;
        ELSIF x =- 10921 THEN
            exp_f := 11;
        ELSIF x =- 10920 THEN
            exp_f := 11;
        ELSIF x =- 10919 THEN
            exp_f := 11;
        ELSIF x =- 10918 THEN
            exp_f := 11;
        ELSIF x =- 10917 THEN
            exp_f := 11;
        ELSIF x =- 10916 THEN
            exp_f := 11;
        ELSIF x =- 10915 THEN
            exp_f := 11;
        ELSIF x =- 10914 THEN
            exp_f := 11;
        ELSIF x =- 10913 THEN
            exp_f := 11;
        ELSIF x =- 10912 THEN
            exp_f := 11;
        ELSIF x =- 10911 THEN
            exp_f := 11;
        ELSIF x =- 10910 THEN
            exp_f := 11;
        ELSIF x =- 10909 THEN
            exp_f := 11;
        ELSIF x =- 10908 THEN
            exp_f := 11;
        ELSIF x =- 10907 THEN
            exp_f := 11;
        ELSIF x =- 10906 THEN
            exp_f := 11;
        ELSIF x =- 10905 THEN
            exp_f := 11;
        ELSIF x =- 10904 THEN
            exp_f := 11;
        ELSIF x =- 10903 THEN
            exp_f := 11;
        ELSIF x =- 10902 THEN
            exp_f := 11;
        ELSIF x =- 10901 THEN
            exp_f := 11;
        ELSIF x =- 10900 THEN
            exp_f := 11;
        ELSIF x =- 10899 THEN
            exp_f := 11;
        ELSIF x =- 10898 THEN
            exp_f := 11;
        ELSIF x =- 10897 THEN
            exp_f := 11;
        ELSIF x =- 10896 THEN
            exp_f := 11;
        ELSIF x =- 10895 THEN
            exp_f := 11;
        ELSIF x =- 10894 THEN
            exp_f := 11;
        ELSIF x =- 10893 THEN
            exp_f := 11;
        ELSIF x =- 10892 THEN
            exp_f := 11;
        ELSIF x =- 10891 THEN
            exp_f := 11;
        ELSIF x =- 10890 THEN
            exp_f := 11;
        ELSIF x =- 10889 THEN
            exp_f := 11;
        ELSIF x =- 10888 THEN
            exp_f := 11;
        ELSIF x =- 10887 THEN
            exp_f := 11;
        ELSIF x =- 10886 THEN
            exp_f := 11;
        ELSIF x =- 10885 THEN
            exp_f := 11;
        ELSIF x =- 10884 THEN
            exp_f := 11;
        ELSIF x =- 10883 THEN
            exp_f := 11;
        ELSIF x =- 10882 THEN
            exp_f := 11;
        ELSIF x =- 10881 THEN
            exp_f := 11;
        ELSIF x =- 10880 THEN
            exp_f := 11;
        ELSIF x =- 10879 THEN
            exp_f := 11;
        ELSIF x =- 10878 THEN
            exp_f := 11;
        ELSIF x =- 10877 THEN
            exp_f := 11;
        ELSIF x =- 10876 THEN
            exp_f := 11;
        ELSIF x =- 10875 THEN
            exp_f := 11;
        ELSIF x =- 10874 THEN
            exp_f := 11;
        ELSIF x =- 10873 THEN
            exp_f := 11;
        ELSIF x =- 10872 THEN
            exp_f := 11;
        ELSIF x =- 10871 THEN
            exp_f := 11;
        ELSIF x =- 10870 THEN
            exp_f := 11;
        ELSIF x =- 10869 THEN
            exp_f := 11;
        ELSIF x =- 10868 THEN
            exp_f := 11;
        ELSIF x =- 10867 THEN
            exp_f := 11;
        ELSIF x =- 10866 THEN
            exp_f := 11;
        ELSIF x =- 10865 THEN
            exp_f := 11;
        ELSIF x =- 10864 THEN
            exp_f := 11;
        ELSIF x =- 10863 THEN
            exp_f := 11;
        ELSIF x =- 10862 THEN
            exp_f := 11;
        ELSIF x =- 10861 THEN
            exp_f := 11;
        ELSIF x =- 10860 THEN
            exp_f := 11;
        ELSIF x =- 10859 THEN
            exp_f := 11;
        ELSIF x =- 10858 THEN
            exp_f := 11;
        ELSIF x =- 10857 THEN
            exp_f := 11;
        ELSIF x =- 10856 THEN
            exp_f := 11;
        ELSIF x =- 10855 THEN
            exp_f := 11;
        ELSIF x =- 10854 THEN
            exp_f := 11;
        ELSIF x =- 10853 THEN
            exp_f := 11;
        ELSIF x =- 10852 THEN
            exp_f := 11;
        ELSIF x =- 10851 THEN
            exp_f := 11;
        ELSIF x =- 10850 THEN
            exp_f := 11;
        ELSIF x =- 10849 THEN
            exp_f := 11;
        ELSIF x =- 10848 THEN
            exp_f := 11;
        ELSIF x =- 10847 THEN
            exp_f := 11;
        ELSIF x =- 10846 THEN
            exp_f := 11;
        ELSIF x =- 10845 THEN
            exp_f := 11;
        ELSIF x =- 10844 THEN
            exp_f := 11;
        ELSIF x =- 10843 THEN
            exp_f := 11;
        ELSIF x =- 10842 THEN
            exp_f := 11;
        ELSIF x =- 10841 THEN
            exp_f := 11;
        ELSIF x =- 10840 THEN
            exp_f := 11;
        ELSIF x =- 10839 THEN
            exp_f := 11;
        ELSIF x =- 10838 THEN
            exp_f := 11;
        ELSIF x =- 10837 THEN
            exp_f := 11;
        ELSIF x =- 10836 THEN
            exp_f := 11;
        ELSIF x =- 10835 THEN
            exp_f := 11;
        ELSIF x =- 10834 THEN
            exp_f := 11;
        ELSIF x =- 10833 THEN
            exp_f := 11;
        ELSIF x =- 10832 THEN
            exp_f := 11;
        ELSIF x =- 10831 THEN
            exp_f := 11;
        ELSIF x =- 10830 THEN
            exp_f := 11;
        ELSIF x =- 10829 THEN
            exp_f := 11;
        ELSIF x =- 10828 THEN
            exp_f := 11;
        ELSIF x =- 10827 THEN
            exp_f := 11;
        ELSIF x =- 10826 THEN
            exp_f := 11;
        ELSIF x =- 10825 THEN
            exp_f := 11;
        ELSIF x =- 10824 THEN
            exp_f := 11;
        ELSIF x =- 10823 THEN
            exp_f := 11;
        ELSIF x =- 10822 THEN
            exp_f := 11;
        ELSIF x =- 10821 THEN
            exp_f := 11;
        ELSIF x =- 10820 THEN
            exp_f := 11;
        ELSIF x =- 10819 THEN
            exp_f := 11;
        ELSIF x =- 10818 THEN
            exp_f := 11;
        ELSIF x =- 10817 THEN
            exp_f := 11;
        ELSIF x =- 10816 THEN
            exp_f := 11;
        ELSIF x =- 10815 THEN
            exp_f := 11;
        ELSIF x =- 10814 THEN
            exp_f := 11;
        ELSIF x =- 10813 THEN
            exp_f := 11;
        ELSIF x =- 10812 THEN
            exp_f := 11;
        ELSIF x =- 10811 THEN
            exp_f := 11;
        ELSIF x =- 10810 THEN
            exp_f := 11;
        ELSIF x =- 10809 THEN
            exp_f := 11;
        ELSIF x =- 10808 THEN
            exp_f := 11;
        ELSIF x =- 10807 THEN
            exp_f := 11;
        ELSIF x =- 10806 THEN
            exp_f := 11;
        ELSIF x =- 10805 THEN
            exp_f := 11;
        ELSIF x =- 10804 THEN
            exp_f := 11;
        ELSIF x =- 10803 THEN
            exp_f := 11;
        ELSIF x =- 10802 THEN
            exp_f := 11;
        ELSIF x =- 10801 THEN
            exp_f := 11;
        ELSIF x =- 10800 THEN
            exp_f := 11;
        ELSIF x =- 10799 THEN
            exp_f := 11;
        ELSIF x =- 10798 THEN
            exp_f := 11;
        ELSIF x =- 10797 THEN
            exp_f := 11;
        ELSIF x =- 10796 THEN
            exp_f := 11;
        ELSIF x =- 10795 THEN
            exp_f := 11;
        ELSIF x =- 10794 THEN
            exp_f := 11;
        ELSIF x =- 10793 THEN
            exp_f := 11;
        ELSIF x =- 10792 THEN
            exp_f := 11;
        ELSIF x =- 10791 THEN
            exp_f := 11;
        ELSIF x =- 10790 THEN
            exp_f := 11;
        ELSIF x =- 10789 THEN
            exp_f := 11;
        ELSIF x =- 10788 THEN
            exp_f := 11;
        ELSIF x =- 10787 THEN
            exp_f := 11;
        ELSIF x =- 10786 THEN
            exp_f := 11;
        ELSIF x =- 10785 THEN
            exp_f := 11;
        ELSIF x =- 10784 THEN
            exp_f := 11;
        ELSIF x =- 10783 THEN
            exp_f := 11;
        ELSIF x =- 10782 THEN
            exp_f := 11;
        ELSIF x =- 10781 THEN
            exp_f := 11;
        ELSIF x =- 10780 THEN
            exp_f := 11;
        ELSIF x =- 10779 THEN
            exp_f := 11;
        ELSIF x =- 10778 THEN
            exp_f := 11;
        ELSIF x =- 10777 THEN
            exp_f := 11;
        ELSIF x =- 10776 THEN
            exp_f := 11;
        ELSIF x =- 10775 THEN
            exp_f := 11;
        ELSIF x =- 10774 THEN
            exp_f := 11;
        ELSIF x =- 10773 THEN
            exp_f := 11;
        ELSIF x =- 10772 THEN
            exp_f := 11;
        ELSIF x =- 10771 THEN
            exp_f := 11;
        ELSIF x =- 10770 THEN
            exp_f := 11;
        ELSIF x =- 10769 THEN
            exp_f := 11;
        ELSIF x =- 10768 THEN
            exp_f := 11;
        ELSIF x =- 10767 THEN
            exp_f := 11;
        ELSIF x =- 10766 THEN
            exp_f := 11;
        ELSIF x =- 10765 THEN
            exp_f := 11;
        ELSIF x =- 10764 THEN
            exp_f := 11;
        ELSIF x =- 10763 THEN
            exp_f := 11;
        ELSIF x =- 10762 THEN
            exp_f := 11;
        ELSIF x =- 10761 THEN
            exp_f := 11;
        ELSIF x =- 10760 THEN
            exp_f := 11;
        ELSIF x =- 10759 THEN
            exp_f := 11;
        ELSIF x =- 10758 THEN
            exp_f := 11;
        ELSIF x =- 10757 THEN
            exp_f := 11;
        ELSIF x =- 10756 THEN
            exp_f := 11;
        ELSIF x =- 10755 THEN
            exp_f := 11;
        ELSIF x =- 10754 THEN
            exp_f := 11;
        ELSIF x =- 10753 THEN
            exp_f := 11;
        ELSIF x =- 10752 THEN
            exp_f := 11;
        ELSIF x =- 10751 THEN
            exp_f := 11;
        ELSIF x =- 10750 THEN
            exp_f := 11;
        ELSIF x =- 10749 THEN
            exp_f := 11;
        ELSIF x =- 10748 THEN
            exp_f := 11;
        ELSIF x =- 10747 THEN
            exp_f := 11;
        ELSIF x =- 10746 THEN
            exp_f := 11;
        ELSIF x =- 10745 THEN
            exp_f := 11;
        ELSIF x =- 10744 THEN
            exp_f := 11;
        ELSIF x =- 10743 THEN
            exp_f := 11;
        ELSIF x =- 10742 THEN
            exp_f := 11;
        ELSIF x =- 10741 THEN
            exp_f := 11;
        ELSIF x =- 10740 THEN
            exp_f := 11;
        ELSIF x =- 10739 THEN
            exp_f := 11;
        ELSIF x =- 10738 THEN
            exp_f := 11;
        ELSIF x =- 10737 THEN
            exp_f := 11;
        ELSIF x =- 10736 THEN
            exp_f := 11;
        ELSIF x =- 10735 THEN
            exp_f := 11;
        ELSIF x =- 10734 THEN
            exp_f := 11;
        ELSIF x =- 10733 THEN
            exp_f := 11;
        ELSIF x =- 10732 THEN
            exp_f := 11;
        ELSIF x =- 10731 THEN
            exp_f := 11;
        ELSIF x =- 10730 THEN
            exp_f := 11;
        ELSIF x =- 10729 THEN
            exp_f := 11;
        ELSIF x =- 10728 THEN
            exp_f := 11;
        ELSIF x =- 10727 THEN
            exp_f := 11;
        ELSIF x =- 10726 THEN
            exp_f := 11;
        ELSIF x =- 10725 THEN
            exp_f := 11;
        ELSIF x =- 10724 THEN
            exp_f := 11;
        ELSIF x =- 10723 THEN
            exp_f := 11;
        ELSIF x =- 10722 THEN
            exp_f := 11;
        ELSIF x =- 10721 THEN
            exp_f := 11;
        ELSIF x =- 10720 THEN
            exp_f := 11;
        ELSIF x =- 10719 THEN
            exp_f := 11;
        ELSIF x =- 10718 THEN
            exp_f := 11;
        ELSIF x =- 10717 THEN
            exp_f := 11;
        ELSIF x =- 10716 THEN
            exp_f := 11;
        ELSIF x =- 10715 THEN
            exp_f := 11;
        ELSIF x =- 10714 THEN
            exp_f := 11;
        ELSIF x =- 10713 THEN
            exp_f := 11;
        ELSIF x =- 10712 THEN
            exp_f := 11;
        ELSIF x =- 10711 THEN
            exp_f := 11;
        ELSIF x =- 10710 THEN
            exp_f := 11;
        ELSIF x =- 10709 THEN
            exp_f := 11;
        ELSIF x =- 10708 THEN
            exp_f := 11;
        ELSIF x =- 10707 THEN
            exp_f := 11;
        ELSIF x =- 10706 THEN
            exp_f := 11;
        ELSIF x =- 10705 THEN
            exp_f := 11;
        ELSIF x =- 10704 THEN
            exp_f := 11;
        ELSIF x =- 10703 THEN
            exp_f := 11;
        ELSIF x =- 10702 THEN
            exp_f := 11;
        ELSIF x =- 10701 THEN
            exp_f := 11;
        ELSIF x =- 10700 THEN
            exp_f := 11;
        ELSIF x =- 10699 THEN
            exp_f := 11;
        ELSIF x =- 10698 THEN
            exp_f := 11;
        ELSIF x =- 10697 THEN
            exp_f := 11;
        ELSIF x =- 10696 THEN
            exp_f := 11;
        ELSIF x =- 10695 THEN
            exp_f := 11;
        ELSIF x =- 10694 THEN
            exp_f := 11;
        ELSIF x =- 10693 THEN
            exp_f := 11;
        ELSIF x =- 10692 THEN
            exp_f := 11;
        ELSIF x =- 10691 THEN
            exp_f := 11;
        ELSIF x =- 10690 THEN
            exp_f := 11;
        ELSIF x =- 10689 THEN
            exp_f := 11;
        ELSIF x =- 10688 THEN
            exp_f := 11;
        ELSIF x =- 10687 THEN
            exp_f := 11;
        ELSIF x =- 10686 THEN
            exp_f := 11;
        ELSIF x =- 10685 THEN
            exp_f := 11;
        ELSIF x =- 10684 THEN
            exp_f := 11;
        ELSIF x =- 10683 THEN
            exp_f := 11;
        ELSIF x =- 10682 THEN
            exp_f := 11;
        ELSIF x =- 10681 THEN
            exp_f := 11;
        ELSIF x =- 10680 THEN
            exp_f := 11;
        ELSIF x =- 10679 THEN
            exp_f := 11;
        ELSIF x =- 10678 THEN
            exp_f := 12;
        ELSIF x =- 10677 THEN
            exp_f := 12;
        ELSIF x =- 10676 THEN
            exp_f := 12;
        ELSIF x =- 10675 THEN
            exp_f := 12;
        ELSIF x =- 10674 THEN
            exp_f := 12;
        ELSIF x =- 10673 THEN
            exp_f := 12;
        ELSIF x =- 10672 THEN
            exp_f := 12;
        ELSIF x =- 10671 THEN
            exp_f := 12;
        ELSIF x =- 10670 THEN
            exp_f := 12;
        ELSIF x =- 10669 THEN
            exp_f := 12;
        ELSIF x =- 10668 THEN
            exp_f := 12;
        ELSIF x =- 10667 THEN
            exp_f := 12;
        ELSIF x =- 10666 THEN
            exp_f := 12;
        ELSIF x =- 10665 THEN
            exp_f := 12;
        ELSIF x =- 10664 THEN
            exp_f := 12;
        ELSIF x =- 10663 THEN
            exp_f := 12;
        ELSIF x =- 10662 THEN
            exp_f := 12;
        ELSIF x =- 10661 THEN
            exp_f := 12;
        ELSIF x =- 10660 THEN
            exp_f := 12;
        ELSIF x =- 10659 THEN
            exp_f := 12;
        ELSIF x =- 10658 THEN
            exp_f := 12;
        ELSIF x =- 10657 THEN
            exp_f := 12;
        ELSIF x =- 10656 THEN
            exp_f := 12;
        ELSIF x =- 10655 THEN
            exp_f := 12;
        ELSIF x =- 10654 THEN
            exp_f := 12;
        ELSIF x =- 10653 THEN
            exp_f := 12;
        ELSIF x =- 10652 THEN
            exp_f := 12;
        ELSIF x =- 10651 THEN
            exp_f := 12;
        ELSIF x =- 10650 THEN
            exp_f := 12;
        ELSIF x =- 10649 THEN
            exp_f := 12;
        ELSIF x =- 10648 THEN
            exp_f := 12;
        ELSIF x =- 10647 THEN
            exp_f := 12;
        ELSIF x =- 10646 THEN
            exp_f := 12;
        ELSIF x =- 10645 THEN
            exp_f := 12;
        ELSIF x =- 10644 THEN
            exp_f := 12;
        ELSIF x =- 10643 THEN
            exp_f := 12;
        ELSIF x =- 10642 THEN
            exp_f := 12;
        ELSIF x =- 10641 THEN
            exp_f := 12;
        ELSIF x =- 10640 THEN
            exp_f := 12;
        ELSIF x =- 10639 THEN
            exp_f := 12;
        ELSIF x =- 10638 THEN
            exp_f := 12;
        ELSIF x =- 10637 THEN
            exp_f := 12;
        ELSIF x =- 10636 THEN
            exp_f := 12;
        ELSIF x =- 10635 THEN
            exp_f := 12;
        ELSIF x =- 10634 THEN
            exp_f := 12;
        ELSIF x =- 10633 THEN
            exp_f := 12;
        ELSIF x =- 10632 THEN
            exp_f := 12;
        ELSIF x =- 10631 THEN
            exp_f := 12;
        ELSIF x =- 10630 THEN
            exp_f := 12;
        ELSIF x =- 10629 THEN
            exp_f := 12;
        ELSIF x =- 10628 THEN
            exp_f := 12;
        ELSIF x =- 10627 THEN
            exp_f := 12;
        ELSIF x =- 10626 THEN
            exp_f := 12;
        ELSIF x =- 10625 THEN
            exp_f := 12;
        ELSIF x =- 10624 THEN
            exp_f := 12;
        ELSIF x =- 10623 THEN
            exp_f := 12;
        ELSIF x =- 10622 THEN
            exp_f := 12;
        ELSIF x =- 10621 THEN
            exp_f := 12;
        ELSIF x =- 10620 THEN
            exp_f := 12;
        ELSIF x =- 10619 THEN
            exp_f := 12;
        ELSIF x =- 10618 THEN
            exp_f := 12;
        ELSIF x =- 10617 THEN
            exp_f := 12;
        ELSIF x =- 10616 THEN
            exp_f := 12;
        ELSIF x =- 10615 THEN
            exp_f := 12;
        ELSIF x =- 10614 THEN
            exp_f := 12;
        ELSIF x =- 10613 THEN
            exp_f := 12;
        ELSIF x =- 10612 THEN
            exp_f := 12;
        ELSIF x =- 10611 THEN
            exp_f := 12;
        ELSIF x =- 10610 THEN
            exp_f := 12;
        ELSIF x =- 10609 THEN
            exp_f := 12;
        ELSIF x =- 10608 THEN
            exp_f := 12;
        ELSIF x =- 10607 THEN
            exp_f := 12;
        ELSIF x =- 10606 THEN
            exp_f := 12;
        ELSIF x =- 10605 THEN
            exp_f := 12;
        ELSIF x =- 10604 THEN
            exp_f := 12;
        ELSIF x =- 10603 THEN
            exp_f := 12;
        ELSIF x =- 10602 THEN
            exp_f := 12;
        ELSIF x =- 10601 THEN
            exp_f := 12;
        ELSIF x =- 10600 THEN
            exp_f := 12;
        ELSIF x =- 10599 THEN
            exp_f := 12;
        ELSIF x =- 10598 THEN
            exp_f := 12;
        ELSIF x =- 10597 THEN
            exp_f := 12;
        ELSIF x =- 10596 THEN
            exp_f := 12;
        ELSIF x =- 10595 THEN
            exp_f := 12;
        ELSIF x =- 10594 THEN
            exp_f := 12;
        ELSIF x =- 10593 THEN
            exp_f := 12;
        ELSIF x =- 10592 THEN
            exp_f := 12;
        ELSIF x =- 10591 THEN
            exp_f := 12;
        ELSIF x =- 10590 THEN
            exp_f := 12;
        ELSIF x =- 10589 THEN
            exp_f := 12;
        ELSIF x =- 10588 THEN
            exp_f := 12;
        ELSIF x =- 10587 THEN
            exp_f := 12;
        ELSIF x =- 10586 THEN
            exp_f := 12;
        ELSIF x =- 10585 THEN
            exp_f := 12;
        ELSIF x =- 10584 THEN
            exp_f := 12;
        ELSIF x =- 10583 THEN
            exp_f := 12;
        ELSIF x =- 10582 THEN
            exp_f := 12;
        ELSIF x =- 10581 THEN
            exp_f := 12;
        ELSIF x =- 10580 THEN
            exp_f := 12;
        ELSIF x =- 10579 THEN
            exp_f := 12;
        ELSIF x =- 10578 THEN
            exp_f := 12;
        ELSIF x =- 10577 THEN
            exp_f := 12;
        ELSIF x =- 10576 THEN
            exp_f := 12;
        ELSIF x =- 10575 THEN
            exp_f := 12;
        ELSIF x =- 10574 THEN
            exp_f := 12;
        ELSIF x =- 10573 THEN
            exp_f := 12;
        ELSIF x =- 10572 THEN
            exp_f := 12;
        ELSIF x =- 10571 THEN
            exp_f := 12;
        ELSIF x =- 10570 THEN
            exp_f := 12;
        ELSIF x =- 10569 THEN
            exp_f := 12;
        ELSIF x =- 10568 THEN
            exp_f := 12;
        ELSIF x =- 10567 THEN
            exp_f := 12;
        ELSIF x =- 10566 THEN
            exp_f := 12;
        ELSIF x =- 10565 THEN
            exp_f := 12;
        ELSIF x =- 10564 THEN
            exp_f := 12;
        ELSIF x =- 10563 THEN
            exp_f := 12;
        ELSIF x =- 10562 THEN
            exp_f := 12;
        ELSIF x =- 10561 THEN
            exp_f := 12;
        ELSIF x =- 10560 THEN
            exp_f := 12;
        ELSIF x =- 10559 THEN
            exp_f := 12;
        ELSIF x =- 10558 THEN
            exp_f := 12;
        ELSIF x =- 10557 THEN
            exp_f := 12;
        ELSIF x =- 10556 THEN
            exp_f := 12;
        ELSIF x =- 10555 THEN
            exp_f := 12;
        ELSIF x =- 10554 THEN
            exp_f := 12;
        ELSIF x =- 10553 THEN
            exp_f := 12;
        ELSIF x =- 10552 THEN
            exp_f := 12;
        ELSIF x =- 10551 THEN
            exp_f := 12;
        ELSIF x =- 10550 THEN
            exp_f := 12;
        ELSIF x =- 10549 THEN
            exp_f := 12;
        ELSIF x =- 10548 THEN
            exp_f := 12;
        ELSIF x =- 10547 THEN
            exp_f := 12;
        ELSIF x =- 10546 THEN
            exp_f := 12;
        ELSIF x =- 10545 THEN
            exp_f := 12;
        ELSIF x =- 10544 THEN
            exp_f := 12;
        ELSIF x =- 10543 THEN
            exp_f := 12;
        ELSIF x =- 10542 THEN
            exp_f := 12;
        ELSIF x =- 10541 THEN
            exp_f := 12;
        ELSIF x =- 10540 THEN
            exp_f := 12;
        ELSIF x =- 10539 THEN
            exp_f := 12;
        ELSIF x =- 10538 THEN
            exp_f := 12;
        ELSIF x =- 10537 THEN
            exp_f := 12;
        ELSIF x =- 10536 THEN
            exp_f := 12;
        ELSIF x =- 10535 THEN
            exp_f := 12;
        ELSIF x =- 10534 THEN
            exp_f := 12;
        ELSIF x =- 10533 THEN
            exp_f := 12;
        ELSIF x =- 10532 THEN
            exp_f := 13;
        ELSIF x =- 10531 THEN
            exp_f := 13;
        ELSIF x =- 10530 THEN
            exp_f := 13;
        ELSIF x =- 10529 THEN
            exp_f := 13;
        ELSIF x =- 10528 THEN
            exp_f := 13;
        ELSIF x =- 10527 THEN
            exp_f := 13;
        ELSIF x =- 10526 THEN
            exp_f := 13;
        ELSIF x =- 10525 THEN
            exp_f := 13;
        ELSIF x =- 10524 THEN
            exp_f := 13;
        ELSIF x =- 10523 THEN
            exp_f := 13;
        ELSIF x =- 10522 THEN
            exp_f := 13;
        ELSIF x =- 10521 THEN
            exp_f := 13;
        ELSIF x =- 10520 THEN
            exp_f := 13;
        ELSIF x =- 10519 THEN
            exp_f := 13;
        ELSIF x =- 10518 THEN
            exp_f := 13;
        ELSIF x =- 10517 THEN
            exp_f := 13;
        ELSIF x =- 10516 THEN
            exp_f := 13;
        ELSIF x =- 10515 THEN
            exp_f := 13;
        ELSIF x =- 10514 THEN
            exp_f := 13;
        ELSIF x =- 10513 THEN
            exp_f := 13;
        ELSIF x =- 10512 THEN
            exp_f := 13;
        ELSIF x =- 10511 THEN
            exp_f := 13;
        ELSIF x =- 10510 THEN
            exp_f := 13;
        ELSIF x =- 10509 THEN
            exp_f := 13;
        ELSIF x =- 10508 THEN
            exp_f := 13;
        ELSIF x =- 10507 THEN
            exp_f := 13;
        ELSIF x =- 10506 THEN
            exp_f := 13;
        ELSIF x =- 10505 THEN
            exp_f := 13;
        ELSIF x =- 10504 THEN
            exp_f := 13;
        ELSIF x =- 10503 THEN
            exp_f := 13;
        ELSIF x =- 10502 THEN
            exp_f := 13;
        ELSIF x =- 10501 THEN
            exp_f := 13;
        ELSIF x =- 10500 THEN
            exp_f := 13;
        ELSIF x =- 10499 THEN
            exp_f := 13;
        ELSIF x =- 10498 THEN
            exp_f := 13;
        ELSIF x =- 10497 THEN
            exp_f := 13;
        ELSIF x =- 10496 THEN
            exp_f := 13;
        ELSIF x =- 10495 THEN
            exp_f := 13;
        ELSIF x =- 10494 THEN
            exp_f := 13;
        ELSIF x =- 10493 THEN
            exp_f := 13;
        ELSIF x =- 10492 THEN
            exp_f := 13;
        ELSIF x =- 10491 THEN
            exp_f := 13;
        ELSIF x =- 10490 THEN
            exp_f := 13;
        ELSIF x =- 10489 THEN
            exp_f := 13;
        ELSIF x =- 10488 THEN
            exp_f := 13;
        ELSIF x =- 10487 THEN
            exp_f := 13;
        ELSIF x =- 10486 THEN
            exp_f := 13;
        ELSIF x =- 10485 THEN
            exp_f := 13;
        ELSIF x =- 10484 THEN
            exp_f := 13;
        ELSIF x =- 10483 THEN
            exp_f := 13;
        ELSIF x =- 10482 THEN
            exp_f := 13;
        ELSIF x =- 10481 THEN
            exp_f := 13;
        ELSIF x =- 10480 THEN
            exp_f := 13;
        ELSIF x =- 10479 THEN
            exp_f := 13;
        ELSIF x =- 10478 THEN
            exp_f := 13;
        ELSIF x =- 10477 THEN
            exp_f := 13;
        ELSIF x =- 10476 THEN
            exp_f := 13;
        ELSIF x =- 10475 THEN
            exp_f := 13;
        ELSIF x =- 10474 THEN
            exp_f := 13;
        ELSIF x =- 10473 THEN
            exp_f := 13;
        ELSIF x =- 10472 THEN
            exp_f := 13;
        ELSIF x =- 10471 THEN
            exp_f := 13;
        ELSIF x =- 10470 THEN
            exp_f := 13;
        ELSIF x =- 10469 THEN
            exp_f := 13;
        ELSIF x =- 10468 THEN
            exp_f := 13;
        ELSIF x =- 10467 THEN
            exp_f := 13;
        ELSIF x =- 10466 THEN
            exp_f := 13;
        ELSIF x =- 10465 THEN
            exp_f := 13;
        ELSIF x =- 10464 THEN
            exp_f := 13;
        ELSIF x =- 10463 THEN
            exp_f := 13;
        ELSIF x =- 10462 THEN
            exp_f := 13;
        ELSIF x =- 10461 THEN
            exp_f := 13;
        ELSIF x =- 10460 THEN
            exp_f := 13;
        ELSIF x =- 10459 THEN
            exp_f := 13;
        ELSIF x =- 10458 THEN
            exp_f := 13;
        ELSIF x =- 10457 THEN
            exp_f := 13;
        ELSIF x =- 10456 THEN
            exp_f := 13;
        ELSIF x =- 10455 THEN
            exp_f := 13;
        ELSIF x =- 10454 THEN
            exp_f := 13;
        ELSIF x =- 10453 THEN
            exp_f := 13;
        ELSIF x =- 10452 THEN
            exp_f := 13;
        ELSIF x =- 10451 THEN
            exp_f := 13;
        ELSIF x =- 10450 THEN
            exp_f := 13;
        ELSIF x =- 10449 THEN
            exp_f := 13;
        ELSIF x =- 10448 THEN
            exp_f := 13;
        ELSIF x =- 10447 THEN
            exp_f := 13;
        ELSIF x =- 10446 THEN
            exp_f := 13;
        ELSIF x =- 10445 THEN
            exp_f := 13;
        ELSIF x =- 10444 THEN
            exp_f := 13;
        ELSIF x =- 10443 THEN
            exp_f := 13;
        ELSIF x =- 10442 THEN
            exp_f := 13;
        ELSIF x =- 10441 THEN
            exp_f := 13;
        ELSIF x =- 10440 THEN
            exp_f := 13;
        ELSIF x =- 10439 THEN
            exp_f := 13;
        ELSIF x =- 10438 THEN
            exp_f := 13;
        ELSIF x =- 10437 THEN
            exp_f := 13;
        ELSIF x =- 10436 THEN
            exp_f := 13;
        ELSIF x =- 10435 THEN
            exp_f := 13;
        ELSIF x =- 10434 THEN
            exp_f := 13;
        ELSIF x =- 10433 THEN
            exp_f := 13;
        ELSIF x =- 10432 THEN
            exp_f := 13;
        ELSIF x =- 10431 THEN
            exp_f := 13;
        ELSIF x =- 10430 THEN
            exp_f := 13;
        ELSIF x =- 10429 THEN
            exp_f := 13;
        ELSIF x =- 10428 THEN
            exp_f := 13;
        ELSIF x =- 10427 THEN
            exp_f := 13;
        ELSIF x =- 10426 THEN
            exp_f := 13;
        ELSIF x =- 10425 THEN
            exp_f := 13;
        ELSIF x =- 10424 THEN
            exp_f := 13;
        ELSIF x =- 10423 THEN
            exp_f := 13;
        ELSIF x =- 10422 THEN
            exp_f := 13;
        ELSIF x =- 10421 THEN
            exp_f := 13;
        ELSIF x =- 10420 THEN
            exp_f := 13;
        ELSIF x =- 10419 THEN
            exp_f := 13;
        ELSIF x =- 10418 THEN
            exp_f := 13;
        ELSIF x =- 10417 THEN
            exp_f := 13;
        ELSIF x =- 10416 THEN
            exp_f := 13;
        ELSIF x =- 10415 THEN
            exp_f := 13;
        ELSIF x =- 10414 THEN
            exp_f := 13;
        ELSIF x =- 10413 THEN
            exp_f := 13;
        ELSIF x =- 10412 THEN
            exp_f := 13;
        ELSIF x =- 10411 THEN
            exp_f := 13;
        ELSIF x =- 10410 THEN
            exp_f := 13;
        ELSIF x =- 10409 THEN
            exp_f := 13;
        ELSIF x =- 10408 THEN
            exp_f := 13;
        ELSIF x =- 10407 THEN
            exp_f := 13;
        ELSIF x =- 10406 THEN
            exp_f := 13;
        ELSIF x =- 10405 THEN
            exp_f := 13;
        ELSIF x =- 10404 THEN
            exp_f := 13;
        ELSIF x =- 10403 THEN
            exp_f := 13;
        ELSIF x =- 10402 THEN
            exp_f := 13;
        ELSIF x =- 10401 THEN
            exp_f := 13;
        ELSIF x =- 10400 THEN
            exp_f := 13;
        ELSIF x =- 10399 THEN
            exp_f := 13;
        ELSIF x =- 10398 THEN
            exp_f := 13;
        ELSIF x =- 10397 THEN
            exp_f := 13;
        ELSIF x =- 10396 THEN
            exp_f := 13;
        ELSIF x =- 10395 THEN
            exp_f := 13;
        ELSIF x =- 10394 THEN
            exp_f := 13;
        ELSIF x =- 10393 THEN
            exp_f := 13;
        ELSIF x =- 10392 THEN
            exp_f := 13;
        ELSIF x =- 10391 THEN
            exp_f := 13;
        ELSIF x =- 10390 THEN
            exp_f := 13;
        ELSIF x =- 10389 THEN
            exp_f := 13;
        ELSIF x =- 10388 THEN
            exp_f := 13;
        ELSIF x =- 10387 THEN
            exp_f := 13;
        ELSIF x =- 10386 THEN
            exp_f := 14;
        ELSIF x =- 10385 THEN
            exp_f := 14;
        ELSIF x =- 10384 THEN
            exp_f := 14;
        ELSIF x =- 10383 THEN
            exp_f := 14;
        ELSIF x =- 10382 THEN
            exp_f := 14;
        ELSIF x =- 10381 THEN
            exp_f := 14;
        ELSIF x =- 10380 THEN
            exp_f := 14;
        ELSIF x =- 10379 THEN
            exp_f := 14;
        ELSIF x =- 10378 THEN
            exp_f := 14;
        ELSIF x =- 10377 THEN
            exp_f := 14;
        ELSIF x =- 10376 THEN
            exp_f := 14;
        ELSIF x =- 10375 THEN
            exp_f := 14;
        ELSIF x =- 10374 THEN
            exp_f := 14;
        ELSIF x =- 10373 THEN
            exp_f := 14;
        ELSIF x =- 10372 THEN
            exp_f := 14;
        ELSIF x =- 10371 THEN
            exp_f := 14;
        ELSIF x =- 10370 THEN
            exp_f := 14;
        ELSIF x =- 10369 THEN
            exp_f := 14;
        ELSIF x =- 10368 THEN
            exp_f := 14;
        ELSIF x =- 10367 THEN
            exp_f := 14;
        ELSIF x =- 10366 THEN
            exp_f := 14;
        ELSIF x =- 10365 THEN
            exp_f := 14;
        ELSIF x =- 10364 THEN
            exp_f := 14;
        ELSIF x =- 10363 THEN
            exp_f := 14;
        ELSIF x =- 10362 THEN
            exp_f := 14;
        ELSIF x =- 10361 THEN
            exp_f := 14;
        ELSIF x =- 10360 THEN
            exp_f := 14;
        ELSIF x =- 10359 THEN
            exp_f := 14;
        ELSIF x =- 10358 THEN
            exp_f := 14;
        ELSIF x =- 10357 THEN
            exp_f := 14;
        ELSIF x =- 10356 THEN
            exp_f := 14;
        ELSIF x =- 10355 THEN
            exp_f := 14;
        ELSIF x =- 10354 THEN
            exp_f := 14;
        ELSIF x =- 10353 THEN
            exp_f := 14;
        ELSIF x =- 10352 THEN
            exp_f := 14;
        ELSIF x =- 10351 THEN
            exp_f := 14;
        ELSIF x =- 10350 THEN
            exp_f := 14;
        ELSIF x =- 10349 THEN
            exp_f := 14;
        ELSIF x =- 10348 THEN
            exp_f := 14;
        ELSIF x =- 10347 THEN
            exp_f := 14;
        ELSIF x =- 10346 THEN
            exp_f := 14;
        ELSIF x =- 10345 THEN
            exp_f := 14;
        ELSIF x =- 10344 THEN
            exp_f := 14;
        ELSIF x =- 10343 THEN
            exp_f := 14;
        ELSIF x =- 10342 THEN
            exp_f := 14;
        ELSIF x =- 10341 THEN
            exp_f := 14;
        ELSIF x =- 10340 THEN
            exp_f := 14;
        ELSIF x =- 10339 THEN
            exp_f := 14;
        ELSIF x =- 10338 THEN
            exp_f := 14;
        ELSIF x =- 10337 THEN
            exp_f := 14;
        ELSIF x =- 10336 THEN
            exp_f := 14;
        ELSIF x =- 10335 THEN
            exp_f := 14;
        ELSIF x =- 10334 THEN
            exp_f := 14;
        ELSIF x =- 10333 THEN
            exp_f := 14;
        ELSIF x =- 10332 THEN
            exp_f := 14;
        ELSIF x =- 10331 THEN
            exp_f := 14;
        ELSIF x =- 10330 THEN
            exp_f := 14;
        ELSIF x =- 10329 THEN
            exp_f := 14;
        ELSIF x =- 10328 THEN
            exp_f := 14;
        ELSIF x =- 10327 THEN
            exp_f := 14;
        ELSIF x =- 10326 THEN
            exp_f := 14;
        ELSIF x =- 10325 THEN
            exp_f := 14;
        ELSIF x =- 10324 THEN
            exp_f := 14;
        ELSIF x =- 10323 THEN
            exp_f := 14;
        ELSIF x =- 10322 THEN
            exp_f := 14;
        ELSIF x =- 10321 THEN
            exp_f := 14;
        ELSIF x =- 10320 THEN
            exp_f := 14;
        ELSIF x =- 10319 THEN
            exp_f := 14;
        ELSIF x =- 10318 THEN
            exp_f := 14;
        ELSIF x =- 10317 THEN
            exp_f := 14;
        ELSIF x =- 10316 THEN
            exp_f := 14;
        ELSIF x =- 10315 THEN
            exp_f := 14;
        ELSIF x =- 10314 THEN
            exp_f := 14;
        ELSIF x =- 10313 THEN
            exp_f := 14;
        ELSIF x =- 10312 THEN
            exp_f := 14;
        ELSIF x =- 10311 THEN
            exp_f := 14;
        ELSIF x =- 10310 THEN
            exp_f := 14;
        ELSIF x =- 10309 THEN
            exp_f := 14;
        ELSIF x =- 10308 THEN
            exp_f := 14;
        ELSIF x =- 10307 THEN
            exp_f := 14;
        ELSIF x =- 10306 THEN
            exp_f := 14;
        ELSIF x =- 10305 THEN
            exp_f := 14;
        ELSIF x =- 10304 THEN
            exp_f := 14;
        ELSIF x =- 10303 THEN
            exp_f := 14;
        ELSIF x =- 10302 THEN
            exp_f := 14;
        ELSIF x =- 10301 THEN
            exp_f := 14;
        ELSIF x =- 10300 THEN
            exp_f := 14;
        ELSIF x =- 10299 THEN
            exp_f := 14;
        ELSIF x =- 10298 THEN
            exp_f := 14;
        ELSIF x =- 10297 THEN
            exp_f := 14;
        ELSIF x =- 10296 THEN
            exp_f := 14;
        ELSIF x =- 10295 THEN
            exp_f := 14;
        ELSIF x =- 10294 THEN
            exp_f := 14;
        ELSIF x =- 10293 THEN
            exp_f := 14;
        ELSIF x =- 10292 THEN
            exp_f := 14;
        ELSIF x =- 10291 THEN
            exp_f := 14;
        ELSIF x =- 10290 THEN
            exp_f := 14;
        ELSIF x =- 10289 THEN
            exp_f := 14;
        ELSIF x =- 10288 THEN
            exp_f := 14;
        ELSIF x =- 10287 THEN
            exp_f := 14;
        ELSIF x =- 10286 THEN
            exp_f := 14;
        ELSIF x =- 10285 THEN
            exp_f := 14;
        ELSIF x =- 10284 THEN
            exp_f := 14;
        ELSIF x =- 10283 THEN
            exp_f := 14;
        ELSIF x =- 10282 THEN
            exp_f := 14;
        ELSIF x =- 10281 THEN
            exp_f := 14;
        ELSIF x =- 10280 THEN
            exp_f := 14;
        ELSIF x =- 10279 THEN
            exp_f := 14;
        ELSIF x =- 10278 THEN
            exp_f := 14;
        ELSIF x =- 10277 THEN
            exp_f := 14;
        ELSIF x =- 10276 THEN
            exp_f := 14;
        ELSIF x =- 10275 THEN
            exp_f := 14;
        ELSIF x =- 10274 THEN
            exp_f := 14;
        ELSIF x =- 10273 THEN
            exp_f := 14;
        ELSIF x =- 10272 THEN
            exp_f := 14;
        ELSIF x =- 10271 THEN
            exp_f := 14;
        ELSIF x =- 10270 THEN
            exp_f := 14;
        ELSIF x =- 10269 THEN
            exp_f := 14;
        ELSIF x =- 10268 THEN
            exp_f := 14;
        ELSIF x =- 10267 THEN
            exp_f := 14;
        ELSIF x =- 10266 THEN
            exp_f := 14;
        ELSIF x =- 10265 THEN
            exp_f := 14;
        ELSIF x =- 10264 THEN
            exp_f := 14;
        ELSIF x =- 10263 THEN
            exp_f := 14;
        ELSIF x =- 10262 THEN
            exp_f := 14;
        ELSIF x =- 10261 THEN
            exp_f := 14;
        ELSIF x =- 10260 THEN
            exp_f := 14;
        ELSIF x =- 10259 THEN
            exp_f := 14;
        ELSIF x =- 10258 THEN
            exp_f := 14;
        ELSIF x =- 10257 THEN
            exp_f := 14;
        ELSIF x =- 10256 THEN
            exp_f := 14;
        ELSIF x =- 10255 THEN
            exp_f := 14;
        ELSIF x =- 10254 THEN
            exp_f := 14;
        ELSIF x =- 10253 THEN
            exp_f := 14;
        ELSIF x =- 10252 THEN
            exp_f := 14;
        ELSIF x =- 10251 THEN
            exp_f := 14;
        ELSIF x =- 10250 THEN
            exp_f := 14;
        ELSIF x =- 10249 THEN
            exp_f := 14;
        ELSIF x =- 10248 THEN
            exp_f := 14;
        ELSIF x =- 10247 THEN
            exp_f := 14;
        ELSIF x =- 10246 THEN
            exp_f := 14;
        ELSIF x =- 10245 THEN
            exp_f := 14;
        ELSIF x =- 10244 THEN
            exp_f := 14;
        ELSIF x =- 10243 THEN
            exp_f := 14;
        ELSIF x =- 10242 THEN
            exp_f := 14;
        ELSIF x =- 10241 THEN
            exp_f := 14;
        ELSIF x =- 10240 THEN
            exp_f := 14;
        ELSIF x =- 10239 THEN
            exp_f := 15;
        ELSIF x =- 10238 THEN
            exp_f := 15;
        ELSIF x =- 10237 THEN
            exp_f := 15;
        ELSIF x =- 10236 THEN
            exp_f := 15;
        ELSIF x =- 10235 THEN
            exp_f := 15;
        ELSIF x =- 10234 THEN
            exp_f := 15;
        ELSIF x =- 10233 THEN
            exp_f := 15;
        ELSIF x =- 10232 THEN
            exp_f := 15;
        ELSIF x =- 10231 THEN
            exp_f := 15;
        ELSIF x =- 10230 THEN
            exp_f := 15;
        ELSIF x =- 10229 THEN
            exp_f := 15;
        ELSIF x =- 10228 THEN
            exp_f := 15;
        ELSIF x =- 10227 THEN
            exp_f := 15;
        ELSIF x =- 10226 THEN
            exp_f := 15;
        ELSIF x =- 10225 THEN
            exp_f := 15;
        ELSIF x =- 10224 THEN
            exp_f := 15;
        ELSIF x =- 10223 THEN
            exp_f := 15;
        ELSIF x =- 10222 THEN
            exp_f := 15;
        ELSIF x =- 10221 THEN
            exp_f := 15;
        ELSIF x =- 10220 THEN
            exp_f := 15;
        ELSIF x =- 10219 THEN
            exp_f := 15;
        ELSIF x =- 10218 THEN
            exp_f := 15;
        ELSIF x =- 10217 THEN
            exp_f := 15;
        ELSIF x =- 10216 THEN
            exp_f := 15;
        ELSIF x =- 10215 THEN
            exp_f := 15;
        ELSIF x =- 10214 THEN
            exp_f := 15;
        ELSIF x =- 10213 THEN
            exp_f := 15;
        ELSIF x =- 10212 THEN
            exp_f := 15;
        ELSIF x =- 10211 THEN
            exp_f := 15;
        ELSIF x =- 10210 THEN
            exp_f := 15;
        ELSIF x =- 10209 THEN
            exp_f := 15;
        ELSIF x =- 10208 THEN
            exp_f := 15;
        ELSIF x =- 10207 THEN
            exp_f := 15;
        ELSIF x =- 10206 THEN
            exp_f := 15;
        ELSIF x =- 10205 THEN
            exp_f := 15;
        ELSIF x =- 10204 THEN
            exp_f := 15;
        ELSIF x =- 10203 THEN
            exp_f := 15;
        ELSIF x =- 10202 THEN
            exp_f := 15;
        ELSIF x =- 10201 THEN
            exp_f := 15;
        ELSIF x =- 10200 THEN
            exp_f := 15;
        ELSIF x =- 10199 THEN
            exp_f := 15;
        ELSIF x =- 10198 THEN
            exp_f := 15;
        ELSIF x =- 10197 THEN
            exp_f := 15;
        ELSIF x =- 10196 THEN
            exp_f := 15;
        ELSIF x =- 10195 THEN
            exp_f := 15;
        ELSIF x =- 10194 THEN
            exp_f := 15;
        ELSIF x =- 10193 THEN
            exp_f := 15;
        ELSIF x =- 10192 THEN
            exp_f := 15;
        ELSIF x =- 10191 THEN
            exp_f := 15;
        ELSIF x =- 10190 THEN
            exp_f := 15;
        ELSIF x =- 10189 THEN
            exp_f := 15;
        ELSIF x =- 10188 THEN
            exp_f := 15;
        ELSIF x =- 10187 THEN
            exp_f := 15;
        ELSIF x =- 10186 THEN
            exp_f := 15;
        ELSIF x =- 10185 THEN
            exp_f := 15;
        ELSIF x =- 10184 THEN
            exp_f := 15;
        ELSIF x =- 10183 THEN
            exp_f := 15;
        ELSIF x =- 10182 THEN
            exp_f := 15;
        ELSIF x =- 10181 THEN
            exp_f := 15;
        ELSIF x =- 10180 THEN
            exp_f := 15;
        ELSIF x =- 10179 THEN
            exp_f := 15;
        ELSIF x =- 10178 THEN
            exp_f := 15;
        ELSIF x =- 10177 THEN
            exp_f := 15;
        ELSIF x =- 10176 THEN
            exp_f := 15;
        ELSIF x =- 10175 THEN
            exp_f := 15;
        ELSIF x =- 10174 THEN
            exp_f := 15;
        ELSIF x =- 10173 THEN
            exp_f := 15;
        ELSIF x =- 10172 THEN
            exp_f := 15;
        ELSIF x =- 10171 THEN
            exp_f := 15;
        ELSIF x =- 10170 THEN
            exp_f := 15;
        ELSIF x =- 10169 THEN
            exp_f := 15;
        ELSIF x =- 10168 THEN
            exp_f := 15;
        ELSIF x =- 10167 THEN
            exp_f := 15;
        ELSIF x =- 10166 THEN
            exp_f := 15;
        ELSIF x =- 10165 THEN
            exp_f := 15;
        ELSIF x =- 10164 THEN
            exp_f := 15;
        ELSIF x =- 10163 THEN
            exp_f := 15;
        ELSIF x =- 10162 THEN
            exp_f := 15;
        ELSIF x =- 10161 THEN
            exp_f := 15;
        ELSIF x =- 10160 THEN
            exp_f := 15;
        ELSIF x =- 10159 THEN
            exp_f := 15;
        ELSIF x =- 10158 THEN
            exp_f := 15;
        ELSIF x =- 10157 THEN
            exp_f := 15;
        ELSIF x =- 10156 THEN
            exp_f := 15;
        ELSIF x =- 10155 THEN
            exp_f := 15;
        ELSIF x =- 10154 THEN
            exp_f := 15;
        ELSIF x =- 10153 THEN
            exp_f := 15;
        ELSIF x =- 10152 THEN
            exp_f := 15;
        ELSIF x =- 10151 THEN
            exp_f := 15;
        ELSIF x =- 10150 THEN
            exp_f := 15;
        ELSIF x =- 10149 THEN
            exp_f := 15;
        ELSIF x =- 10148 THEN
            exp_f := 15;
        ELSIF x =- 10147 THEN
            exp_f := 15;
        ELSIF x =- 10146 THEN
            exp_f := 15;
        ELSIF x =- 10145 THEN
            exp_f := 15;
        ELSIF x =- 10144 THEN
            exp_f := 15;
        ELSIF x =- 10143 THEN
            exp_f := 15;
        ELSIF x =- 10142 THEN
            exp_f := 15;
        ELSIF x =- 10141 THEN
            exp_f := 15;
        ELSIF x =- 10140 THEN
            exp_f := 15;
        ELSIF x =- 10139 THEN
            exp_f := 15;
        ELSIF x =- 10138 THEN
            exp_f := 15;
        ELSIF x =- 10137 THEN
            exp_f := 15;
        ELSIF x =- 10136 THEN
            exp_f := 15;
        ELSIF x =- 10135 THEN
            exp_f := 15;
        ELSIF x =- 10134 THEN
            exp_f := 15;
        ELSIF x =- 10133 THEN
            exp_f := 15;
        ELSIF x =- 10132 THEN
            exp_f := 15;
        ELSIF x =- 10131 THEN
            exp_f := 15;
        ELSIF x =- 10130 THEN
            exp_f := 15;
        ELSIF x =- 10129 THEN
            exp_f := 15;
        ELSIF x =- 10128 THEN
            exp_f := 15;
        ELSIF x =- 10127 THEN
            exp_f := 15;
        ELSIF x =- 10126 THEN
            exp_f := 15;
        ELSIF x =- 10125 THEN
            exp_f := 15;
        ELSIF x =- 10124 THEN
            exp_f := 15;
        ELSIF x =- 10123 THEN
            exp_f := 15;
        ELSIF x =- 10122 THEN
            exp_f := 15;
        ELSIF x =- 10121 THEN
            exp_f := 15;
        ELSIF x =- 10120 THEN
            exp_f := 15;
        ELSIF x =- 10119 THEN
            exp_f := 15;
        ELSIF x =- 10118 THEN
            exp_f := 15;
        ELSIF x =- 10117 THEN
            exp_f := 15;
        ELSIF x =- 10116 THEN
            exp_f := 15;
        ELSIF x =- 10115 THEN
            exp_f := 15;
        ELSIF x =- 10114 THEN
            exp_f := 15;
        ELSIF x =- 10113 THEN
            exp_f := 15;
        ELSIF x =- 10112 THEN
            exp_f := 15;
        ELSIF x =- 10111 THEN
            exp_f := 15;
        ELSIF x =- 10110 THEN
            exp_f := 15;
        ELSIF x =- 10109 THEN
            exp_f := 15;
        ELSIF x =- 10108 THEN
            exp_f := 15;
        ELSIF x =- 10107 THEN
            exp_f := 15;
        ELSIF x =- 10106 THEN
            exp_f := 15;
        ELSIF x =- 10105 THEN
            exp_f := 15;
        ELSIF x =- 10104 THEN
            exp_f := 15;
        ELSIF x =- 10103 THEN
            exp_f := 15;
        ELSIF x =- 10102 THEN
            exp_f := 15;
        ELSIF x =- 10101 THEN
            exp_f := 15;
        ELSIF x =- 10100 THEN
            exp_f := 15;
        ELSIF x =- 10099 THEN
            exp_f := 15;
        ELSIF x =- 10098 THEN
            exp_f := 15;
        ELSIF x =- 10097 THEN
            exp_f := 15;
        ELSIF x =- 10096 THEN
            exp_f := 15;
        ELSIF x =- 10095 THEN
            exp_f := 15;
        ELSIF x =- 10094 THEN
            exp_f := 15;
        ELSIF x =- 10093 THEN
            exp_f := 15;
        ELSIF x =- 10092 THEN
            exp_f := 15;
        ELSIF x =- 10091 THEN
            exp_f := 15;
        ELSIF x =- 10090 THEN
            exp_f := 15;
        ELSIF x =- 10089 THEN
            exp_f := 15;
        ELSIF x =- 10088 THEN
            exp_f := 15;
        ELSIF x =- 10087 THEN
            exp_f := 15;
        ELSIF x =- 10086 THEN
            exp_f := 15;
        ELSIF x =- 10085 THEN
            exp_f := 15;
        ELSIF x =- 10084 THEN
            exp_f := 15;
        ELSIF x =- 10083 THEN
            exp_f := 15;
        ELSIF x =- 10082 THEN
            exp_f := 16;
        ELSIF x =- 10081 THEN
            exp_f := 16;
        ELSIF x =- 10080 THEN
            exp_f := 16;
        ELSIF x =- 10079 THEN
            exp_f := 16;
        ELSIF x =- 10078 THEN
            exp_f := 16;
        ELSIF x =- 10077 THEN
            exp_f := 16;
        ELSIF x =- 10076 THEN
            exp_f := 16;
        ELSIF x =- 10075 THEN
            exp_f := 16;
        ELSIF x =- 10074 THEN
            exp_f := 16;
        ELSIF x =- 10073 THEN
            exp_f := 16;
        ELSIF x =- 10072 THEN
            exp_f := 16;
        ELSIF x =- 10071 THEN
            exp_f := 16;
        ELSIF x =- 10070 THEN
            exp_f := 16;
        ELSIF x =- 10069 THEN
            exp_f := 16;
        ELSIF x =- 10068 THEN
            exp_f := 16;
        ELSIF x =- 10067 THEN
            exp_f := 16;
        ELSIF x =- 10066 THEN
            exp_f := 16;
        ELSIF x =- 10065 THEN
            exp_f := 16;
        ELSIF x =- 10064 THEN
            exp_f := 16;
        ELSIF x =- 10063 THEN
            exp_f := 16;
        ELSIF x =- 10062 THEN
            exp_f := 16;
        ELSIF x =- 10061 THEN
            exp_f := 16;
        ELSIF x =- 10060 THEN
            exp_f := 16;
        ELSIF x =- 10059 THEN
            exp_f := 16;
        ELSIF x =- 10058 THEN
            exp_f := 16;
        ELSIF x =- 10057 THEN
            exp_f := 16;
        ELSIF x =- 10056 THEN
            exp_f := 16;
        ELSIF x =- 10055 THEN
            exp_f := 16;
        ELSIF x =- 10054 THEN
            exp_f := 16;
        ELSIF x =- 10053 THEN
            exp_f := 16;
        ELSIF x =- 10052 THEN
            exp_f := 16;
        ELSIF x =- 10051 THEN
            exp_f := 16;
        ELSIF x =- 10050 THEN
            exp_f := 16;
        ELSIF x =- 10049 THEN
            exp_f := 16;
        ELSIF x =- 10048 THEN
            exp_f := 16;
        ELSIF x =- 10047 THEN
            exp_f := 16;
        ELSIF x =- 10046 THEN
            exp_f := 16;
        ELSIF x =- 10045 THEN
            exp_f := 16;
        ELSIF x =- 10044 THEN
            exp_f := 16;
        ELSIF x =- 10043 THEN
            exp_f := 16;
        ELSIF x =- 10042 THEN
            exp_f := 16;
        ELSIF x =- 10041 THEN
            exp_f := 16;
        ELSIF x =- 10040 THEN
            exp_f := 16;
        ELSIF x =- 10039 THEN
            exp_f := 16;
        ELSIF x =- 10038 THEN
            exp_f := 16;
        ELSIF x =- 10037 THEN
            exp_f := 16;
        ELSIF x =- 10036 THEN
            exp_f := 16;
        ELSIF x =- 10035 THEN
            exp_f := 16;
        ELSIF x =- 10034 THEN
            exp_f := 16;
        ELSIF x =- 10033 THEN
            exp_f := 16;
        ELSIF x =- 10032 THEN
            exp_f := 16;
        ELSIF x =- 10031 THEN
            exp_f := 16;
        ELSIF x =- 10030 THEN
            exp_f := 16;
        ELSIF x =- 10029 THEN
            exp_f := 16;
        ELSIF x =- 10028 THEN
            exp_f := 16;
        ELSIF x =- 10027 THEN
            exp_f := 16;
        ELSIF x =- 10026 THEN
            exp_f := 16;
        ELSIF x =- 10025 THEN
            exp_f := 16;
        ELSIF x =- 10024 THEN
            exp_f := 16;
        ELSIF x =- 10023 THEN
            exp_f := 16;
        ELSIF x =- 10022 THEN
            exp_f := 16;
        ELSIF x =- 10021 THEN
            exp_f := 16;
        ELSIF x =- 10020 THEN
            exp_f := 16;
        ELSIF x =- 10019 THEN
            exp_f := 16;
        ELSIF x =- 10018 THEN
            exp_f := 16;
        ELSIF x =- 10017 THEN
            exp_f := 16;
        ELSIF x =- 10016 THEN
            exp_f := 16;
        ELSIF x =- 10015 THEN
            exp_f := 16;
        ELSIF x =- 10014 THEN
            exp_f := 16;
        ELSIF x =- 10013 THEN
            exp_f := 16;
        ELSIF x =- 10012 THEN
            exp_f := 16;
        ELSIF x =- 10011 THEN
            exp_f := 16;
        ELSIF x =- 10010 THEN
            exp_f := 16;
        ELSIF x =- 10009 THEN
            exp_f := 16;
        ELSIF x =- 10008 THEN
            exp_f := 16;
        ELSIF x =- 10007 THEN
            exp_f := 16;
        ELSIF x =- 10006 THEN
            exp_f := 16;
        ELSIF x =- 10005 THEN
            exp_f := 16;
        ELSIF x =- 10004 THEN
            exp_f := 16;
        ELSIF x =- 10003 THEN
            exp_f := 16;
        ELSIF x =- 10002 THEN
            exp_f := 16;
        ELSIF x =- 10001 THEN
            exp_f := 16;
        ELSIF x =- 10000 THEN
            exp_f := 16;
        ELSIF x =- 9999 THEN
            exp_f := 16;
        ELSIF x =- 9998 THEN
            exp_f := 16;
        ELSIF x =- 9997 THEN
            exp_f := 16;
        ELSIF x =- 9996 THEN
            exp_f := 16;
        ELSIF x =- 9995 THEN
            exp_f := 16;
        ELSIF x =- 9994 THEN
            exp_f := 16;
        ELSIF x =- 9993 THEN
            exp_f := 16;
        ELSIF x =- 9992 THEN
            exp_f := 16;
        ELSIF x =- 9991 THEN
            exp_f := 16;
        ELSIF x =- 9990 THEN
            exp_f := 16;
        ELSIF x =- 9989 THEN
            exp_f := 16;
        ELSIF x =- 9988 THEN
            exp_f := 16;
        ELSIF x =- 9987 THEN
            exp_f := 16;
        ELSIF x =- 9986 THEN
            exp_f := 16;
        ELSIF x =- 9985 THEN
            exp_f := 16;
        ELSIF x =- 9984 THEN
            exp_f := 16;
        ELSIF x =- 9983 THEN
            exp_f := 16;
        ELSIF x =- 9982 THEN
            exp_f := 16;
        ELSIF x =- 9981 THEN
            exp_f := 16;
        ELSIF x =- 9980 THEN
            exp_f := 16;
        ELSIF x =- 9979 THEN
            exp_f := 16;
        ELSIF x =- 9978 THEN
            exp_f := 16;
        ELSIF x =- 9977 THEN
            exp_f := 16;
        ELSIF x =- 9976 THEN
            exp_f := 16;
        ELSIF x =- 9975 THEN
            exp_f := 16;
        ELSIF x =- 9974 THEN
            exp_f := 16;
        ELSIF x =- 9973 THEN
            exp_f := 16;
        ELSIF x =- 9972 THEN
            exp_f := 16;
        ELSIF x =- 9971 THEN
            exp_f := 16;
        ELSIF x =- 9970 THEN
            exp_f := 16;
        ELSIF x =- 9969 THEN
            exp_f := 16;
        ELSIF x =- 9968 THEN
            exp_f := 16;
        ELSIF x =- 9967 THEN
            exp_f := 16;
        ELSIF x =- 9966 THEN
            exp_f := 16;
        ELSIF x =- 9965 THEN
            exp_f := 16;
        ELSIF x =- 9964 THEN
            exp_f := 16;
        ELSIF x =- 9963 THEN
            exp_f := 16;
        ELSIF x =- 9962 THEN
            exp_f := 16;
        ELSIF x =- 9961 THEN
            exp_f := 16;
        ELSIF x =- 9960 THEN
            exp_f := 16;
        ELSIF x =- 9959 THEN
            exp_f := 16;
        ELSIF x =- 9958 THEN
            exp_f := 16;
        ELSIF x =- 9957 THEN
            exp_f := 16;
        ELSIF x =- 9956 THEN
            exp_f := 16;
        ELSIF x =- 9955 THEN
            exp_f := 16;
        ELSIF x =- 9954 THEN
            exp_f := 16;
        ELSIF x =- 9953 THEN
            exp_f := 16;
        ELSIF x =- 9952 THEN
            exp_f := 16;
        ELSIF x =- 9951 THEN
            exp_f := 16;
        ELSIF x =- 9950 THEN
            exp_f := 16;
        ELSIF x =- 9949 THEN
            exp_f := 16;
        ELSIF x =- 9948 THEN
            exp_f := 16;
        ELSIF x =- 9947 THEN
            exp_f := 16;
        ELSIF x =- 9946 THEN
            exp_f := 16;
        ELSIF x =- 9945 THEN
            exp_f := 16;
        ELSIF x =- 9944 THEN
            exp_f := 16;
        ELSIF x =- 9943 THEN
            exp_f := 16;
        ELSIF x =- 9942 THEN
            exp_f := 16;
        ELSIF x =- 9941 THEN
            exp_f := 16;
        ELSIF x =- 9940 THEN
            exp_f := 16;
        ELSIF x =- 9939 THEN
            exp_f := 16;
        ELSIF x =- 9938 THEN
            exp_f := 16;
        ELSIF x =- 9937 THEN
            exp_f := 16;
        ELSIF x =- 9936 THEN
            exp_f := 16;
        ELSIF x =- 9935 THEN
            exp_f := 16;
        ELSIF x =- 9934 THEN
            exp_f := 16;
        ELSIF x =- 9933 THEN
            exp_f := 16;
        ELSIF x =- 9932 THEN
            exp_f := 16;
        ELSIF x =- 9931 THEN
            exp_f := 16;
        ELSIF x =- 9930 THEN
            exp_f := 16;
        ELSIF x =- 9929 THEN
            exp_f := 16;
        ELSIF x =- 9928 THEN
            exp_f := 16;
        ELSIF x =- 9927 THEN
            exp_f := 16;
        ELSIF x =- 9926 THEN
            exp_f := 16;
        ELSIF x =- 9925 THEN
            exp_f := 16;
        ELSIF x =- 9924 THEN
            exp_f := 17;
        ELSIF x =- 9923 THEN
            exp_f := 17;
        ELSIF x =- 9922 THEN
            exp_f := 17;
        ELSIF x =- 9921 THEN
            exp_f := 17;
        ELSIF x =- 9920 THEN
            exp_f := 17;
        ELSIF x =- 9919 THEN
            exp_f := 17;
        ELSIF x =- 9918 THEN
            exp_f := 17;
        ELSIF x =- 9917 THEN
            exp_f := 17;
        ELSIF x =- 9916 THEN
            exp_f := 17;
        ELSIF x =- 9915 THEN
            exp_f := 17;
        ELSIF x =- 9914 THEN
            exp_f := 17;
        ELSIF x =- 9913 THEN
            exp_f := 17;
        ELSIF x =- 9912 THEN
            exp_f := 17;
        ELSIF x =- 9911 THEN
            exp_f := 17;
        ELSIF x =- 9910 THEN
            exp_f := 17;
        ELSIF x =- 9909 THEN
            exp_f := 17;
        ELSIF x =- 9908 THEN
            exp_f := 17;
        ELSIF x =- 9907 THEN
            exp_f := 17;
        ELSIF x =- 9906 THEN
            exp_f := 17;
        ELSIF x =- 9905 THEN
            exp_f := 17;
        ELSIF x =- 9904 THEN
            exp_f := 17;
        ELSIF x =- 9903 THEN
            exp_f := 17;
        ELSIF x =- 9902 THEN
            exp_f := 17;
        ELSIF x =- 9901 THEN
            exp_f := 17;
        ELSIF x =- 9900 THEN
            exp_f := 17;
        ELSIF x =- 9899 THEN
            exp_f := 17;
        ELSIF x =- 9898 THEN
            exp_f := 17;
        ELSIF x =- 9897 THEN
            exp_f := 17;
        ELSIF x =- 9896 THEN
            exp_f := 17;
        ELSIF x =- 9895 THEN
            exp_f := 17;
        ELSIF x =- 9894 THEN
            exp_f := 17;
        ELSIF x =- 9893 THEN
            exp_f := 17;
        ELSIF x =- 9892 THEN
            exp_f := 17;
        ELSIF x =- 9891 THEN
            exp_f := 17;
        ELSIF x =- 9890 THEN
            exp_f := 17;
        ELSIF x =- 9889 THEN
            exp_f := 17;
        ELSIF x =- 9888 THEN
            exp_f := 17;
        ELSIF x =- 9887 THEN
            exp_f := 17;
        ELSIF x =- 9886 THEN
            exp_f := 17;
        ELSIF x =- 9885 THEN
            exp_f := 17;
        ELSIF x =- 9884 THEN
            exp_f := 17;
        ELSIF x =- 9883 THEN
            exp_f := 17;
        ELSIF x =- 9882 THEN
            exp_f := 17;
        ELSIF x =- 9881 THEN
            exp_f := 17;
        ELSIF x =- 9880 THEN
            exp_f := 17;
        ELSIF x =- 9879 THEN
            exp_f := 17;
        ELSIF x =- 9878 THEN
            exp_f := 17;
        ELSIF x =- 9877 THEN
            exp_f := 17;
        ELSIF x =- 9876 THEN
            exp_f := 17;
        ELSIF x =- 9875 THEN
            exp_f := 17;
        ELSIF x =- 9874 THEN
            exp_f := 17;
        ELSIF x =- 9873 THEN
            exp_f := 17;
        ELSIF x =- 9872 THEN
            exp_f := 17;
        ELSIF x =- 9871 THEN
            exp_f := 17;
        ELSIF x =- 9870 THEN
            exp_f := 17;
        ELSIF x =- 9869 THEN
            exp_f := 17;
        ELSIF x =- 9868 THEN
            exp_f := 17;
        ELSIF x =- 9867 THEN
            exp_f := 17;
        ELSIF x =- 9866 THEN
            exp_f := 17;
        ELSIF x =- 9865 THEN
            exp_f := 17;
        ELSIF x =- 9864 THEN
            exp_f := 17;
        ELSIF x =- 9863 THEN
            exp_f := 17;
        ELSIF x =- 9862 THEN
            exp_f := 17;
        ELSIF x =- 9861 THEN
            exp_f := 17;
        ELSIF x =- 9860 THEN
            exp_f := 17;
        ELSIF x =- 9859 THEN
            exp_f := 17;
        ELSIF x =- 9858 THEN
            exp_f := 17;
        ELSIF x =- 9857 THEN
            exp_f := 17;
        ELSIF x =- 9856 THEN
            exp_f := 17;
        ELSIF x =- 9855 THEN
            exp_f := 17;
        ELSIF x =- 9854 THEN
            exp_f := 17;
        ELSIF x =- 9853 THEN
            exp_f := 17;
        ELSIF x =- 9852 THEN
            exp_f := 17;
        ELSIF x =- 9851 THEN
            exp_f := 17;
        ELSIF x =- 9850 THEN
            exp_f := 17;
        ELSIF x =- 9849 THEN
            exp_f := 17;
        ELSIF x =- 9848 THEN
            exp_f := 17;
        ELSIF x =- 9847 THEN
            exp_f := 17;
        ELSIF x =- 9846 THEN
            exp_f := 17;
        ELSIF x =- 9845 THEN
            exp_f := 17;
        ELSIF x =- 9844 THEN
            exp_f := 17;
        ELSIF x =- 9843 THEN
            exp_f := 17;
        ELSIF x =- 9842 THEN
            exp_f := 17;
        ELSIF x =- 9841 THEN
            exp_f := 17;
        ELSIF x =- 9840 THEN
            exp_f := 17;
        ELSIF x =- 9839 THEN
            exp_f := 17;
        ELSIF x =- 9838 THEN
            exp_f := 17;
        ELSIF x =- 9837 THEN
            exp_f := 17;
        ELSIF x =- 9836 THEN
            exp_f := 17;
        ELSIF x =- 9835 THEN
            exp_f := 17;
        ELSIF x =- 9834 THEN
            exp_f := 17;
        ELSIF x =- 9833 THEN
            exp_f := 17;
        ELSIF x =- 9832 THEN
            exp_f := 17;
        ELSIF x =- 9831 THEN
            exp_f := 17;
        ELSIF x =- 9830 THEN
            exp_f := 17;
        ELSIF x =- 9829 THEN
            exp_f := 17;
        ELSIF x =- 9828 THEN
            exp_f := 17;
        ELSIF x =- 9827 THEN
            exp_f := 17;
        ELSIF x =- 9826 THEN
            exp_f := 17;
        ELSIF x =- 9825 THEN
            exp_f := 17;
        ELSIF x =- 9824 THEN
            exp_f := 17;
        ELSIF x =- 9823 THEN
            exp_f := 17;
        ELSIF x =- 9822 THEN
            exp_f := 17;
        ELSIF x =- 9821 THEN
            exp_f := 17;
        ELSIF x =- 9820 THEN
            exp_f := 17;
        ELSIF x =- 9819 THEN
            exp_f := 17;
        ELSIF x =- 9818 THEN
            exp_f := 17;
        ELSIF x =- 9817 THEN
            exp_f := 17;
        ELSIF x =- 9816 THEN
            exp_f := 17;
        ELSIF x =- 9815 THEN
            exp_f := 17;
        ELSIF x =- 9814 THEN
            exp_f := 17;
        ELSIF x =- 9813 THEN
            exp_f := 17;
        ELSIF x =- 9812 THEN
            exp_f := 17;
        ELSIF x =- 9811 THEN
            exp_f := 17;
        ELSIF x =- 9810 THEN
            exp_f := 17;
        ELSIF x =- 9809 THEN
            exp_f := 17;
        ELSIF x =- 9808 THEN
            exp_f := 17;
        ELSIF x =- 9807 THEN
            exp_f := 17;
        ELSIF x =- 9806 THEN
            exp_f := 17;
        ELSIF x =- 9805 THEN
            exp_f := 17;
        ELSIF x =- 9804 THEN
            exp_f := 17;
        ELSIF x =- 9803 THEN
            exp_f := 17;
        ELSIF x =- 9802 THEN
            exp_f := 17;
        ELSIF x =- 9801 THEN
            exp_f := 17;
        ELSIF x =- 9800 THEN
            exp_f := 17;
        ELSIF x =- 9799 THEN
            exp_f := 17;
        ELSIF x =- 9798 THEN
            exp_f := 17;
        ELSIF x =- 9797 THEN
            exp_f := 17;
        ELSIF x =- 9796 THEN
            exp_f := 17;
        ELSIF x =- 9795 THEN
            exp_f := 17;
        ELSIF x =- 9794 THEN
            exp_f := 17;
        ELSIF x =- 9793 THEN
            exp_f := 17;
        ELSIF x =- 9792 THEN
            exp_f := 17;
        ELSIF x =- 9791 THEN
            exp_f := 17;
        ELSIF x =- 9790 THEN
            exp_f := 17;
        ELSIF x =- 9789 THEN
            exp_f := 17;
        ELSIF x =- 9788 THEN
            exp_f := 17;
        ELSIF x =- 9787 THEN
            exp_f := 17;
        ELSIF x =- 9786 THEN
            exp_f := 17;
        ELSIF x =- 9785 THEN
            exp_f := 17;
        ELSIF x =- 9784 THEN
            exp_f := 17;
        ELSIF x =- 9783 THEN
            exp_f := 17;
        ELSIF x =- 9782 THEN
            exp_f := 17;
        ELSIF x =- 9781 THEN
            exp_f := 17;
        ELSIF x =- 9780 THEN
            exp_f := 17;
        ELSIF x =- 9779 THEN
            exp_f := 17;
        ELSIF x =- 9778 THEN
            exp_f := 17;
        ELSIF x =- 9777 THEN
            exp_f := 17;
        ELSIF x =- 9776 THEN
            exp_f := 17;
        ELSIF x =- 9775 THEN
            exp_f := 17;
        ELSIF x =- 9774 THEN
            exp_f := 17;
        ELSIF x =- 9773 THEN
            exp_f := 17;
        ELSIF x =- 9772 THEN
            exp_f := 17;
        ELSIF x =- 9771 THEN
            exp_f := 17;
        ELSIF x =- 9770 THEN
            exp_f := 17;
        ELSIF x =- 9769 THEN
            exp_f := 17;
        ELSIF x =- 9768 THEN
            exp_f := 17;
        ELSIF x =- 9767 THEN
            exp_f := 18;
        ELSIF x =- 9766 THEN
            exp_f := 18;
        ELSIF x =- 9765 THEN
            exp_f := 18;
        ELSIF x =- 9764 THEN
            exp_f := 18;
        ELSIF x =- 9763 THEN
            exp_f := 18;
        ELSIF x =- 9762 THEN
            exp_f := 18;
        ELSIF x =- 9761 THEN
            exp_f := 18;
        ELSIF x =- 9760 THEN
            exp_f := 18;
        ELSIF x =- 9759 THEN
            exp_f := 18;
        ELSIF x =- 9758 THEN
            exp_f := 18;
        ELSIF x =- 9757 THEN
            exp_f := 18;
        ELSIF x =- 9756 THEN
            exp_f := 18;
        ELSIF x =- 9755 THEN
            exp_f := 18;
        ELSIF x =- 9754 THEN
            exp_f := 18;
        ELSIF x =- 9753 THEN
            exp_f := 18;
        ELSIF x =- 9752 THEN
            exp_f := 18;
        ELSIF x =- 9751 THEN
            exp_f := 18;
        ELSIF x =- 9750 THEN
            exp_f := 18;
        ELSIF x =- 9749 THEN
            exp_f := 18;
        ELSIF x =- 9748 THEN
            exp_f := 18;
        ELSIF x =- 9747 THEN
            exp_f := 18;
        ELSIF x =- 9746 THEN
            exp_f := 18;
        ELSIF x =- 9745 THEN
            exp_f := 18;
        ELSIF x =- 9744 THEN
            exp_f := 18;
        ELSIF x =- 9743 THEN
            exp_f := 18;
        ELSIF x =- 9742 THEN
            exp_f := 18;
        ELSIF x =- 9741 THEN
            exp_f := 18;
        ELSIF x =- 9740 THEN
            exp_f := 18;
        ELSIF x =- 9739 THEN
            exp_f := 18;
        ELSIF x =- 9738 THEN
            exp_f := 18;
        ELSIF x =- 9737 THEN
            exp_f := 18;
        ELSIF x =- 9736 THEN
            exp_f := 18;
        ELSIF x =- 9735 THEN
            exp_f := 18;
        ELSIF x =- 9734 THEN
            exp_f := 18;
        ELSIF x =- 9733 THEN
            exp_f := 18;
        ELSIF x =- 9732 THEN
            exp_f := 18;
        ELSIF x =- 9731 THEN
            exp_f := 18;
        ELSIF x =- 9730 THEN
            exp_f := 18;
        ELSIF x =- 9729 THEN
            exp_f := 18;
        ELSIF x =- 9728 THEN
            exp_f := 18;
        ELSIF x =- 9727 THEN
            exp_f := 18;
        ELSIF x =- 9726 THEN
            exp_f := 18;
        ELSIF x =- 9725 THEN
            exp_f := 18;
        ELSIF x =- 9724 THEN
            exp_f := 18;
        ELSIF x =- 9723 THEN
            exp_f := 18;
        ELSIF x =- 9722 THEN
            exp_f := 18;
        ELSIF x =- 9721 THEN
            exp_f := 18;
        ELSIF x =- 9720 THEN
            exp_f := 18;
        ELSIF x =- 9719 THEN
            exp_f := 18;
        ELSIF x =- 9718 THEN
            exp_f := 18;
        ELSIF x =- 9717 THEN
            exp_f := 18;
        ELSIF x =- 9716 THEN
            exp_f := 18;
        ELSIF x =- 9715 THEN
            exp_f := 18;
        ELSIF x =- 9714 THEN
            exp_f := 18;
        ELSIF x =- 9713 THEN
            exp_f := 18;
        ELSIF x =- 9712 THEN
            exp_f := 18;
        ELSIF x =- 9711 THEN
            exp_f := 18;
        ELSIF x =- 9710 THEN
            exp_f := 18;
        ELSIF x =- 9709 THEN
            exp_f := 18;
        ELSIF x =- 9708 THEN
            exp_f := 18;
        ELSIF x =- 9707 THEN
            exp_f := 18;
        ELSIF x =- 9706 THEN
            exp_f := 18;
        ELSIF x =- 9705 THEN
            exp_f := 18;
        ELSIF x =- 9704 THEN
            exp_f := 18;
        ELSIF x =- 9703 THEN
            exp_f := 18;
        ELSIF x =- 9702 THEN
            exp_f := 18;
        ELSIF x =- 9701 THEN
            exp_f := 18;
        ELSIF x =- 9700 THEN
            exp_f := 18;
        ELSIF x =- 9699 THEN
            exp_f := 18;
        ELSIF x =- 9698 THEN
            exp_f := 18;
        ELSIF x =- 9697 THEN
            exp_f := 18;
        ELSIF x =- 9696 THEN
            exp_f := 18;
        ELSIF x =- 9695 THEN
            exp_f := 18;
        ELSIF x =- 9694 THEN
            exp_f := 18;
        ELSIF x =- 9693 THEN
            exp_f := 18;
        ELSIF x =- 9692 THEN
            exp_f := 18;
        ELSIF x =- 9691 THEN
            exp_f := 18;
        ELSIF x =- 9690 THEN
            exp_f := 18;
        ELSIF x =- 9689 THEN
            exp_f := 18;
        ELSIF x =- 9688 THEN
            exp_f := 18;
        ELSIF x =- 9687 THEN
            exp_f := 18;
        ELSIF x =- 9686 THEN
            exp_f := 18;
        ELSIF x =- 9685 THEN
            exp_f := 18;
        ELSIF x =- 9684 THEN
            exp_f := 18;
        ELSIF x =- 9683 THEN
            exp_f := 18;
        ELSIF x =- 9682 THEN
            exp_f := 18;
        ELSIF x =- 9681 THEN
            exp_f := 18;
        ELSIF x =- 9680 THEN
            exp_f := 18;
        ELSIF x =- 9679 THEN
            exp_f := 18;
        ELSIF x =- 9678 THEN
            exp_f := 18;
        ELSIF x =- 9677 THEN
            exp_f := 18;
        ELSIF x =- 9676 THEN
            exp_f := 18;
        ELSIF x =- 9675 THEN
            exp_f := 18;
        ELSIF x =- 9674 THEN
            exp_f := 18;
        ELSIF x =- 9673 THEN
            exp_f := 18;
        ELSIF x =- 9672 THEN
            exp_f := 18;
        ELSIF x =- 9671 THEN
            exp_f := 18;
        ELSIF x =- 9670 THEN
            exp_f := 18;
        ELSIF x =- 9669 THEN
            exp_f := 18;
        ELSIF x =- 9668 THEN
            exp_f := 18;
        ELSIF x =- 9667 THEN
            exp_f := 18;
        ELSIF x =- 9666 THEN
            exp_f := 18;
        ELSIF x =- 9665 THEN
            exp_f := 18;
        ELSIF x =- 9664 THEN
            exp_f := 18;
        ELSIF x =- 9663 THEN
            exp_f := 18;
        ELSIF x =- 9662 THEN
            exp_f := 18;
        ELSIF x =- 9661 THEN
            exp_f := 18;
        ELSIF x =- 9660 THEN
            exp_f := 18;
        ELSIF x =- 9659 THEN
            exp_f := 18;
        ELSIF x =- 9658 THEN
            exp_f := 18;
        ELSIF x =- 9657 THEN
            exp_f := 18;
        ELSIF x =- 9656 THEN
            exp_f := 18;
        ELSIF x =- 9655 THEN
            exp_f := 18;
        ELSIF x =- 9654 THEN
            exp_f := 19;
        ELSIF x =- 9653 THEN
            exp_f := 19;
        ELSIF x =- 9652 THEN
            exp_f := 19;
        ELSIF x =- 9651 THEN
            exp_f := 19;
        ELSIF x =- 9650 THEN
            exp_f := 19;
        ELSIF x =- 9649 THEN
            exp_f := 19;
        ELSIF x =- 9648 THEN
            exp_f := 19;
        ELSIF x =- 9647 THEN
            exp_f := 19;
        ELSIF x =- 9646 THEN
            exp_f := 19;
        ELSIF x =- 9645 THEN
            exp_f := 19;
        ELSIF x =- 9644 THEN
            exp_f := 19;
        ELSIF x =- 9643 THEN
            exp_f := 19;
        ELSIF x =- 9642 THEN
            exp_f := 19;
        ELSIF x =- 9641 THEN
            exp_f := 19;
        ELSIF x =- 9640 THEN
            exp_f := 19;
        ELSIF x =- 9639 THEN
            exp_f := 19;
        ELSIF x =- 9638 THEN
            exp_f := 19;
        ELSIF x =- 9637 THEN
            exp_f := 19;
        ELSIF x =- 9636 THEN
            exp_f := 19;
        ELSIF x =- 9635 THEN
            exp_f := 19;
        ELSIF x =- 9634 THEN
            exp_f := 19;
        ELSIF x =- 9633 THEN
            exp_f := 19;
        ELSIF x =- 9632 THEN
            exp_f := 19;
        ELSIF x =- 9631 THEN
            exp_f := 19;
        ELSIF x =- 9630 THEN
            exp_f := 19;
        ELSIF x =- 9629 THEN
            exp_f := 19;
        ELSIF x =- 9628 THEN
            exp_f := 19;
        ELSIF x =- 9627 THEN
            exp_f := 19;
        ELSIF x =- 9626 THEN
            exp_f := 19;
        ELSIF x =- 9625 THEN
            exp_f := 19;
        ELSIF x =- 9624 THEN
            exp_f := 19;
        ELSIF x =- 9623 THEN
            exp_f := 19;
        ELSIF x =- 9622 THEN
            exp_f := 19;
        ELSIF x =- 9621 THEN
            exp_f := 19;
        ELSIF x =- 9620 THEN
            exp_f := 19;
        ELSIF x =- 9619 THEN
            exp_f := 19;
        ELSIF x =- 9618 THEN
            exp_f := 19;
        ELSIF x =- 9617 THEN
            exp_f := 19;
        ELSIF x =- 9616 THEN
            exp_f := 19;
        ELSIF x =- 9615 THEN
            exp_f := 19;
        ELSIF x =- 9614 THEN
            exp_f := 19;
        ELSIF x =- 9613 THEN
            exp_f := 19;
        ELSIF x =- 9612 THEN
            exp_f := 19;
        ELSIF x =- 9611 THEN
            exp_f := 19;
        ELSIF x =- 9610 THEN
            exp_f := 19;
        ELSIF x =- 9609 THEN
            exp_f := 19;
        ELSIF x =- 9608 THEN
            exp_f := 19;
        ELSIF x =- 9607 THEN
            exp_f := 19;
        ELSIF x =- 9606 THEN
            exp_f := 19;
        ELSIF x =- 9605 THEN
            exp_f := 19;
        ELSIF x =- 9604 THEN
            exp_f := 19;
        ELSIF x =- 9603 THEN
            exp_f := 19;
        ELSIF x =- 9602 THEN
            exp_f := 19;
        ELSIF x =- 9601 THEN
            exp_f := 19;
        ELSIF x =- 9600 THEN
            exp_f := 19;
        ELSIF x =- 9599 THEN
            exp_f := 19;
        ELSIF x =- 9598 THEN
            exp_f := 19;
        ELSIF x =- 9597 THEN
            exp_f := 19;
        ELSIF x =- 9596 THEN
            exp_f := 19;
        ELSIF x =- 9595 THEN
            exp_f := 19;
        ELSIF x =- 9594 THEN
            exp_f := 19;
        ELSIF x =- 9593 THEN
            exp_f := 19;
        ELSIF x =- 9592 THEN
            exp_f := 19;
        ELSIF x =- 9591 THEN
            exp_f := 19;
        ELSIF x =- 9590 THEN
            exp_f := 19;
        ELSIF x =- 9589 THEN
            exp_f := 19;
        ELSIF x =- 9588 THEN
            exp_f := 19;
        ELSIF x =- 9587 THEN
            exp_f := 19;
        ELSIF x =- 9586 THEN
            exp_f := 19;
        ELSIF x =- 9585 THEN
            exp_f := 19;
        ELSIF x =- 9584 THEN
            exp_f := 19;
        ELSIF x =- 9583 THEN
            exp_f := 19;
        ELSIF x =- 9582 THEN
            exp_f := 19;
        ELSIF x =- 9581 THEN
            exp_f := 19;
        ELSIF x =- 9580 THEN
            exp_f := 19;
        ELSIF x =- 9579 THEN
            exp_f := 19;
        ELSIF x =- 9578 THEN
            exp_f := 19;
        ELSIF x =- 9577 THEN
            exp_f := 19;
        ELSIF x =- 9576 THEN
            exp_f := 19;
        ELSIF x =- 9575 THEN
            exp_f := 19;
        ELSIF x =- 9574 THEN
            exp_f := 19;
        ELSIF x =- 9573 THEN
            exp_f := 19;
        ELSIF x =- 9572 THEN
            exp_f := 19;
        ELSIF x =- 9571 THEN
            exp_f := 19;
        ELSIF x =- 9570 THEN
            exp_f := 19;
        ELSIF x =- 9569 THEN
            exp_f := 19;
        ELSIF x =- 9568 THEN
            exp_f := 19;
        ELSIF x =- 9567 THEN
            exp_f := 19;
        ELSIF x =- 9566 THEN
            exp_f := 19;
        ELSIF x =- 9565 THEN
            exp_f := 19;
        ELSIF x =- 9564 THEN
            exp_f := 19;
        ELSIF x =- 9563 THEN
            exp_f := 19;
        ELSIF x =- 9562 THEN
            exp_f := 19;
        ELSIF x =- 9561 THEN
            exp_f := 19;
        ELSIF x =- 9560 THEN
            exp_f := 19;
        ELSIF x =- 9559 THEN
            exp_f := 19;
        ELSIF x =- 9558 THEN
            exp_f := 19;
        ELSIF x =- 9557 THEN
            exp_f := 20;
        ELSIF x =- 9556 THEN
            exp_f := 20;
        ELSIF x =- 9555 THEN
            exp_f := 20;
        ELSIF x =- 9554 THEN
            exp_f := 20;
        ELSIF x =- 9553 THEN
            exp_f := 20;
        ELSIF x =- 9552 THEN
            exp_f := 20;
        ELSIF x =- 9551 THEN
            exp_f := 20;
        ELSIF x =- 9550 THEN
            exp_f := 20;
        ELSIF x =- 9549 THEN
            exp_f := 20;
        ELSIF x =- 9548 THEN
            exp_f := 20;
        ELSIF x =- 9547 THEN
            exp_f := 20;
        ELSIF x =- 9546 THEN
            exp_f := 20;
        ELSIF x =- 9545 THEN
            exp_f := 20;
        ELSIF x =- 9544 THEN
            exp_f := 20;
        ELSIF x =- 9543 THEN
            exp_f := 20;
        ELSIF x =- 9542 THEN
            exp_f := 20;
        ELSIF x =- 9541 THEN
            exp_f := 20;
        ELSIF x =- 9540 THEN
            exp_f := 20;
        ELSIF x =- 9539 THEN
            exp_f := 20;
        ELSIF x =- 9538 THEN
            exp_f := 20;
        ELSIF x =- 9537 THEN
            exp_f := 20;
        ELSIF x =- 9536 THEN
            exp_f := 20;
        ELSIF x =- 9535 THEN
            exp_f := 20;
        ELSIF x =- 9534 THEN
            exp_f := 20;
        ELSIF x =- 9533 THEN
            exp_f := 20;
        ELSIF x =- 9532 THEN
            exp_f := 20;
        ELSIF x =- 9531 THEN
            exp_f := 20;
        ELSIF x =- 9530 THEN
            exp_f := 20;
        ELSIF x =- 9529 THEN
            exp_f := 20;
        ELSIF x =- 9528 THEN
            exp_f := 20;
        ELSIF x =- 9527 THEN
            exp_f := 20;
        ELSIF x =- 9526 THEN
            exp_f := 20;
        ELSIF x =- 9525 THEN
            exp_f := 20;
        ELSIF x =- 9524 THEN
            exp_f := 20;
        ELSIF x =- 9523 THEN
            exp_f := 20;
        ELSIF x =- 9522 THEN
            exp_f := 20;
        ELSIF x =- 9521 THEN
            exp_f := 20;
        ELSIF x =- 9520 THEN
            exp_f := 20;
        ELSIF x =- 9519 THEN
            exp_f := 20;
        ELSIF x =- 9518 THEN
            exp_f := 20;
        ELSIF x =- 9517 THEN
            exp_f := 20;
        ELSIF x =- 9516 THEN
            exp_f := 20;
        ELSIF x =- 9515 THEN
            exp_f := 20;
        ELSIF x =- 9514 THEN
            exp_f := 20;
        ELSIF x =- 9513 THEN
            exp_f := 20;
        ELSIF x =- 9512 THEN
            exp_f := 20;
        ELSIF x =- 9511 THEN
            exp_f := 20;
        ELSIF x =- 9510 THEN
            exp_f := 20;
        ELSIF x =- 9509 THEN
            exp_f := 20;
        ELSIF x =- 9508 THEN
            exp_f := 20;
        ELSIF x =- 9507 THEN
            exp_f := 20;
        ELSIF x =- 9506 THEN
            exp_f := 20;
        ELSIF x =- 9505 THEN
            exp_f := 20;
        ELSIF x =- 9504 THEN
            exp_f := 20;
        ELSIF x =- 9503 THEN
            exp_f := 20;
        ELSIF x =- 9502 THEN
            exp_f := 20;
        ELSIF x =- 9501 THEN
            exp_f := 20;
        ELSIF x =- 9500 THEN
            exp_f := 20;
        ELSIF x =- 9499 THEN
            exp_f := 20;
        ELSIF x =- 9498 THEN
            exp_f := 20;
        ELSIF x =- 9497 THEN
            exp_f := 20;
        ELSIF x =- 9496 THEN
            exp_f := 20;
        ELSIF x =- 9495 THEN
            exp_f := 20;
        ELSIF x =- 9494 THEN
            exp_f := 20;
        ELSIF x =- 9493 THEN
            exp_f := 20;
        ELSIF x =- 9492 THEN
            exp_f := 20;
        ELSIF x =- 9491 THEN
            exp_f := 20;
        ELSIF x =- 9490 THEN
            exp_f := 20;
        ELSIF x =- 9489 THEN
            exp_f := 20;
        ELSIF x =- 9488 THEN
            exp_f := 20;
        ELSIF x =- 9487 THEN
            exp_f := 20;
        ELSIF x =- 9486 THEN
            exp_f := 20;
        ELSIF x =- 9485 THEN
            exp_f := 20;
        ELSIF x =- 9484 THEN
            exp_f := 20;
        ELSIF x =- 9483 THEN
            exp_f := 20;
        ELSIF x =- 9482 THEN
            exp_f := 20;
        ELSIF x =- 9481 THEN
            exp_f := 20;
        ELSIF x =- 9480 THEN
            exp_f := 20;
        ELSIF x =- 9479 THEN
            exp_f := 20;
        ELSIF x =- 9478 THEN
            exp_f := 20;
        ELSIF x =- 9477 THEN
            exp_f := 20;
        ELSIF x =- 9476 THEN
            exp_f := 20;
        ELSIF x =- 9475 THEN
            exp_f := 20;
        ELSIF x =- 9474 THEN
            exp_f := 20;
        ELSIF x =- 9473 THEN
            exp_f := 20;
        ELSIF x =- 9472 THEN
            exp_f := 20;
        ELSIF x =- 9471 THEN
            exp_f := 20;
        ELSIF x =- 9470 THEN
            exp_f := 20;
        ELSIF x =- 9469 THEN
            exp_f := 20;
        ELSIF x =- 9468 THEN
            exp_f := 20;
        ELSIF x =- 9467 THEN
            exp_f := 20;
        ELSIF x =- 9466 THEN
            exp_f := 20;
        ELSIF x =- 9465 THEN
            exp_f := 20;
        ELSIF x =- 9464 THEN
            exp_f := 20;
        ELSIF x =- 9463 THEN
            exp_f := 20;
        ELSIF x =- 9462 THEN
            exp_f := 20;
        ELSIF x =- 9461 THEN
            exp_f := 20;
        ELSIF x =- 9460 THEN
            exp_f := 20;
        ELSIF x =- 9459 THEN
            exp_f := 21;
        ELSIF x =- 9458 THEN
            exp_f := 21;
        ELSIF x =- 9457 THEN
            exp_f := 21;
        ELSIF x =- 9456 THEN
            exp_f := 21;
        ELSIF x =- 9455 THEN
            exp_f := 21;
        ELSIF x =- 9454 THEN
            exp_f := 21;
        ELSIF x =- 9453 THEN
            exp_f := 21;
        ELSIF x =- 9452 THEN
            exp_f := 21;
        ELSIF x =- 9451 THEN
            exp_f := 21;
        ELSIF x =- 9450 THEN
            exp_f := 21;
        ELSIF x =- 9449 THEN
            exp_f := 21;
        ELSIF x =- 9448 THEN
            exp_f := 21;
        ELSIF x =- 9447 THEN
            exp_f := 21;
        ELSIF x =- 9446 THEN
            exp_f := 21;
        ELSIF x =- 9445 THEN
            exp_f := 21;
        ELSIF x =- 9444 THEN
            exp_f := 21;
        ELSIF x =- 9443 THEN
            exp_f := 21;
        ELSIF x =- 9442 THEN
            exp_f := 21;
        ELSIF x =- 9441 THEN
            exp_f := 21;
        ELSIF x =- 9440 THEN
            exp_f := 21;
        ELSIF x =- 9439 THEN
            exp_f := 21;
        ELSIF x =- 9438 THEN
            exp_f := 21;
        ELSIF x =- 9437 THEN
            exp_f := 21;
        ELSIF x =- 9436 THEN
            exp_f := 21;
        ELSIF x =- 9435 THEN
            exp_f := 21;
        ELSIF x =- 9434 THEN
            exp_f := 21;
        ELSIF x =- 9433 THEN
            exp_f := 21;
        ELSIF x =- 9432 THEN
            exp_f := 21;
        ELSIF x =- 9431 THEN
            exp_f := 21;
        ELSIF x =- 9430 THEN
            exp_f := 21;
        ELSIF x =- 9429 THEN
            exp_f := 21;
        ELSIF x =- 9428 THEN
            exp_f := 21;
        ELSIF x =- 9427 THEN
            exp_f := 21;
        ELSIF x =- 9426 THEN
            exp_f := 21;
        ELSIF x =- 9425 THEN
            exp_f := 21;
        ELSIF x =- 9424 THEN
            exp_f := 21;
        ELSIF x =- 9423 THEN
            exp_f := 21;
        ELSIF x =- 9422 THEN
            exp_f := 21;
        ELSIF x =- 9421 THEN
            exp_f := 21;
        ELSIF x =- 9420 THEN
            exp_f := 21;
        ELSIF x =- 9419 THEN
            exp_f := 21;
        ELSIF x =- 9418 THEN
            exp_f := 21;
        ELSIF x =- 9417 THEN
            exp_f := 21;
        ELSIF x =- 9416 THEN
            exp_f := 21;
        ELSIF x =- 9415 THEN
            exp_f := 21;
        ELSIF x =- 9414 THEN
            exp_f := 21;
        ELSIF x =- 9413 THEN
            exp_f := 21;
        ELSIF x =- 9412 THEN
            exp_f := 21;
        ELSIF x =- 9411 THEN
            exp_f := 21;
        ELSIF x =- 9410 THEN
            exp_f := 21;
        ELSIF x =- 9409 THEN
            exp_f := 21;
        ELSIF x =- 9408 THEN
            exp_f := 21;
        ELSIF x =- 9407 THEN
            exp_f := 21;
        ELSIF x =- 9406 THEN
            exp_f := 21;
        ELSIF x =- 9405 THEN
            exp_f := 21;
        ELSIF x =- 9404 THEN
            exp_f := 21;
        ELSIF x =- 9403 THEN
            exp_f := 21;
        ELSIF x =- 9402 THEN
            exp_f := 21;
        ELSIF x =- 9401 THEN
            exp_f := 21;
        ELSIF x =- 9400 THEN
            exp_f := 21;
        ELSIF x =- 9399 THEN
            exp_f := 21;
        ELSIF x =- 9398 THEN
            exp_f := 21;
        ELSIF x =- 9397 THEN
            exp_f := 21;
        ELSIF x =- 9396 THEN
            exp_f := 21;
        ELSIF x =- 9395 THEN
            exp_f := 21;
        ELSIF x =- 9394 THEN
            exp_f := 21;
        ELSIF x =- 9393 THEN
            exp_f := 21;
        ELSIF x =- 9392 THEN
            exp_f := 21;
        ELSIF x =- 9391 THEN
            exp_f := 21;
        ELSIF x =- 9390 THEN
            exp_f := 21;
        ELSIF x =- 9389 THEN
            exp_f := 21;
        ELSIF x =- 9388 THEN
            exp_f := 21;
        ELSIF x =- 9387 THEN
            exp_f := 21;
        ELSIF x =- 9386 THEN
            exp_f := 21;
        ELSIF x =- 9385 THEN
            exp_f := 21;
        ELSIF x =- 9384 THEN
            exp_f := 21;
        ELSIF x =- 9383 THEN
            exp_f := 21;
        ELSIF x =- 9382 THEN
            exp_f := 21;
        ELSIF x =- 9381 THEN
            exp_f := 21;
        ELSIF x =- 9380 THEN
            exp_f := 21;
        ELSIF x =- 9379 THEN
            exp_f := 21;
        ELSIF x =- 9378 THEN
            exp_f := 21;
        ELSIF x =- 9377 THEN
            exp_f := 21;
        ELSIF x =- 9376 THEN
            exp_f := 21;
        ELSIF x =- 9375 THEN
            exp_f := 21;
        ELSIF x =- 9374 THEN
            exp_f := 21;
        ELSIF x =- 9373 THEN
            exp_f := 21;
        ELSIF x =- 9372 THEN
            exp_f := 21;
        ELSIF x =- 9371 THEN
            exp_f := 21;
        ELSIF x =- 9370 THEN
            exp_f := 21;
        ELSIF x =- 9369 THEN
            exp_f := 21;
        ELSIF x =- 9368 THEN
            exp_f := 21;
        ELSIF x =- 9367 THEN
            exp_f := 21;
        ELSIF x =- 9366 THEN
            exp_f := 21;
        ELSIF x =- 9365 THEN
            exp_f := 21;
        ELSIF x =- 9364 THEN
            exp_f := 21;
        ELSIF x =- 9363 THEN
            exp_f := 21;
        ELSIF x =- 9362 THEN
            exp_f := 22;
        ELSIF x =- 9361 THEN
            exp_f := 22;
        ELSIF x =- 9360 THEN
            exp_f := 22;
        ELSIF x =- 9359 THEN
            exp_f := 22;
        ELSIF x =- 9358 THEN
            exp_f := 22;
        ELSIF x =- 9357 THEN
            exp_f := 22;
        ELSIF x =- 9356 THEN
            exp_f := 22;
        ELSIF x =- 9355 THEN
            exp_f := 22;
        ELSIF x =- 9354 THEN
            exp_f := 22;
        ELSIF x =- 9353 THEN
            exp_f := 22;
        ELSIF x =- 9352 THEN
            exp_f := 22;
        ELSIF x =- 9351 THEN
            exp_f := 22;
        ELSIF x =- 9350 THEN
            exp_f := 22;
        ELSIF x =- 9349 THEN
            exp_f := 22;
        ELSIF x =- 9348 THEN
            exp_f := 22;
        ELSIF x =- 9347 THEN
            exp_f := 22;
        ELSIF x =- 9346 THEN
            exp_f := 22;
        ELSIF x =- 9345 THEN
            exp_f := 22;
        ELSIF x =- 9344 THEN
            exp_f := 22;
        ELSIF x =- 9343 THEN
            exp_f := 22;
        ELSIF x =- 9342 THEN
            exp_f := 22;
        ELSIF x =- 9341 THEN
            exp_f := 22;
        ELSIF x =- 9340 THEN
            exp_f := 22;
        ELSIF x =- 9339 THEN
            exp_f := 22;
        ELSIF x =- 9338 THEN
            exp_f := 22;
        ELSIF x =- 9337 THEN
            exp_f := 22;
        ELSIF x =- 9336 THEN
            exp_f := 22;
        ELSIF x =- 9335 THEN
            exp_f := 22;
        ELSIF x =- 9334 THEN
            exp_f := 22;
        ELSIF x =- 9333 THEN
            exp_f := 22;
        ELSIF x =- 9332 THEN
            exp_f := 22;
        ELSIF x =- 9331 THEN
            exp_f := 22;
        ELSIF x =- 9330 THEN
            exp_f := 22;
        ELSIF x =- 9329 THEN
            exp_f := 22;
        ELSIF x =- 9328 THEN
            exp_f := 22;
        ELSIF x =- 9327 THEN
            exp_f := 22;
        ELSIF x =- 9326 THEN
            exp_f := 22;
        ELSIF x =- 9325 THEN
            exp_f := 22;
        ELSIF x =- 9324 THEN
            exp_f := 22;
        ELSIF x =- 9323 THEN
            exp_f := 22;
        ELSIF x =- 9322 THEN
            exp_f := 22;
        ELSIF x =- 9321 THEN
            exp_f := 22;
        ELSIF x =- 9320 THEN
            exp_f := 22;
        ELSIF x =- 9319 THEN
            exp_f := 22;
        ELSIF x =- 9318 THEN
            exp_f := 22;
        ELSIF x =- 9317 THEN
            exp_f := 22;
        ELSIF x =- 9316 THEN
            exp_f := 22;
        ELSIF x =- 9315 THEN
            exp_f := 22;
        ELSIF x =- 9314 THEN
            exp_f := 22;
        ELSIF x =- 9313 THEN
            exp_f := 22;
        ELSIF x =- 9312 THEN
            exp_f := 22;
        ELSIF x =- 9311 THEN
            exp_f := 22;
        ELSIF x =- 9310 THEN
            exp_f := 22;
        ELSIF x =- 9309 THEN
            exp_f := 22;
        ELSIF x =- 9308 THEN
            exp_f := 22;
        ELSIF x =- 9307 THEN
            exp_f := 22;
        ELSIF x =- 9306 THEN
            exp_f := 22;
        ELSIF x =- 9305 THEN
            exp_f := 22;
        ELSIF x =- 9304 THEN
            exp_f := 22;
        ELSIF x =- 9303 THEN
            exp_f := 22;
        ELSIF x =- 9302 THEN
            exp_f := 22;
        ELSIF x =- 9301 THEN
            exp_f := 22;
        ELSIF x =- 9300 THEN
            exp_f := 22;
        ELSIF x =- 9299 THEN
            exp_f := 22;
        ELSIF x =- 9298 THEN
            exp_f := 22;
        ELSIF x =- 9297 THEN
            exp_f := 22;
        ELSIF x =- 9296 THEN
            exp_f := 22;
        ELSIF x =- 9295 THEN
            exp_f := 22;
        ELSIF x =- 9294 THEN
            exp_f := 22;
        ELSIF x =- 9293 THEN
            exp_f := 22;
        ELSIF x =- 9292 THEN
            exp_f := 22;
        ELSIF x =- 9291 THEN
            exp_f := 22;
        ELSIF x =- 9290 THEN
            exp_f := 22;
        ELSIF x =- 9289 THEN
            exp_f := 22;
        ELSIF x =- 9288 THEN
            exp_f := 22;
        ELSIF x =- 9287 THEN
            exp_f := 22;
        ELSIF x =- 9286 THEN
            exp_f := 22;
        ELSIF x =- 9285 THEN
            exp_f := 22;
        ELSIF x =- 9284 THEN
            exp_f := 22;
        ELSIF x =- 9283 THEN
            exp_f := 22;
        ELSIF x =- 9282 THEN
            exp_f := 22;
        ELSIF x =- 9281 THEN
            exp_f := 22;
        ELSIF x =- 9280 THEN
            exp_f := 22;
        ELSIF x =- 9279 THEN
            exp_f := 22;
        ELSIF x =- 9278 THEN
            exp_f := 22;
        ELSIF x =- 9277 THEN
            exp_f := 22;
        ELSIF x =- 9276 THEN
            exp_f := 22;
        ELSIF x =- 9275 THEN
            exp_f := 22;
        ELSIF x =- 9274 THEN
            exp_f := 22;
        ELSIF x =- 9273 THEN
            exp_f := 22;
        ELSIF x =- 9272 THEN
            exp_f := 22;
        ELSIF x =- 9271 THEN
            exp_f := 22;
        ELSIF x =- 9270 THEN
            exp_f := 22;
        ELSIF x =- 9269 THEN
            exp_f := 22;
        ELSIF x =- 9268 THEN
            exp_f := 22;
        ELSIF x =- 9267 THEN
            exp_f := 22;
        ELSIF x =- 9266 THEN
            exp_f := 22;
        ELSIF x =- 9265 THEN
            exp_f := 22;
        ELSIF x =- 9264 THEN
            exp_f := 23;
        ELSIF x =- 9263 THEN
            exp_f := 23;
        ELSIF x =- 9262 THEN
            exp_f := 23;
        ELSIF x =- 9261 THEN
            exp_f := 23;
        ELSIF x =- 9260 THEN
            exp_f := 23;
        ELSIF x =- 9259 THEN
            exp_f := 23;
        ELSIF x =- 9258 THEN
            exp_f := 23;
        ELSIF x =- 9257 THEN
            exp_f := 23;
        ELSIF x =- 9256 THEN
            exp_f := 23;
        ELSIF x =- 9255 THEN
            exp_f := 23;
        ELSIF x =- 9254 THEN
            exp_f := 23;
        ELSIF x =- 9253 THEN
            exp_f := 23;
        ELSIF x =- 9252 THEN
            exp_f := 23;
        ELSIF x =- 9251 THEN
            exp_f := 23;
        ELSIF x =- 9250 THEN
            exp_f := 23;
        ELSIF x =- 9249 THEN
            exp_f := 23;
        ELSIF x =- 9248 THEN
            exp_f := 23;
        ELSIF x =- 9247 THEN
            exp_f := 23;
        ELSIF x =- 9246 THEN
            exp_f := 23;
        ELSIF x =- 9245 THEN
            exp_f := 23;
        ELSIF x =- 9244 THEN
            exp_f := 23;
        ELSIF x =- 9243 THEN
            exp_f := 23;
        ELSIF x =- 9242 THEN
            exp_f := 23;
        ELSIF x =- 9241 THEN
            exp_f := 23;
        ELSIF x =- 9240 THEN
            exp_f := 23;
        ELSIF x =- 9239 THEN
            exp_f := 23;
        ELSIF x =- 9238 THEN
            exp_f := 23;
        ELSIF x =- 9237 THEN
            exp_f := 23;
        ELSIF x =- 9236 THEN
            exp_f := 23;
        ELSIF x =- 9235 THEN
            exp_f := 23;
        ELSIF x =- 9234 THEN
            exp_f := 23;
        ELSIF x =- 9233 THEN
            exp_f := 23;
        ELSIF x =- 9232 THEN
            exp_f := 23;
        ELSIF x =- 9231 THEN
            exp_f := 23;
        ELSIF x =- 9230 THEN
            exp_f := 23;
        ELSIF x =- 9229 THEN
            exp_f := 23;
        ELSIF x =- 9228 THEN
            exp_f := 23;
        ELSIF x =- 9227 THEN
            exp_f := 23;
        ELSIF x =- 9226 THEN
            exp_f := 23;
        ELSIF x =- 9225 THEN
            exp_f := 23;
        ELSIF x =- 9224 THEN
            exp_f := 23;
        ELSIF x =- 9223 THEN
            exp_f := 23;
        ELSIF x =- 9222 THEN
            exp_f := 23;
        ELSIF x =- 9221 THEN
            exp_f := 23;
        ELSIF x =- 9220 THEN
            exp_f := 23;
        ELSIF x =- 9219 THEN
            exp_f := 23;
        ELSIF x =- 9218 THEN
            exp_f := 23;
        ELSIF x =- 9217 THEN
            exp_f := 23;
        ELSIF x =- 9216 THEN
            exp_f := 23;
        ELSIF x =- 9215 THEN
            exp_f := 23;
        ELSIF x =- 9214 THEN
            exp_f := 23;
        ELSIF x =- 9213 THEN
            exp_f := 23;
        ELSIF x =- 9212 THEN
            exp_f := 23;
        ELSIF x =- 9211 THEN
            exp_f := 23;
        ELSIF x =- 9210 THEN
            exp_f := 23;
        ELSIF x =- 9209 THEN
            exp_f := 23;
        ELSIF x =- 9208 THEN
            exp_f := 23;
        ELSIF x =- 9207 THEN
            exp_f := 23;
        ELSIF x =- 9206 THEN
            exp_f := 23;
        ELSIF x =- 9205 THEN
            exp_f := 23;
        ELSIF x =- 9204 THEN
            exp_f := 23;
        ELSIF x =- 9203 THEN
            exp_f := 23;
        ELSIF x =- 9202 THEN
            exp_f := 23;
        ELSIF x =- 9201 THEN
            exp_f := 23;
        ELSIF x =- 9200 THEN
            exp_f := 23;
        ELSIF x =- 9199 THEN
            exp_f := 23;
        ELSIF x =- 9198 THEN
            exp_f := 23;
        ELSIF x =- 9197 THEN
            exp_f := 23;
        ELSIF x =- 9196 THEN
            exp_f := 23;
        ELSIF x =- 9195 THEN
            exp_f := 23;
        ELSIF x =- 9194 THEN
            exp_f := 23;
        ELSIF x =- 9193 THEN
            exp_f := 23;
        ELSIF x =- 9192 THEN
            exp_f := 23;
        ELSIF x =- 9191 THEN
            exp_f := 23;
        ELSIF x =- 9190 THEN
            exp_f := 23;
        ELSIF x =- 9189 THEN
            exp_f := 23;
        ELSIF x =- 9188 THEN
            exp_f := 23;
        ELSIF x =- 9187 THEN
            exp_f := 23;
        ELSIF x =- 9186 THEN
            exp_f := 23;
        ELSIF x =- 9185 THEN
            exp_f := 23;
        ELSIF x =- 9184 THEN
            exp_f := 23;
        ELSIF x =- 9183 THEN
            exp_f := 23;
        ELSIF x =- 9182 THEN
            exp_f := 23;
        ELSIF x =- 9181 THEN
            exp_f := 23;
        ELSIF x =- 9180 THEN
            exp_f := 23;
        ELSIF x =- 9179 THEN
            exp_f := 23;
        ELSIF x =- 9178 THEN
            exp_f := 23;
        ELSIF x =- 9177 THEN
            exp_f := 23;
        ELSIF x =- 9176 THEN
            exp_f := 23;
        ELSIF x =- 9175 THEN
            exp_f := 24;
        ELSIF x =- 9174 THEN
            exp_f := 24;
        ELSIF x =- 9173 THEN
            exp_f := 24;
        ELSIF x =- 9172 THEN
            exp_f := 24;
        ELSIF x =- 9171 THEN
            exp_f := 24;
        ELSIF x =- 9170 THEN
            exp_f := 24;
        ELSIF x =- 9169 THEN
            exp_f := 24;
        ELSIF x =- 9168 THEN
            exp_f := 24;
        ELSIF x =- 9167 THEN
            exp_f := 24;
        ELSIF x =- 9166 THEN
            exp_f := 24;
        ELSIF x =- 9165 THEN
            exp_f := 24;
        ELSIF x =- 9164 THEN
            exp_f := 24;
        ELSIF x =- 9163 THEN
            exp_f := 24;
        ELSIF x =- 9162 THEN
            exp_f := 24;
        ELSIF x =- 9161 THEN
            exp_f := 24;
        ELSIF x =- 9160 THEN
            exp_f := 24;
        ELSIF x =- 9159 THEN
            exp_f := 24;
        ELSIF x =- 9158 THEN
            exp_f := 24;
        ELSIF x =- 9157 THEN
            exp_f := 24;
        ELSIF x =- 9156 THEN
            exp_f := 24;
        ELSIF x =- 9155 THEN
            exp_f := 24;
        ELSIF x =- 9154 THEN
            exp_f := 24;
        ELSIF x =- 9153 THEN
            exp_f := 24;
        ELSIF x =- 9152 THEN
            exp_f := 24;
        ELSIF x =- 9151 THEN
            exp_f := 24;
        ELSIF x =- 9150 THEN
            exp_f := 24;
        ELSIF x =- 9149 THEN
            exp_f := 24;
        ELSIF x =- 9148 THEN
            exp_f := 24;
        ELSIF x =- 9147 THEN
            exp_f := 24;
        ELSIF x =- 9146 THEN
            exp_f := 24;
        ELSIF x =- 9145 THEN
            exp_f := 24;
        ELSIF x =- 9144 THEN
            exp_f := 24;
        ELSIF x =- 9143 THEN
            exp_f := 24;
        ELSIF x =- 9142 THEN
            exp_f := 24;
        ELSIF x =- 9141 THEN
            exp_f := 24;
        ELSIF x =- 9140 THEN
            exp_f := 24;
        ELSIF x =- 9139 THEN
            exp_f := 24;
        ELSIF x =- 9138 THEN
            exp_f := 24;
        ELSIF x =- 9137 THEN
            exp_f := 24;
        ELSIF x =- 9136 THEN
            exp_f := 24;
        ELSIF x =- 9135 THEN
            exp_f := 24;
        ELSIF x =- 9134 THEN
            exp_f := 24;
        ELSIF x =- 9133 THEN
            exp_f := 24;
        ELSIF x =- 9132 THEN
            exp_f := 24;
        ELSIF x =- 9131 THEN
            exp_f := 24;
        ELSIF x =- 9130 THEN
            exp_f := 24;
        ELSIF x =- 9129 THEN
            exp_f := 24;
        ELSIF x =- 9128 THEN
            exp_f := 24;
        ELSIF x =- 9127 THEN
            exp_f := 24;
        ELSIF x =- 9126 THEN
            exp_f := 24;
        ELSIF x =- 9125 THEN
            exp_f := 24;
        ELSIF x =- 9124 THEN
            exp_f := 24;
        ELSIF x =- 9123 THEN
            exp_f := 24;
        ELSIF x =- 9122 THEN
            exp_f := 24;
        ELSIF x =- 9121 THEN
            exp_f := 24;
        ELSIF x =- 9120 THEN
            exp_f := 24;
        ELSIF x =- 9119 THEN
            exp_f := 24;
        ELSIF x =- 9118 THEN
            exp_f := 24;
        ELSIF x =- 9117 THEN
            exp_f := 24;
        ELSIF x =- 9116 THEN
            exp_f := 24;
        ELSIF x =- 9115 THEN
            exp_f := 24;
        ELSIF x =- 9114 THEN
            exp_f := 24;
        ELSIF x =- 9113 THEN
            exp_f := 24;
        ELSIF x =- 9112 THEN
            exp_f := 24;
        ELSIF x =- 9111 THEN
            exp_f := 24;
        ELSIF x =- 9110 THEN
            exp_f := 24;
        ELSIF x =- 9109 THEN
            exp_f := 24;
        ELSIF x =- 9108 THEN
            exp_f := 24;
        ELSIF x =- 9107 THEN
            exp_f := 24;
        ELSIF x =- 9106 THEN
            exp_f := 24;
        ELSIF x =- 9105 THEN
            exp_f := 24;
        ELSIF x =- 9104 THEN
            exp_f := 24;
        ELSIF x =- 9103 THEN
            exp_f := 24;
        ELSIF x =- 9102 THEN
            exp_f := 24;
        ELSIF x =- 9101 THEN
            exp_f := 24;
        ELSIF x =- 9100 THEN
            exp_f := 24;
        ELSIF x =- 9099 THEN
            exp_f := 24;
        ELSIF x =- 9098 THEN
            exp_f := 24;
        ELSIF x =- 9097 THEN
            exp_f := 24;
        ELSIF x =- 9096 THEN
            exp_f := 24;
        ELSIF x =- 9095 THEN
            exp_f := 24;
        ELSIF x =- 9094 THEN
            exp_f := 24;
        ELSIF x =- 9093 THEN
            exp_f := 25;
        ELSIF x =- 9092 THEN
            exp_f := 25;
        ELSIF x =- 9091 THEN
            exp_f := 25;
        ELSIF x =- 9090 THEN
            exp_f := 25;
        ELSIF x =- 9089 THEN
            exp_f := 25;
        ELSIF x =- 9088 THEN
            exp_f := 25;
        ELSIF x =- 9087 THEN
            exp_f := 25;
        ELSIF x =- 9086 THEN
            exp_f := 25;
        ELSIF x =- 9085 THEN
            exp_f := 25;
        ELSIF x =- 9084 THEN
            exp_f := 25;
        ELSIF x =- 9083 THEN
            exp_f := 25;
        ELSIF x =- 9082 THEN
            exp_f := 25;
        ELSIF x =- 9081 THEN
            exp_f := 25;
        ELSIF x =- 9080 THEN
            exp_f := 25;
        ELSIF x =- 9079 THEN
            exp_f := 25;
        ELSIF x =- 9078 THEN
            exp_f := 25;
        ELSIF x =- 9077 THEN
            exp_f := 25;
        ELSIF x =- 9076 THEN
            exp_f := 25;
        ELSIF x =- 9075 THEN
            exp_f := 25;
        ELSIF x =- 9074 THEN
            exp_f := 25;
        ELSIF x =- 9073 THEN
            exp_f := 25;
        ELSIF x =- 9072 THEN
            exp_f := 25;
        ELSIF x =- 9071 THEN
            exp_f := 25;
        ELSIF x =- 9070 THEN
            exp_f := 25;
        ELSIF x =- 9069 THEN
            exp_f := 25;
        ELSIF x =- 9068 THEN
            exp_f := 25;
        ELSIF x =- 9067 THEN
            exp_f := 25;
        ELSIF x =- 9066 THEN
            exp_f := 25;
        ELSIF x =- 9065 THEN
            exp_f := 25;
        ELSIF x =- 9064 THEN
            exp_f := 25;
        ELSIF x =- 9063 THEN
            exp_f := 25;
        ELSIF x =- 9062 THEN
            exp_f := 25;
        ELSIF x =- 9061 THEN
            exp_f := 25;
        ELSIF x =- 9060 THEN
            exp_f := 25;
        ELSIF x =- 9059 THEN
            exp_f := 25;
        ELSIF x =- 9058 THEN
            exp_f := 25;
        ELSIF x =- 9057 THEN
            exp_f := 25;
        ELSIF x =- 9056 THEN
            exp_f := 25;
        ELSIF x =- 9055 THEN
            exp_f := 25;
        ELSIF x =- 9054 THEN
            exp_f := 25;
        ELSIF x =- 9053 THEN
            exp_f := 25;
        ELSIF x =- 9052 THEN
            exp_f := 25;
        ELSIF x =- 9051 THEN
            exp_f := 25;
        ELSIF x =- 9050 THEN
            exp_f := 25;
        ELSIF x =- 9049 THEN
            exp_f := 25;
        ELSIF x =- 9048 THEN
            exp_f := 25;
        ELSIF x =- 9047 THEN
            exp_f := 25;
        ELSIF x =- 9046 THEN
            exp_f := 25;
        ELSIF x =- 9045 THEN
            exp_f := 25;
        ELSIF x =- 9044 THEN
            exp_f := 25;
        ELSIF x =- 9043 THEN
            exp_f := 25;
        ELSIF x =- 9042 THEN
            exp_f := 25;
        ELSIF x =- 9041 THEN
            exp_f := 25;
        ELSIF x =- 9040 THEN
            exp_f := 25;
        ELSIF x =- 9039 THEN
            exp_f := 25;
        ELSIF x =- 9038 THEN
            exp_f := 25;
        ELSIF x =- 9037 THEN
            exp_f := 25;
        ELSIF x =- 9036 THEN
            exp_f := 25;
        ELSIF x =- 9035 THEN
            exp_f := 25;
        ELSIF x =- 9034 THEN
            exp_f := 25;
        ELSIF x =- 9033 THEN
            exp_f := 25;
        ELSIF x =- 9032 THEN
            exp_f := 25;
        ELSIF x =- 9031 THEN
            exp_f := 25;
        ELSIF x =- 9030 THEN
            exp_f := 25;
        ELSIF x =- 9029 THEN
            exp_f := 25;
        ELSIF x =- 9028 THEN
            exp_f := 25;
        ELSIF x =- 9027 THEN
            exp_f := 25;
        ELSIF x =- 9026 THEN
            exp_f := 25;
        ELSIF x =- 9025 THEN
            exp_f := 25;
        ELSIF x =- 9024 THEN
            exp_f := 25;
        ELSIF x =- 9023 THEN
            exp_f := 25;
        ELSIF x =- 9022 THEN
            exp_f := 25;
        ELSIF x =- 9021 THEN
            exp_f := 25;
        ELSIF x =- 9020 THEN
            exp_f := 25;
        ELSIF x =- 9019 THEN
            exp_f := 25;
        ELSIF x =- 9018 THEN
            exp_f := 25;
        ELSIF x =- 9017 THEN
            exp_f := 25;
        ELSIF x =- 9016 THEN
            exp_f := 25;
        ELSIF x =- 9015 THEN
            exp_f := 25;
        ELSIF x =- 9014 THEN
            exp_f := 25;
        ELSIF x =- 9013 THEN
            exp_f := 25;
        ELSIF x =- 9012 THEN
            exp_f := 25;
        ELSIF x =- 9011 THEN
            exp_f := 26;
        ELSIF x =- 9010 THEN
            exp_f := 26;
        ELSIF x =- 9009 THEN
            exp_f := 26;
        ELSIF x =- 9008 THEN
            exp_f := 26;
        ELSIF x =- 9007 THEN
            exp_f := 26;
        ELSIF x =- 9006 THEN
            exp_f := 26;
        ELSIF x =- 9005 THEN
            exp_f := 26;
        ELSIF x =- 9004 THEN
            exp_f := 26;
        ELSIF x =- 9003 THEN
            exp_f := 26;
        ELSIF x =- 9002 THEN
            exp_f := 26;
        ELSIF x =- 9001 THEN
            exp_f := 26;
        ELSIF x =- 9000 THEN
            exp_f := 26;
        ELSIF x =- 8999 THEN
            exp_f := 26;
        ELSIF x =- 8998 THEN
            exp_f := 26;
        ELSIF x =- 8997 THEN
            exp_f := 26;
        ELSIF x =- 8996 THEN
            exp_f := 26;
        ELSIF x =- 8995 THEN
            exp_f := 26;
        ELSIF x =- 8994 THEN
            exp_f := 26;
        ELSIF x =- 8993 THEN
            exp_f := 26;
        ELSIF x =- 8992 THEN
            exp_f := 26;
        ELSIF x =- 8991 THEN
            exp_f := 26;
        ELSIF x =- 8990 THEN
            exp_f := 26;
        ELSIF x =- 8989 THEN
            exp_f := 26;
        ELSIF x =- 8988 THEN
            exp_f := 26;
        ELSIF x =- 8987 THEN
            exp_f := 26;
        ELSIF x =- 8986 THEN
            exp_f := 26;
        ELSIF x =- 8985 THEN
            exp_f := 26;
        ELSIF x =- 8984 THEN
            exp_f := 26;
        ELSIF x =- 8983 THEN
            exp_f := 26;
        ELSIF x =- 8982 THEN
            exp_f := 26;
        ELSIF x =- 8981 THEN
            exp_f := 26;
        ELSIF x =- 8980 THEN
            exp_f := 26;
        ELSIF x =- 8979 THEN
            exp_f := 26;
        ELSIF x =- 8978 THEN
            exp_f := 26;
        ELSIF x =- 8977 THEN
            exp_f := 26;
        ELSIF x =- 8976 THEN
            exp_f := 26;
        ELSIF x =- 8975 THEN
            exp_f := 26;
        ELSIF x =- 8974 THEN
            exp_f := 26;
        ELSIF x =- 8973 THEN
            exp_f := 26;
        ELSIF x =- 8972 THEN
            exp_f := 26;
        ELSIF x =- 8971 THEN
            exp_f := 26;
        ELSIF x =- 8970 THEN
            exp_f := 26;
        ELSIF x =- 8969 THEN
            exp_f := 26;
        ELSIF x =- 8968 THEN
            exp_f := 26;
        ELSIF x =- 8967 THEN
            exp_f := 26;
        ELSIF x =- 8966 THEN
            exp_f := 26;
        ELSIF x =- 8965 THEN
            exp_f := 26;
        ELSIF x =- 8964 THEN
            exp_f := 26;
        ELSIF x =- 8963 THEN
            exp_f := 26;
        ELSIF x =- 8962 THEN
            exp_f := 26;
        ELSIF x =- 8961 THEN
            exp_f := 26;
        ELSIF x =- 8960 THEN
            exp_f := 26;
        ELSIF x =- 8959 THEN
            exp_f := 26;
        ELSIF x =- 8958 THEN
            exp_f := 26;
        ELSIF x =- 8957 THEN
            exp_f := 26;
        ELSIF x =- 8956 THEN
            exp_f := 26;
        ELSIF x =- 8955 THEN
            exp_f := 26;
        ELSIF x =- 8954 THEN
            exp_f := 26;
        ELSIF x =- 8953 THEN
            exp_f := 26;
        ELSIF x =- 8952 THEN
            exp_f := 26;
        ELSIF x =- 8951 THEN
            exp_f := 26;
        ELSIF x =- 8950 THEN
            exp_f := 26;
        ELSIF x =- 8949 THEN
            exp_f := 26;
        ELSIF x =- 8948 THEN
            exp_f := 26;
        ELSIF x =- 8947 THEN
            exp_f := 26;
        ELSIF x =- 8946 THEN
            exp_f := 26;
        ELSIF x =- 8945 THEN
            exp_f := 26;
        ELSIF x =- 8944 THEN
            exp_f := 26;
        ELSIF x =- 8943 THEN
            exp_f := 26;
        ELSIF x =- 8942 THEN
            exp_f := 26;
        ELSIF x =- 8941 THEN
            exp_f := 26;
        ELSIF x =- 8940 THEN
            exp_f := 26;
        ELSIF x =- 8939 THEN
            exp_f := 26;
        ELSIF x =- 8938 THEN
            exp_f := 26;
        ELSIF x =- 8937 THEN
            exp_f := 26;
        ELSIF x =- 8936 THEN
            exp_f := 26;
        ELSIF x =- 8935 THEN
            exp_f := 26;
        ELSIF x =- 8934 THEN
            exp_f := 26;
        ELSIF x =- 8933 THEN
            exp_f := 26;
        ELSIF x =- 8932 THEN
            exp_f := 26;
        ELSIF x =- 8931 THEN
            exp_f := 26;
        ELSIF x =- 8930 THEN
            exp_f := 26;
        ELSIF x =- 8929 THEN
            exp_f := 27;
        ELSIF x =- 8928 THEN
            exp_f := 27;
        ELSIF x =- 8927 THEN
            exp_f := 27;
        ELSIF x =- 8926 THEN
            exp_f := 27;
        ELSIF x =- 8925 THEN
            exp_f := 27;
        ELSIF x =- 8924 THEN
            exp_f := 27;
        ELSIF x =- 8923 THEN
            exp_f := 27;
        ELSIF x =- 8922 THEN
            exp_f := 27;
        ELSIF x =- 8921 THEN
            exp_f := 27;
        ELSIF x =- 8920 THEN
            exp_f := 27;
        ELSIF x =- 8919 THEN
            exp_f := 27;
        ELSIF x =- 8918 THEN
            exp_f := 27;
        ELSIF x =- 8917 THEN
            exp_f := 27;
        ELSIF x =- 8916 THEN
            exp_f := 27;
        ELSIF x =- 8915 THEN
            exp_f := 27;
        ELSIF x =- 8914 THEN
            exp_f := 27;
        ELSIF x =- 8913 THEN
            exp_f := 27;
        ELSIF x =- 8912 THEN
            exp_f := 27;
        ELSIF x =- 8911 THEN
            exp_f := 27;
        ELSIF x =- 8910 THEN
            exp_f := 27;
        ELSIF x =- 8909 THEN
            exp_f := 27;
        ELSIF x =- 8908 THEN
            exp_f := 27;
        ELSIF x =- 8907 THEN
            exp_f := 27;
        ELSIF x =- 8906 THEN
            exp_f := 27;
        ELSIF x =- 8905 THEN
            exp_f := 27;
        ELSIF x =- 8904 THEN
            exp_f := 27;
        ELSIF x =- 8903 THEN
            exp_f := 27;
        ELSIF x =- 8902 THEN
            exp_f := 27;
        ELSIF x =- 8901 THEN
            exp_f := 27;
        ELSIF x =- 8900 THEN
            exp_f := 27;
        ELSIF x =- 8899 THEN
            exp_f := 27;
        ELSIF x =- 8898 THEN
            exp_f := 27;
        ELSIF x =- 8897 THEN
            exp_f := 27;
        ELSIF x =- 8896 THEN
            exp_f := 27;
        ELSIF x =- 8895 THEN
            exp_f := 27;
        ELSIF x =- 8894 THEN
            exp_f := 27;
        ELSIF x =- 8893 THEN
            exp_f := 27;
        ELSIF x =- 8892 THEN
            exp_f := 27;
        ELSIF x =- 8891 THEN
            exp_f := 27;
        ELSIF x =- 8890 THEN
            exp_f := 27;
        ELSIF x =- 8889 THEN
            exp_f := 27;
        ELSIF x =- 8888 THEN
            exp_f := 27;
        ELSIF x =- 8887 THEN
            exp_f := 27;
        ELSIF x =- 8886 THEN
            exp_f := 27;
        ELSIF x =- 8885 THEN
            exp_f := 27;
        ELSIF x =- 8884 THEN
            exp_f := 27;
        ELSIF x =- 8883 THEN
            exp_f := 27;
        ELSIF x =- 8882 THEN
            exp_f := 27;
        ELSIF x =- 8881 THEN
            exp_f := 27;
        ELSIF x =- 8880 THEN
            exp_f := 27;
        ELSIF x =- 8879 THEN
            exp_f := 27;
        ELSIF x =- 8878 THEN
            exp_f := 27;
        ELSIF x =- 8877 THEN
            exp_f := 27;
        ELSIF x =- 8876 THEN
            exp_f := 27;
        ELSIF x =- 8875 THEN
            exp_f := 27;
        ELSIF x =- 8874 THEN
            exp_f := 27;
        ELSIF x =- 8873 THEN
            exp_f := 27;
        ELSIF x =- 8872 THEN
            exp_f := 27;
        ELSIF x =- 8871 THEN
            exp_f := 27;
        ELSIF x =- 8870 THEN
            exp_f := 27;
        ELSIF x =- 8869 THEN
            exp_f := 27;
        ELSIF x =- 8868 THEN
            exp_f := 27;
        ELSIF x =- 8867 THEN
            exp_f := 27;
        ELSIF x =- 8866 THEN
            exp_f := 27;
        ELSIF x =- 8865 THEN
            exp_f := 27;
        ELSIF x =- 8864 THEN
            exp_f := 27;
        ELSIF x =- 8863 THEN
            exp_f := 27;
        ELSIF x =- 8862 THEN
            exp_f := 27;
        ELSIF x =- 8861 THEN
            exp_f := 27;
        ELSIF x =- 8860 THEN
            exp_f := 27;
        ELSIF x =- 8859 THEN
            exp_f := 27;
        ELSIF x =- 8858 THEN
            exp_f := 27;
        ELSIF x =- 8857 THEN
            exp_f := 27;
        ELSIF x =- 8856 THEN
            exp_f := 27;
        ELSIF x =- 8855 THEN
            exp_f := 27;
        ELSIF x =- 8854 THEN
            exp_f := 27;
        ELSIF x =- 8853 THEN
            exp_f := 27;
        ELSIF x =- 8852 THEN
            exp_f := 27;
        ELSIF x =- 8851 THEN
            exp_f := 27;
        ELSIF x =- 8850 THEN
            exp_f := 27;
        ELSIF x =- 8849 THEN
            exp_f := 27;
        ELSIF x =- 8848 THEN
            exp_f := 27;
        ELSIF x =- 8847 THEN
            exp_f := 28;
        ELSIF x =- 8846 THEN
            exp_f := 28;
        ELSIF x =- 8845 THEN
            exp_f := 28;
        ELSIF x =- 8844 THEN
            exp_f := 28;
        ELSIF x =- 8843 THEN
            exp_f := 28;
        ELSIF x =- 8842 THEN
            exp_f := 28;
        ELSIF x =- 8841 THEN
            exp_f := 28;
        ELSIF x =- 8840 THEN
            exp_f := 28;
        ELSIF x =- 8839 THEN
            exp_f := 28;
        ELSIF x =- 8838 THEN
            exp_f := 28;
        ELSIF x =- 8837 THEN
            exp_f := 28;
        ELSIF x =- 8836 THEN
            exp_f := 28;
        ELSIF x =- 8835 THEN
            exp_f := 28;
        ELSIF x =- 8834 THEN
            exp_f := 28;
        ELSIF x =- 8833 THEN
            exp_f := 28;
        ELSIF x =- 8832 THEN
            exp_f := 28;
        ELSIF x =- 8831 THEN
            exp_f := 28;
        ELSIF x =- 8830 THEN
            exp_f := 28;
        ELSIF x =- 8829 THEN
            exp_f := 28;
        ELSIF x =- 8828 THEN
            exp_f := 28;
        ELSIF x =- 8827 THEN
            exp_f := 28;
        ELSIF x =- 8826 THEN
            exp_f := 28;
        ELSIF x =- 8825 THEN
            exp_f := 28;
        ELSIF x =- 8824 THEN
            exp_f := 28;
        ELSIF x =- 8823 THEN
            exp_f := 28;
        ELSIF x =- 8822 THEN
            exp_f := 28;
        ELSIF x =- 8821 THEN
            exp_f := 28;
        ELSIF x =- 8820 THEN
            exp_f := 28;
        ELSIF x =- 8819 THEN
            exp_f := 28;
        ELSIF x =- 8818 THEN
            exp_f := 28;
        ELSIF x =- 8817 THEN
            exp_f := 28;
        ELSIF x =- 8816 THEN
            exp_f := 28;
        ELSIF x =- 8815 THEN
            exp_f := 28;
        ELSIF x =- 8814 THEN
            exp_f := 28;
        ELSIF x =- 8813 THEN
            exp_f := 28;
        ELSIF x =- 8812 THEN
            exp_f := 28;
        ELSIF x =- 8811 THEN
            exp_f := 28;
        ELSIF x =- 8810 THEN
            exp_f := 28;
        ELSIF x =- 8809 THEN
            exp_f := 28;
        ELSIF x =- 8808 THEN
            exp_f := 28;
        ELSIF x =- 8807 THEN
            exp_f := 28;
        ELSIF x =- 8806 THEN
            exp_f := 28;
        ELSIF x =- 8805 THEN
            exp_f := 28;
        ELSIF x =- 8804 THEN
            exp_f := 28;
        ELSIF x =- 8803 THEN
            exp_f := 28;
        ELSIF x =- 8802 THEN
            exp_f := 28;
        ELSIF x =- 8801 THEN
            exp_f := 28;
        ELSIF x =- 8800 THEN
            exp_f := 28;
        ELSIF x =- 8799 THEN
            exp_f := 28;
        ELSIF x =- 8798 THEN
            exp_f := 28;
        ELSIF x =- 8797 THEN
            exp_f := 28;
        ELSIF x =- 8796 THEN
            exp_f := 28;
        ELSIF x =- 8795 THEN
            exp_f := 28;
        ELSIF x =- 8794 THEN
            exp_f := 28;
        ELSIF x =- 8793 THEN
            exp_f := 28;
        ELSIF x =- 8792 THEN
            exp_f := 28;
        ELSIF x =- 8791 THEN
            exp_f := 28;
        ELSIF x =- 8790 THEN
            exp_f := 28;
        ELSIF x =- 8789 THEN
            exp_f := 28;
        ELSIF x =- 8788 THEN
            exp_f := 28;
        ELSIF x =- 8787 THEN
            exp_f := 28;
        ELSIF x =- 8786 THEN
            exp_f := 28;
        ELSIF x =- 8785 THEN
            exp_f := 28;
        ELSIF x =- 8784 THEN
            exp_f := 28;
        ELSIF x =- 8783 THEN
            exp_f := 28;
        ELSIF x =- 8782 THEN
            exp_f := 28;
        ELSIF x =- 8781 THEN
            exp_f := 28;
        ELSIF x =- 8780 THEN
            exp_f := 28;
        ELSIF x =- 8779 THEN
            exp_f := 28;
        ELSIF x =- 8778 THEN
            exp_f := 28;
        ELSIF x =- 8777 THEN
            exp_f := 28;
        ELSIF x =- 8776 THEN
            exp_f := 28;
        ELSIF x =- 8775 THEN
            exp_f := 28;
        ELSIF x =- 8774 THEN
            exp_f := 28;
        ELSIF x =- 8773 THEN
            exp_f := 28;
        ELSIF x =- 8772 THEN
            exp_f := 28;
        ELSIF x =- 8771 THEN
            exp_f := 28;
        ELSIF x =- 8770 THEN
            exp_f := 28;
        ELSIF x =- 8769 THEN
            exp_f := 28;
        ELSIF x =- 8768 THEN
            exp_f := 28;
        ELSIF x =- 8767 THEN
            exp_f := 28;
        ELSIF x =- 8766 THEN
            exp_f := 28;
        ELSIF x =- 8765 THEN
            exp_f := 29;
        ELSIF x =- 8764 THEN
            exp_f := 29;
        ELSIF x =- 8763 THEN
            exp_f := 29;
        ELSIF x =- 8762 THEN
            exp_f := 29;
        ELSIF x =- 8761 THEN
            exp_f := 29;
        ELSIF x =- 8760 THEN
            exp_f := 29;
        ELSIF x =- 8759 THEN
            exp_f := 29;
        ELSIF x =- 8758 THEN
            exp_f := 29;
        ELSIF x =- 8757 THEN
            exp_f := 29;
        ELSIF x =- 8756 THEN
            exp_f := 29;
        ELSIF x =- 8755 THEN
            exp_f := 29;
        ELSIF x =- 8754 THEN
            exp_f := 29;
        ELSIF x =- 8753 THEN
            exp_f := 29;
        ELSIF x =- 8752 THEN
            exp_f := 29;
        ELSIF x =- 8751 THEN
            exp_f := 29;
        ELSIF x =- 8750 THEN
            exp_f := 29;
        ELSIF x =- 8749 THEN
            exp_f := 29;
        ELSIF x =- 8748 THEN
            exp_f := 29;
        ELSIF x =- 8747 THEN
            exp_f := 29;
        ELSIF x =- 8746 THEN
            exp_f := 29;
        ELSIF x =- 8745 THEN
            exp_f := 29;
        ELSIF x =- 8744 THEN
            exp_f := 29;
        ELSIF x =- 8743 THEN
            exp_f := 29;
        ELSIF x =- 8742 THEN
            exp_f := 29;
        ELSIF x =- 8741 THEN
            exp_f := 29;
        ELSIF x =- 8740 THEN
            exp_f := 29;
        ELSIF x =- 8739 THEN
            exp_f := 29;
        ELSIF x =- 8738 THEN
            exp_f := 29;
        ELSIF x =- 8737 THEN
            exp_f := 29;
        ELSIF x =- 8736 THEN
            exp_f := 29;
        ELSIF x =- 8735 THEN
            exp_f := 29;
        ELSIF x =- 8734 THEN
            exp_f := 29;
        ELSIF x =- 8733 THEN
            exp_f := 29;
        ELSIF x =- 8732 THEN
            exp_f := 29;
        ELSIF x =- 8731 THEN
            exp_f := 29;
        ELSIF x =- 8730 THEN
            exp_f := 29;
        ELSIF x =- 8729 THEN
            exp_f := 29;
        ELSIF x =- 8728 THEN
            exp_f := 29;
        ELSIF x =- 8727 THEN
            exp_f := 29;
        ELSIF x =- 8726 THEN
            exp_f := 29;
        ELSIF x =- 8725 THEN
            exp_f := 29;
        ELSIF x =- 8724 THEN
            exp_f := 29;
        ELSIF x =- 8723 THEN
            exp_f := 29;
        ELSIF x =- 8722 THEN
            exp_f := 29;
        ELSIF x =- 8721 THEN
            exp_f := 29;
        ELSIF x =- 8720 THEN
            exp_f := 29;
        ELSIF x =- 8719 THEN
            exp_f := 29;
        ELSIF x =- 8718 THEN
            exp_f := 29;
        ELSIF x =- 8717 THEN
            exp_f := 29;
        ELSIF x =- 8716 THEN
            exp_f := 29;
        ELSIF x =- 8715 THEN
            exp_f := 29;
        ELSIF x =- 8714 THEN
            exp_f := 29;
        ELSIF x =- 8713 THEN
            exp_f := 29;
        ELSIF x =- 8712 THEN
            exp_f := 29;
        ELSIF x =- 8711 THEN
            exp_f := 29;
        ELSIF x =- 8710 THEN
            exp_f := 29;
        ELSIF x =- 8709 THEN
            exp_f := 29;
        ELSIF x =- 8708 THEN
            exp_f := 29;
        ELSIF x =- 8707 THEN
            exp_f := 29;
        ELSIF x =- 8706 THEN
            exp_f := 29;
        ELSIF x =- 8705 THEN
            exp_f := 29;
        ELSIF x =- 8704 THEN
            exp_f := 29;
        ELSIF x =- 8703 THEN
            exp_f := 29;
        ELSIF x =- 8702 THEN
            exp_f := 29;
        ELSIF x =- 8701 THEN
            exp_f := 29;
        ELSIF x =- 8700 THEN
            exp_f := 29;
        ELSIF x =- 8699 THEN
            exp_f := 29;
        ELSIF x =- 8698 THEN
            exp_f := 29;
        ELSIF x =- 8697 THEN
            exp_f := 29;
        ELSIF x =- 8696 THEN
            exp_f := 29;
        ELSIF x =- 8695 THEN
            exp_f := 29;
        ELSIF x =- 8694 THEN
            exp_f := 29;
        ELSIF x =- 8693 THEN
            exp_f := 29;
        ELSIF x =- 8692 THEN
            exp_f := 29;
        ELSIF x =- 8691 THEN
            exp_f := 29;
        ELSIF x =- 8690 THEN
            exp_f := 29;
        ELSIF x =- 8689 THEN
            exp_f := 29;
        ELSIF x =- 8688 THEN
            exp_f := 29;
        ELSIF x =- 8687 THEN
            exp_f := 29;
        ELSIF x =- 8686 THEN
            exp_f := 29;
        ELSIF x =- 8685 THEN
            exp_f := 29;
        ELSIF x =- 8684 THEN
            exp_f := 29;
        ELSIF x =- 8683 THEN
            exp_f := 29;
        ELSIF x =- 8682 THEN
            exp_f := 29;
        ELSIF x =- 8681 THEN
            exp_f := 29;
        ELSIF x =- 8680 THEN
            exp_f := 29;
        ELSIF x =- 8679 THEN
            exp_f := 29;
        ELSIF x =- 8678 THEN
            exp_f := 29;
        ELSIF x =- 8677 THEN
            exp_f := 29;
        ELSIF x =- 8676 THEN
            exp_f := 29;
        ELSIF x =- 8675 THEN
            exp_f := 29;
        ELSIF x =- 8674 THEN
            exp_f := 29;
        ELSIF x =- 8673 THEN
            exp_f := 30;
        ELSIF x =- 8672 THEN
            exp_f := 30;
        ELSIF x =- 8671 THEN
            exp_f := 30;
        ELSIF x =- 8670 THEN
            exp_f := 30;
        ELSIF x =- 8669 THEN
            exp_f := 30;
        ELSIF x =- 8668 THEN
            exp_f := 30;
        ELSIF x =- 8667 THEN
            exp_f := 30;
        ELSIF x =- 8666 THEN
            exp_f := 30;
        ELSIF x =- 8665 THEN
            exp_f := 30;
        ELSIF x =- 8664 THEN
            exp_f := 30;
        ELSIF x =- 8663 THEN
            exp_f := 30;
        ELSIF x =- 8662 THEN
            exp_f := 30;
        ELSIF x =- 8661 THEN
            exp_f := 30;
        ELSIF x =- 8660 THEN
            exp_f := 30;
        ELSIF x =- 8659 THEN
            exp_f := 30;
        ELSIF x =- 8658 THEN
            exp_f := 30;
        ELSIF x =- 8657 THEN
            exp_f := 30;
        ELSIF x =- 8656 THEN
            exp_f := 30;
        ELSIF x =- 8655 THEN
            exp_f := 30;
        ELSIF x =- 8654 THEN
            exp_f := 30;
        ELSIF x =- 8653 THEN
            exp_f := 30;
        ELSIF x =- 8652 THEN
            exp_f := 30;
        ELSIF x =- 8651 THEN
            exp_f := 30;
        ELSIF x =- 8650 THEN
            exp_f := 30;
        ELSIF x =- 8649 THEN
            exp_f := 30;
        ELSIF x =- 8648 THEN
            exp_f := 30;
        ELSIF x =- 8647 THEN
            exp_f := 30;
        ELSIF x =- 8646 THEN
            exp_f := 30;
        ELSIF x =- 8645 THEN
            exp_f := 30;
        ELSIF x =- 8644 THEN
            exp_f := 30;
        ELSIF x =- 8643 THEN
            exp_f := 30;
        ELSIF x =- 8642 THEN
            exp_f := 30;
        ELSIF x =- 8641 THEN
            exp_f := 30;
        ELSIF x =- 8640 THEN
            exp_f := 30;
        ELSIF x =- 8639 THEN
            exp_f := 30;
        ELSIF x =- 8638 THEN
            exp_f := 30;
        ELSIF x =- 8637 THEN
            exp_f := 30;
        ELSIF x =- 8636 THEN
            exp_f := 30;
        ELSIF x =- 8635 THEN
            exp_f := 30;
        ELSIF x =- 8634 THEN
            exp_f := 30;
        ELSIF x =- 8633 THEN
            exp_f := 30;
        ELSIF x =- 8632 THEN
            exp_f := 30;
        ELSIF x =- 8631 THEN
            exp_f := 30;
        ELSIF x =- 8630 THEN
            exp_f := 30;
        ELSIF x =- 8629 THEN
            exp_f := 30;
        ELSIF x =- 8628 THEN
            exp_f := 30;
        ELSIF x =- 8627 THEN
            exp_f := 30;
        ELSIF x =- 8626 THEN
            exp_f := 30;
        ELSIF x =- 8625 THEN
            exp_f := 30;
        ELSIF x =- 8624 THEN
            exp_f := 30;
        ELSIF x =- 8623 THEN
            exp_f := 30;
        ELSIF x =- 8622 THEN
            exp_f := 30;
        ELSIF x =- 8621 THEN
            exp_f := 30;
        ELSIF x =- 8620 THEN
            exp_f := 30;
        ELSIF x =- 8619 THEN
            exp_f := 30;
        ELSIF x =- 8618 THEN
            exp_f := 30;
        ELSIF x =- 8617 THEN
            exp_f := 30;
        ELSIF x =- 8616 THEN
            exp_f := 30;
        ELSIF x =- 8615 THEN
            exp_f := 30;
        ELSIF x =- 8614 THEN
            exp_f := 30;
        ELSIF x =- 8613 THEN
            exp_f := 31;
        ELSIF x =- 8612 THEN
            exp_f := 31;
        ELSIF x =- 8611 THEN
            exp_f := 31;
        ELSIF x =- 8610 THEN
            exp_f := 31;
        ELSIF x =- 8609 THEN
            exp_f := 31;
        ELSIF x =- 8608 THEN
            exp_f := 31;
        ELSIF x =- 8607 THEN
            exp_f := 31;
        ELSIF x =- 8606 THEN
            exp_f := 31;
        ELSIF x =- 8605 THEN
            exp_f := 31;
        ELSIF x =- 8604 THEN
            exp_f := 31;
        ELSIF x =- 8603 THEN
            exp_f := 31;
        ELSIF x =- 8602 THEN
            exp_f := 31;
        ELSIF x =- 8601 THEN
            exp_f := 31;
        ELSIF x =- 8600 THEN
            exp_f := 31;
        ELSIF x =- 8599 THEN
            exp_f := 31;
        ELSIF x =- 8598 THEN
            exp_f := 31;
        ELSIF x =- 8597 THEN
            exp_f := 31;
        ELSIF x =- 8596 THEN
            exp_f := 31;
        ELSIF x =- 8595 THEN
            exp_f := 31;
        ELSIF x =- 8594 THEN
            exp_f := 31;
        ELSIF x =- 8593 THEN
            exp_f := 31;
        ELSIF x =- 8592 THEN
            exp_f := 31;
        ELSIF x =- 8591 THEN
            exp_f := 31;
        ELSIF x =- 8590 THEN
            exp_f := 31;
        ELSIF x =- 8589 THEN
            exp_f := 31;
        ELSIF x =- 8588 THEN
            exp_f := 31;
        ELSIF x =- 8587 THEN
            exp_f := 31;
        ELSIF x =- 8586 THEN
            exp_f := 31;
        ELSIF x =- 8585 THEN
            exp_f := 31;
        ELSIF x =- 8584 THEN
            exp_f := 31;
        ELSIF x =- 8583 THEN
            exp_f := 31;
        ELSIF x =- 8582 THEN
            exp_f := 31;
        ELSIF x =- 8581 THEN
            exp_f := 31;
        ELSIF x =- 8580 THEN
            exp_f := 31;
        ELSIF x =- 8579 THEN
            exp_f := 31;
        ELSIF x =- 8578 THEN
            exp_f := 31;
        ELSIF x =- 8577 THEN
            exp_f := 31;
        ELSIF x =- 8576 THEN
            exp_f := 31;
        ELSIF x =- 8575 THEN
            exp_f := 31;
        ELSIF x =- 8574 THEN
            exp_f := 31;
        ELSIF x =- 8573 THEN
            exp_f := 31;
        ELSIF x =- 8572 THEN
            exp_f := 31;
        ELSIF x =- 8571 THEN
            exp_f := 31;
        ELSIF x =- 8570 THEN
            exp_f := 31;
        ELSIF x =- 8569 THEN
            exp_f := 31;
        ELSIF x =- 8568 THEN
            exp_f := 31;
        ELSIF x =- 8567 THEN
            exp_f := 31;
        ELSIF x =- 8566 THEN
            exp_f := 31;
        ELSIF x =- 8565 THEN
            exp_f := 31;
        ELSIF x =- 8564 THEN
            exp_f := 31;
        ELSIF x =- 8563 THEN
            exp_f := 31;
        ELSIF x =- 8562 THEN
            exp_f := 31;
        ELSIF x =- 8561 THEN
            exp_f := 31;
        ELSIF x =- 8560 THEN
            exp_f := 31;
        ELSIF x =- 8559 THEN
            exp_f := 31;
        ELSIF x =- 8558 THEN
            exp_f := 31;
        ELSIF x =- 8557 THEN
            exp_f := 31;
        ELSIF x =- 8556 THEN
            exp_f := 31;
        ELSIF x =- 8555 THEN
            exp_f := 31;
        ELSIF x =- 8554 THEN
            exp_f := 31;
        ELSIF x =- 8553 THEN
            exp_f := 32;
        ELSIF x =- 8552 THEN
            exp_f := 32;
        ELSIF x =- 8551 THEN
            exp_f := 32;
        ELSIF x =- 8550 THEN
            exp_f := 32;
        ELSIF x =- 8549 THEN
            exp_f := 32;
        ELSIF x =- 8548 THEN
            exp_f := 32;
        ELSIF x =- 8547 THEN
            exp_f := 32;
        ELSIF x =- 8546 THEN
            exp_f := 32;
        ELSIF x =- 8545 THEN
            exp_f := 32;
        ELSIF x =- 8544 THEN
            exp_f := 32;
        ELSIF x =- 8543 THEN
            exp_f := 32;
        ELSIF x =- 8542 THEN
            exp_f := 32;
        ELSIF x =- 8541 THEN
            exp_f := 32;
        ELSIF x =- 8540 THEN
            exp_f := 32;
        ELSIF x =- 8539 THEN
            exp_f := 32;
        ELSIF x =- 8538 THEN
            exp_f := 32;
        ELSIF x =- 8537 THEN
            exp_f := 32;
        ELSIF x =- 8536 THEN
            exp_f := 32;
        ELSIF x =- 8535 THEN
            exp_f := 32;
        ELSIF x =- 8534 THEN
            exp_f := 32;
        ELSIF x =- 8533 THEN
            exp_f := 32;
        ELSIF x =- 8532 THEN
            exp_f := 32;
        ELSIF x =- 8531 THEN
            exp_f := 32;
        ELSIF x =- 8530 THEN
            exp_f := 32;
        ELSIF x =- 8529 THEN
            exp_f := 32;
        ELSIF x =- 8528 THEN
            exp_f := 32;
        ELSIF x =- 8527 THEN
            exp_f := 32;
        ELSIF x =- 8526 THEN
            exp_f := 32;
        ELSIF x =- 8525 THEN
            exp_f := 32;
        ELSIF x =- 8524 THEN
            exp_f := 32;
        ELSIF x =- 8523 THEN
            exp_f := 32;
        ELSIF x =- 8522 THEN
            exp_f := 32;
        ELSIF x =- 8521 THEN
            exp_f := 32;
        ELSIF x =- 8520 THEN
            exp_f := 32;
        ELSIF x =- 8519 THEN
            exp_f := 32;
        ELSIF x =- 8518 THEN
            exp_f := 32;
        ELSIF x =- 8517 THEN
            exp_f := 32;
        ELSIF x =- 8516 THEN
            exp_f := 32;
        ELSIF x =- 8515 THEN
            exp_f := 32;
        ELSIF x =- 8514 THEN
            exp_f := 32;
        ELSIF x =- 8513 THEN
            exp_f := 32;
        ELSIF x =- 8512 THEN
            exp_f := 32;
        ELSIF x =- 8511 THEN
            exp_f := 32;
        ELSIF x =- 8510 THEN
            exp_f := 32;
        ELSIF x =- 8509 THEN
            exp_f := 32;
        ELSIF x =- 8508 THEN
            exp_f := 32;
        ELSIF x =- 8507 THEN
            exp_f := 32;
        ELSIF x =- 8506 THEN
            exp_f := 32;
        ELSIF x =- 8505 THEN
            exp_f := 32;
        ELSIF x =- 8504 THEN
            exp_f := 32;
        ELSIF x =- 8503 THEN
            exp_f := 32;
        ELSIF x =- 8502 THEN
            exp_f := 32;
        ELSIF x =- 8501 THEN
            exp_f := 32;
        ELSIF x =- 8500 THEN
            exp_f := 32;
        ELSIF x =- 8499 THEN
            exp_f := 32;
        ELSIF x =- 8498 THEN
            exp_f := 32;
        ELSIF x =- 8497 THEN
            exp_f := 32;
        ELSIF x =- 8496 THEN
            exp_f := 32;
        ELSIF x =- 8495 THEN
            exp_f := 32;
        ELSIF x =- 8494 THEN
            exp_f := 32;
        ELSIF x =- 8493 THEN
            exp_f := 33;
        ELSIF x =- 8492 THEN
            exp_f := 33;
        ELSIF x =- 8491 THEN
            exp_f := 33;
        ELSIF x =- 8490 THEN
            exp_f := 33;
        ELSIF x =- 8489 THEN
            exp_f := 33;
        ELSIF x =- 8488 THEN
            exp_f := 33;
        ELSIF x =- 8487 THEN
            exp_f := 33;
        ELSIF x =- 8486 THEN
            exp_f := 33;
        ELSIF x =- 8485 THEN
            exp_f := 33;
        ELSIF x =- 8484 THEN
            exp_f := 33;
        ELSIF x =- 8483 THEN
            exp_f := 33;
        ELSIF x =- 8482 THEN
            exp_f := 33;
        ELSIF x =- 8481 THEN
            exp_f := 33;
        ELSIF x =- 8480 THEN
            exp_f := 33;
        ELSIF x =- 8479 THEN
            exp_f := 33;
        ELSIF x =- 8478 THEN
            exp_f := 33;
        ELSIF x =- 8477 THEN
            exp_f := 33;
        ELSIF x =- 8476 THEN
            exp_f := 33;
        ELSIF x =- 8475 THEN
            exp_f := 33;
        ELSIF x =- 8474 THEN
            exp_f := 33;
        ELSIF x =- 8473 THEN
            exp_f := 33;
        ELSIF x =- 8472 THEN
            exp_f := 33;
        ELSIF x =- 8471 THEN
            exp_f := 33;
        ELSIF x =- 8470 THEN
            exp_f := 33;
        ELSIF x =- 8469 THEN
            exp_f := 33;
        ELSIF x =- 8468 THEN
            exp_f := 33;
        ELSIF x =- 8467 THEN
            exp_f := 33;
        ELSIF x =- 8466 THEN
            exp_f := 33;
        ELSIF x =- 8465 THEN
            exp_f := 33;
        ELSIF x =- 8464 THEN
            exp_f := 33;
        ELSIF x =- 8463 THEN
            exp_f := 33;
        ELSIF x =- 8462 THEN
            exp_f := 33;
        ELSIF x =- 8461 THEN
            exp_f := 33;
        ELSIF x =- 8460 THEN
            exp_f := 33;
        ELSIF x =- 8459 THEN
            exp_f := 33;
        ELSIF x =- 8458 THEN
            exp_f := 33;
        ELSIF x =- 8457 THEN
            exp_f := 33;
        ELSIF x =- 8456 THEN
            exp_f := 33;
        ELSIF x =- 8455 THEN
            exp_f := 33;
        ELSIF x =- 8454 THEN
            exp_f := 33;
        ELSIF x =- 8453 THEN
            exp_f := 33;
        ELSIF x =- 8452 THEN
            exp_f := 33;
        ELSIF x =- 8451 THEN
            exp_f := 33;
        ELSIF x =- 8450 THEN
            exp_f := 33;
        ELSIF x =- 8449 THEN
            exp_f := 33;
        ELSIF x =- 8448 THEN
            exp_f := 33;
        ELSIF x =- 8447 THEN
            exp_f := 33;
        ELSIF x =- 8446 THEN
            exp_f := 33;
        ELSIF x =- 8445 THEN
            exp_f := 33;
        ELSIF x =- 8444 THEN
            exp_f := 33;
        ELSIF x =- 8443 THEN
            exp_f := 33;
        ELSIF x =- 8442 THEN
            exp_f := 33;
        ELSIF x =- 8441 THEN
            exp_f := 33;
        ELSIF x =- 8440 THEN
            exp_f := 33;
        ELSIF x =- 8439 THEN
            exp_f := 33;
        ELSIF x =- 8438 THEN
            exp_f := 33;
        ELSIF x =- 8437 THEN
            exp_f := 33;
        ELSIF x =- 8436 THEN
            exp_f := 33;
        ELSIF x =- 8435 THEN
            exp_f := 33;
        ELSIF x =- 8434 THEN
            exp_f := 33;
        ELSIF x =- 8433 THEN
            exp_f := 33;
        ELSIF x =- 8432 THEN
            exp_f := 34;
        ELSIF x =- 8431 THEN
            exp_f := 34;
        ELSIF x =- 8430 THEN
            exp_f := 34;
        ELSIF x =- 8429 THEN
            exp_f := 34;
        ELSIF x =- 8428 THEN
            exp_f := 34;
        ELSIF x =- 8427 THEN
            exp_f := 34;
        ELSIF x =- 8426 THEN
            exp_f := 34;
        ELSIF x =- 8425 THEN
            exp_f := 34;
        ELSIF x =- 8424 THEN
            exp_f := 34;
        ELSIF x =- 8423 THEN
            exp_f := 34;
        ELSIF x =- 8422 THEN
            exp_f := 34;
        ELSIF x =- 8421 THEN
            exp_f := 34;
        ELSIF x =- 8420 THEN
            exp_f := 34;
        ELSIF x =- 8419 THEN
            exp_f := 34;
        ELSIF x =- 8418 THEN
            exp_f := 34;
        ELSIF x =- 8417 THEN
            exp_f := 34;
        ELSIF x =- 8416 THEN
            exp_f := 34;
        ELSIF x =- 8415 THEN
            exp_f := 34;
        ELSIF x =- 8414 THEN
            exp_f := 34;
        ELSIF x =- 8413 THEN
            exp_f := 34;
        ELSIF x =- 8412 THEN
            exp_f := 34;
        ELSIF x =- 8411 THEN
            exp_f := 34;
        ELSIF x =- 8410 THEN
            exp_f := 34;
        ELSIF x =- 8409 THEN
            exp_f := 34;
        ELSIF x =- 8408 THEN
            exp_f := 34;
        ELSIF x =- 8407 THEN
            exp_f := 34;
        ELSIF x =- 8406 THEN
            exp_f := 34;
        ELSIF x =- 8405 THEN
            exp_f := 34;
        ELSIF x =- 8404 THEN
            exp_f := 34;
        ELSIF x =- 8403 THEN
            exp_f := 34;
        ELSIF x =- 8402 THEN
            exp_f := 34;
        ELSIF x =- 8401 THEN
            exp_f := 34;
        ELSIF x =- 8400 THEN
            exp_f := 34;
        ELSIF x =- 8399 THEN
            exp_f := 34;
        ELSIF x =- 8398 THEN
            exp_f := 34;
        ELSIF x =- 8397 THEN
            exp_f := 34;
        ELSIF x =- 8396 THEN
            exp_f := 34;
        ELSIF x =- 8395 THEN
            exp_f := 34;
        ELSIF x =- 8394 THEN
            exp_f := 34;
        ELSIF x =- 8393 THEN
            exp_f := 34;
        ELSIF x =- 8392 THEN
            exp_f := 34;
        ELSIF x =- 8391 THEN
            exp_f := 34;
        ELSIF x =- 8390 THEN
            exp_f := 34;
        ELSIF x =- 8389 THEN
            exp_f := 34;
        ELSIF x =- 8388 THEN
            exp_f := 34;
        ELSIF x =- 8387 THEN
            exp_f := 34;
        ELSIF x =- 8386 THEN
            exp_f := 34;
        ELSIF x =- 8385 THEN
            exp_f := 34;
        ELSIF x =- 8384 THEN
            exp_f := 34;
        ELSIF x =- 8383 THEN
            exp_f := 34;
        ELSIF x =- 8382 THEN
            exp_f := 34;
        ELSIF x =- 8381 THEN
            exp_f := 34;
        ELSIF x =- 8380 THEN
            exp_f := 34;
        ELSIF x =- 8379 THEN
            exp_f := 34;
        ELSIF x =- 8378 THEN
            exp_f := 34;
        ELSIF x =- 8377 THEN
            exp_f := 34;
        ELSIF x =- 8376 THEN
            exp_f := 34;
        ELSIF x =- 8375 THEN
            exp_f := 34;
        ELSIF x =- 8374 THEN
            exp_f := 34;
        ELSIF x =- 8373 THEN
            exp_f := 34;
        ELSIF x =- 8372 THEN
            exp_f := 35;
        ELSIF x =- 8371 THEN
            exp_f := 35;
        ELSIF x =- 8370 THEN
            exp_f := 35;
        ELSIF x =- 8369 THEN
            exp_f := 35;
        ELSIF x =- 8368 THEN
            exp_f := 35;
        ELSIF x =- 8367 THEN
            exp_f := 35;
        ELSIF x =- 8366 THEN
            exp_f := 35;
        ELSIF x =- 8365 THEN
            exp_f := 35;
        ELSIF x =- 8364 THEN
            exp_f := 35;
        ELSIF x =- 8363 THEN
            exp_f := 35;
        ELSIF x =- 8362 THEN
            exp_f := 35;
        ELSIF x =- 8361 THEN
            exp_f := 35;
        ELSIF x =- 8360 THEN
            exp_f := 35;
        ELSIF x =- 8359 THEN
            exp_f := 35;
        ELSIF x =- 8358 THEN
            exp_f := 35;
        ELSIF x =- 8357 THEN
            exp_f := 35;
        ELSIF x =- 8356 THEN
            exp_f := 35;
        ELSIF x =- 8355 THEN
            exp_f := 35;
        ELSIF x =- 8354 THEN
            exp_f := 35;
        ELSIF x =- 8353 THEN
            exp_f := 35;
        ELSIF x =- 8352 THEN
            exp_f := 35;
        ELSIF x =- 8351 THEN
            exp_f := 35;
        ELSIF x =- 8350 THEN
            exp_f := 35;
        ELSIF x =- 8349 THEN
            exp_f := 35;
        ELSIF x =- 8348 THEN
            exp_f := 35;
        ELSIF x =- 8347 THEN
            exp_f := 35;
        ELSIF x =- 8346 THEN
            exp_f := 35;
        ELSIF x =- 8345 THEN
            exp_f := 35;
        ELSIF x =- 8344 THEN
            exp_f := 35;
        ELSIF x =- 8343 THEN
            exp_f := 35;
        ELSIF x =- 8342 THEN
            exp_f := 35;
        ELSIF x =- 8341 THEN
            exp_f := 35;
        ELSIF x =- 8340 THEN
            exp_f := 35;
        ELSIF x =- 8339 THEN
            exp_f := 35;
        ELSIF x =- 8338 THEN
            exp_f := 35;
        ELSIF x =- 8337 THEN
            exp_f := 35;
        ELSIF x =- 8336 THEN
            exp_f := 35;
        ELSIF x =- 8335 THEN
            exp_f := 35;
        ELSIF x =- 8334 THEN
            exp_f := 35;
        ELSIF x =- 8333 THEN
            exp_f := 35;
        ELSIF x =- 8332 THEN
            exp_f := 35;
        ELSIF x =- 8331 THEN
            exp_f := 35;
        ELSIF x =- 8330 THEN
            exp_f := 35;
        ELSIF x =- 8329 THEN
            exp_f := 35;
        ELSIF x =- 8328 THEN
            exp_f := 35;
        ELSIF x =- 8327 THEN
            exp_f := 35;
        ELSIF x =- 8326 THEN
            exp_f := 35;
        ELSIF x =- 8325 THEN
            exp_f := 35;
        ELSIF x =- 8324 THEN
            exp_f := 35;
        ELSIF x =- 8323 THEN
            exp_f := 35;
        ELSIF x =- 8322 THEN
            exp_f := 35;
        ELSIF x =- 8321 THEN
            exp_f := 35;
        ELSIF x =- 8320 THEN
            exp_f := 35;
        ELSIF x =- 8319 THEN
            exp_f := 35;
        ELSIF x =- 8318 THEN
            exp_f := 35;
        ELSIF x =- 8317 THEN
            exp_f := 35;
        ELSIF x =- 8316 THEN
            exp_f := 35;
        ELSIF x =- 8315 THEN
            exp_f := 35;
        ELSIF x =- 8314 THEN
            exp_f := 35;
        ELSIF x =- 8313 THEN
            exp_f := 35;
        ELSIF x =- 8312 THEN
            exp_f := 36;
        ELSIF x =- 8311 THEN
            exp_f := 36;
        ELSIF x =- 8310 THEN
            exp_f := 36;
        ELSIF x =- 8309 THEN
            exp_f := 36;
        ELSIF x =- 8308 THEN
            exp_f := 36;
        ELSIF x =- 8307 THEN
            exp_f := 36;
        ELSIF x =- 8306 THEN
            exp_f := 36;
        ELSIF x =- 8305 THEN
            exp_f := 36;
        ELSIF x =- 8304 THEN
            exp_f := 36;
        ELSIF x =- 8303 THEN
            exp_f := 36;
        ELSIF x =- 8302 THEN
            exp_f := 36;
        ELSIF x =- 8301 THEN
            exp_f := 36;
        ELSIF x =- 8300 THEN
            exp_f := 36;
        ELSIF x =- 8299 THEN
            exp_f := 36;
        ELSIF x =- 8298 THEN
            exp_f := 36;
        ELSIF x =- 8297 THEN
            exp_f := 36;
        ELSIF x =- 8296 THEN
            exp_f := 36;
        ELSIF x =- 8295 THEN
            exp_f := 36;
        ELSIF x =- 8294 THEN
            exp_f := 36;
        ELSIF x =- 8293 THEN
            exp_f := 36;
        ELSIF x =- 8292 THEN
            exp_f := 36;
        ELSIF x =- 8291 THEN
            exp_f := 36;
        ELSIF x =- 8290 THEN
            exp_f := 36;
        ELSIF x =- 8289 THEN
            exp_f := 36;
        ELSIF x =- 8288 THEN
            exp_f := 36;
        ELSIF x =- 8287 THEN
            exp_f := 36;
        ELSIF x =- 8286 THEN
            exp_f := 36;
        ELSIF x =- 8285 THEN
            exp_f := 36;
        ELSIF x =- 8284 THEN
            exp_f := 36;
        ELSIF x =- 8283 THEN
            exp_f := 36;
        ELSIF x =- 8282 THEN
            exp_f := 36;
        ELSIF x =- 8281 THEN
            exp_f := 36;
        ELSIF x =- 8280 THEN
            exp_f := 36;
        ELSIF x =- 8279 THEN
            exp_f := 36;
        ELSIF x =- 8278 THEN
            exp_f := 36;
        ELSIF x =- 8277 THEN
            exp_f := 36;
        ELSIF x =- 8276 THEN
            exp_f := 36;
        ELSIF x =- 8275 THEN
            exp_f := 36;
        ELSIF x =- 8274 THEN
            exp_f := 36;
        ELSIF x =- 8273 THEN
            exp_f := 36;
        ELSIF x =- 8272 THEN
            exp_f := 36;
        ELSIF x =- 8271 THEN
            exp_f := 36;
        ELSIF x =- 8270 THEN
            exp_f := 36;
        ELSIF x =- 8269 THEN
            exp_f := 36;
        ELSIF x =- 8268 THEN
            exp_f := 36;
        ELSIF x =- 8267 THEN
            exp_f := 36;
        ELSIF x =- 8266 THEN
            exp_f := 36;
        ELSIF x =- 8265 THEN
            exp_f := 36;
        ELSIF x =- 8264 THEN
            exp_f := 36;
        ELSIF x =- 8263 THEN
            exp_f := 36;
        ELSIF x =- 8262 THEN
            exp_f := 36;
        ELSIF x =- 8261 THEN
            exp_f := 36;
        ELSIF x =- 8260 THEN
            exp_f := 36;
        ELSIF x =- 8259 THEN
            exp_f := 36;
        ELSIF x =- 8258 THEN
            exp_f := 36;
        ELSIF x =- 8257 THEN
            exp_f := 36;
        ELSIF x =- 8256 THEN
            exp_f := 36;
        ELSIF x =- 8255 THEN
            exp_f := 36;
        ELSIF x =- 8254 THEN
            exp_f := 36;
        ELSIF x =- 8253 THEN
            exp_f := 36;
        ELSIF x =- 8252 THEN
            exp_f := 37;
        ELSIF x =- 8251 THEN
            exp_f := 37;
        ELSIF x =- 8250 THEN
            exp_f := 37;
        ELSIF x =- 8249 THEN
            exp_f := 37;
        ELSIF x =- 8248 THEN
            exp_f := 37;
        ELSIF x =- 8247 THEN
            exp_f := 37;
        ELSIF x =- 8246 THEN
            exp_f := 37;
        ELSIF x =- 8245 THEN
            exp_f := 37;
        ELSIF x =- 8244 THEN
            exp_f := 37;
        ELSIF x =- 8243 THEN
            exp_f := 37;
        ELSIF x =- 8242 THEN
            exp_f := 37;
        ELSIF x =- 8241 THEN
            exp_f := 37;
        ELSIF x =- 8240 THEN
            exp_f := 37;
        ELSIF x =- 8239 THEN
            exp_f := 37;
        ELSIF x =- 8238 THEN
            exp_f := 37;
        ELSIF x =- 8237 THEN
            exp_f := 37;
        ELSIF x =- 8236 THEN
            exp_f := 37;
        ELSIF x =- 8235 THEN
            exp_f := 37;
        ELSIF x =- 8234 THEN
            exp_f := 37;
        ELSIF x =- 8233 THEN
            exp_f := 37;
        ELSIF x =- 8232 THEN
            exp_f := 37;
        ELSIF x =- 8231 THEN
            exp_f := 37;
        ELSIF x =- 8230 THEN
            exp_f := 37;
        ELSIF x =- 8229 THEN
            exp_f := 37;
        ELSIF x =- 8228 THEN
            exp_f := 37;
        ELSIF x =- 8227 THEN
            exp_f := 37;
        ELSIF x =- 8226 THEN
            exp_f := 37;
        ELSIF x =- 8225 THEN
            exp_f := 37;
        ELSIF x =- 8224 THEN
            exp_f := 37;
        ELSIF x =- 8223 THEN
            exp_f := 37;
        ELSIF x =- 8222 THEN
            exp_f := 37;
        ELSIF x =- 8221 THEN
            exp_f := 37;
        ELSIF x =- 8220 THEN
            exp_f := 37;
        ELSIF x =- 8219 THEN
            exp_f := 37;
        ELSIF x =- 8218 THEN
            exp_f := 37;
        ELSIF x =- 8217 THEN
            exp_f := 37;
        ELSIF x =- 8216 THEN
            exp_f := 37;
        ELSIF x =- 8215 THEN
            exp_f := 37;
        ELSIF x =- 8214 THEN
            exp_f := 37;
        ELSIF x =- 8213 THEN
            exp_f := 37;
        ELSIF x =- 8212 THEN
            exp_f := 37;
        ELSIF x =- 8211 THEN
            exp_f := 37;
        ELSIF x =- 8210 THEN
            exp_f := 37;
        ELSIF x =- 8209 THEN
            exp_f := 37;
        ELSIF x =- 8208 THEN
            exp_f := 37;
        ELSIF x =- 8207 THEN
            exp_f := 37;
        ELSIF x =- 8206 THEN
            exp_f := 37;
        ELSIF x =- 8205 THEN
            exp_f := 37;
        ELSIF x =- 8204 THEN
            exp_f := 37;
        ELSIF x =- 8203 THEN
            exp_f := 37;
        ELSIF x =- 8202 THEN
            exp_f := 37;
        ELSIF x =- 8201 THEN
            exp_f := 37;
        ELSIF x =- 8200 THEN
            exp_f := 37;
        ELSIF x =- 8199 THEN
            exp_f := 37;
        ELSIF x =- 8198 THEN
            exp_f := 37;
        ELSIF x =- 8197 THEN
            exp_f := 37;
        ELSIF x =- 8196 THEN
            exp_f := 37;
        ELSIF x =- 8195 THEN
            exp_f := 37;
        ELSIF x =- 8194 THEN
            exp_f := 37;
        ELSIF x =- 8193 THEN
            exp_f := 37;
        ELSIF x =- 8192 THEN
            exp_f := 37;
        ELSIF x =- 8191 THEN
            exp_f := 38;
        ELSIF x =- 8190 THEN
            exp_f := 38;
        ELSIF x =- 8189 THEN
            exp_f := 38;
        ELSIF x =- 8188 THEN
            exp_f := 38;
        ELSIF x =- 8187 THEN
            exp_f := 38;
        ELSIF x =- 8186 THEN
            exp_f := 38;
        ELSIF x =- 8185 THEN
            exp_f := 38;
        ELSIF x =- 8184 THEN
            exp_f := 38;
        ELSIF x =- 8183 THEN
            exp_f := 38;
        ELSIF x =- 8182 THEN
            exp_f := 38;
        ELSIF x =- 8181 THEN
            exp_f := 38;
        ELSIF x =- 8180 THEN
            exp_f := 38;
        ELSIF x =- 8179 THEN
            exp_f := 38;
        ELSIF x =- 8178 THEN
            exp_f := 38;
        ELSIF x =- 8177 THEN
            exp_f := 38;
        ELSIF x =- 8176 THEN
            exp_f := 38;
        ELSIF x =- 8175 THEN
            exp_f := 38;
        ELSIF x =- 8174 THEN
            exp_f := 38;
        ELSIF x =- 8173 THEN
            exp_f := 38;
        ELSIF x =- 8172 THEN
            exp_f := 38;
        ELSIF x =- 8171 THEN
            exp_f := 38;
        ELSIF x =- 8170 THEN
            exp_f := 38;
        ELSIF x =- 8169 THEN
            exp_f := 38;
        ELSIF x =- 8168 THEN
            exp_f := 38;
        ELSIF x =- 8167 THEN
            exp_f := 38;
        ELSIF x =- 8166 THEN
            exp_f := 38;
        ELSIF x =- 8165 THEN
            exp_f := 38;
        ELSIF x =- 8164 THEN
            exp_f := 38;
        ELSIF x =- 8163 THEN
            exp_f := 38;
        ELSIF x =- 8162 THEN
            exp_f := 38;
        ELSIF x =- 8161 THEN
            exp_f := 38;
        ELSIF x =- 8160 THEN
            exp_f := 38;
        ELSIF x =- 8159 THEN
            exp_f := 38;
        ELSIF x =- 8158 THEN
            exp_f := 38;
        ELSIF x =- 8157 THEN
            exp_f := 38;
        ELSIF x =- 8156 THEN
            exp_f := 38;
        ELSIF x =- 8155 THEN
            exp_f := 38;
        ELSIF x =- 8154 THEN
            exp_f := 38;
        ELSIF x =- 8153 THEN
            exp_f := 38;
        ELSIF x =- 8152 THEN
            exp_f := 38;
        ELSIF x =- 8151 THEN
            exp_f := 38;
        ELSIF x =- 8150 THEN
            exp_f := 38;
        ELSIF x =- 8149 THEN
            exp_f := 38;
        ELSIF x =- 8148 THEN
            exp_f := 38;
        ELSIF x =- 8147 THEN
            exp_f := 38;
        ELSIF x =- 8146 THEN
            exp_f := 38;
        ELSIF x =- 8145 THEN
            exp_f := 38;
        ELSIF x =- 8144 THEN
            exp_f := 38;
        ELSIF x =- 8143 THEN
            exp_f := 38;
        ELSIF x =- 8142 THEN
            exp_f := 38;
        ELSIF x =- 8141 THEN
            exp_f := 38;
        ELSIF x =- 8140 THEN
            exp_f := 38;
        ELSIF x =- 8139 THEN
            exp_f := 39;
        ELSIF x =- 8138 THEN
            exp_f := 39;
        ELSIF x =- 8137 THEN
            exp_f := 39;
        ELSIF x =- 8136 THEN
            exp_f := 39;
        ELSIF x =- 8135 THEN
            exp_f := 39;
        ELSIF x =- 8134 THEN
            exp_f := 39;
        ELSIF x =- 8133 THEN
            exp_f := 39;
        ELSIF x =- 8132 THEN
            exp_f := 39;
        ELSIF x =- 8131 THEN
            exp_f := 39;
        ELSIF x =- 8130 THEN
            exp_f := 39;
        ELSIF x =- 8129 THEN
            exp_f := 39;
        ELSIF x =- 8128 THEN
            exp_f := 39;
        ELSIF x =- 8127 THEN
            exp_f := 39;
        ELSIF x =- 8126 THEN
            exp_f := 39;
        ELSIF x =- 8125 THEN
            exp_f := 39;
        ELSIF x =- 8124 THEN
            exp_f := 39;
        ELSIF x =- 8123 THEN
            exp_f := 39;
        ELSIF x =- 8122 THEN
            exp_f := 39;
        ELSIF x =- 8121 THEN
            exp_f := 39;
        ELSIF x =- 8120 THEN
            exp_f := 39;
        ELSIF x =- 8119 THEN
            exp_f := 39;
        ELSIF x =- 8118 THEN
            exp_f := 39;
        ELSIF x =- 8117 THEN
            exp_f := 39;
        ELSIF x =- 8116 THEN
            exp_f := 39;
        ELSIF x =- 8115 THEN
            exp_f := 39;
        ELSIF x =- 8114 THEN
            exp_f := 39;
        ELSIF x =- 8113 THEN
            exp_f := 39;
        ELSIF x =- 8112 THEN
            exp_f := 39;
        ELSIF x =- 8111 THEN
            exp_f := 39;
        ELSIF x =- 8110 THEN
            exp_f := 39;
        ELSIF x =- 8109 THEN
            exp_f := 39;
        ELSIF x =- 8108 THEN
            exp_f := 39;
        ELSIF x =- 8107 THEN
            exp_f := 39;
        ELSIF x =- 8106 THEN
            exp_f := 39;
        ELSIF x =- 8105 THEN
            exp_f := 39;
        ELSIF x =- 8104 THEN
            exp_f := 39;
        ELSIF x =- 8103 THEN
            exp_f := 39;
        ELSIF x =- 8102 THEN
            exp_f := 39;
        ELSIF x =- 8101 THEN
            exp_f := 39;
        ELSIF x =- 8100 THEN
            exp_f := 39;
        ELSIF x =- 8099 THEN
            exp_f := 39;
        ELSIF x =- 8098 THEN
            exp_f := 39;
        ELSIF x =- 8097 THEN
            exp_f := 39;
        ELSIF x =- 8096 THEN
            exp_f := 39;
        ELSIF x =- 8095 THEN
            exp_f := 39;
        ELSIF x =- 8094 THEN
            exp_f := 39;
        ELSIF x =- 8093 THEN
            exp_f := 39;
        ELSIF x =- 8092 THEN
            exp_f := 39;
        ELSIF x =- 8091 THEN
            exp_f := 39;
        ELSIF x =- 8090 THEN
            exp_f := 39;
        ELSIF x =- 8089 THEN
            exp_f := 39;
        ELSIF x =- 8088 THEN
            exp_f := 39;
        ELSIF x =- 8087 THEN
            exp_f := 39;
        ELSIF x =- 8086 THEN
            exp_f := 40;
        ELSIF x =- 8085 THEN
            exp_f := 40;
        ELSIF x =- 8084 THEN
            exp_f := 40;
        ELSIF x =- 8083 THEN
            exp_f := 40;
        ELSIF x =- 8082 THEN
            exp_f := 40;
        ELSIF x =- 8081 THEN
            exp_f := 40;
        ELSIF x =- 8080 THEN
            exp_f := 40;
        ELSIF x =- 8079 THEN
            exp_f := 40;
        ELSIF x =- 8078 THEN
            exp_f := 40;
        ELSIF x =- 8077 THEN
            exp_f := 40;
        ELSIF x =- 8076 THEN
            exp_f := 40;
        ELSIF x =- 8075 THEN
            exp_f := 40;
        ELSIF x =- 8074 THEN
            exp_f := 40;
        ELSIF x =- 8073 THEN
            exp_f := 40;
        ELSIF x =- 8072 THEN
            exp_f := 40;
        ELSIF x =- 8071 THEN
            exp_f := 40;
        ELSIF x =- 8070 THEN
            exp_f := 40;
        ELSIF x =- 8069 THEN
            exp_f := 40;
        ELSIF x =- 8068 THEN
            exp_f := 40;
        ELSIF x =- 8067 THEN
            exp_f := 40;
        ELSIF x =- 8066 THEN
            exp_f := 40;
        ELSIF x =- 8065 THEN
            exp_f := 40;
        ELSIF x =- 8064 THEN
            exp_f := 40;
        ELSIF x =- 8063 THEN
            exp_f := 40;
        ELSIF x =- 8062 THEN
            exp_f := 40;
        ELSIF x =- 8061 THEN
            exp_f := 40;
        ELSIF x =- 8060 THEN
            exp_f := 40;
        ELSIF x =- 8059 THEN
            exp_f := 40;
        ELSIF x =- 8058 THEN
            exp_f := 40;
        ELSIF x =- 8057 THEN
            exp_f := 40;
        ELSIF x =- 8056 THEN
            exp_f := 40;
        ELSIF x =- 8055 THEN
            exp_f := 40;
        ELSIF x =- 8054 THEN
            exp_f := 40;
        ELSIF x =- 8053 THEN
            exp_f := 40;
        ELSIF x =- 8052 THEN
            exp_f := 40;
        ELSIF x =- 8051 THEN
            exp_f := 40;
        ELSIF x =- 8050 THEN
            exp_f := 40;
        ELSIF x =- 8049 THEN
            exp_f := 40;
        ELSIF x =- 8048 THEN
            exp_f := 40;
        ELSIF x =- 8047 THEN
            exp_f := 40;
        ELSIF x =- 8046 THEN
            exp_f := 40;
        ELSIF x =- 8045 THEN
            exp_f := 40;
        ELSIF x =- 8044 THEN
            exp_f := 40;
        ELSIF x =- 8043 THEN
            exp_f := 40;
        ELSIF x =- 8042 THEN
            exp_f := 40;
        ELSIF x =- 8041 THEN
            exp_f := 40;
        ELSIF x =- 8040 THEN
            exp_f := 40;
        ELSIF x =- 8039 THEN
            exp_f := 40;
        ELSIF x =- 8038 THEN
            exp_f := 40;
        ELSIF x =- 8037 THEN
            exp_f := 40;
        ELSIF x =- 8036 THEN
            exp_f := 40;
        ELSIF x =- 8035 THEN
            exp_f := 40;
        ELSIF x =- 8034 THEN
            exp_f := 41;
        ELSIF x =- 8033 THEN
            exp_f := 41;
        ELSIF x =- 8032 THEN
            exp_f := 41;
        ELSIF x =- 8031 THEN
            exp_f := 41;
        ELSIF x =- 8030 THEN
            exp_f := 41;
        ELSIF x =- 8029 THEN
            exp_f := 41;
        ELSIF x =- 8028 THEN
            exp_f := 41;
        ELSIF x =- 8027 THEN
            exp_f := 41;
        ELSIF x =- 8026 THEN
            exp_f := 41;
        ELSIF x =- 8025 THEN
            exp_f := 41;
        ELSIF x =- 8024 THEN
            exp_f := 41;
        ELSIF x =- 8023 THEN
            exp_f := 41;
        ELSIF x =- 8022 THEN
            exp_f := 41;
        ELSIF x =- 8021 THEN
            exp_f := 41;
        ELSIF x =- 8020 THEN
            exp_f := 41;
        ELSIF x =- 8019 THEN
            exp_f := 41;
        ELSIF x =- 8018 THEN
            exp_f := 41;
        ELSIF x =- 8017 THEN
            exp_f := 41;
        ELSIF x =- 8016 THEN
            exp_f := 41;
        ELSIF x =- 8015 THEN
            exp_f := 41;
        ELSIF x =- 8014 THEN
            exp_f := 41;
        ELSIF x =- 8013 THEN
            exp_f := 41;
        ELSIF x =- 8012 THEN
            exp_f := 41;
        ELSIF x =- 8011 THEN
            exp_f := 41;
        ELSIF x =- 8010 THEN
            exp_f := 41;
        ELSIF x =- 8009 THEN
            exp_f := 41;
        ELSIF x =- 8008 THEN
            exp_f := 41;
        ELSIF x =- 8007 THEN
            exp_f := 41;
        ELSIF x =- 8006 THEN
            exp_f := 41;
        ELSIF x =- 8005 THEN
            exp_f := 41;
        ELSIF x =- 8004 THEN
            exp_f := 41;
        ELSIF x =- 8003 THEN
            exp_f := 41;
        ELSIF x =- 8002 THEN
            exp_f := 41;
        ELSIF x =- 8001 THEN
            exp_f := 41;
        ELSIF x =- 8000 THEN
            exp_f := 41;
        ELSIF x =- 7999 THEN
            exp_f := 41;
        ELSIF x =- 7998 THEN
            exp_f := 41;
        ELSIF x =- 7997 THEN
            exp_f := 41;
        ELSIF x =- 7996 THEN
            exp_f := 41;
        ELSIF x =- 7995 THEN
            exp_f := 41;
        ELSIF x =- 7994 THEN
            exp_f := 41;
        ELSIF x =- 7993 THEN
            exp_f := 41;
        ELSIF x =- 7992 THEN
            exp_f := 41;
        ELSIF x =- 7991 THEN
            exp_f := 41;
        ELSIF x =- 7990 THEN
            exp_f := 41;
        ELSIF x =- 7989 THEN
            exp_f := 41;
        ELSIF x =- 7988 THEN
            exp_f := 41;
        ELSIF x =- 7987 THEN
            exp_f := 41;
        ELSIF x =- 7986 THEN
            exp_f := 41;
        ELSIF x =- 7985 THEN
            exp_f := 41;
        ELSIF x =- 7984 THEN
            exp_f := 41;
        ELSIF x =- 7983 THEN
            exp_f := 41;
        ELSIF x =- 7982 THEN
            exp_f := 41;
        ELSIF x =- 7981 THEN
            exp_f := 42;
        ELSIF x =- 7980 THEN
            exp_f := 42;
        ELSIF x =- 7979 THEN
            exp_f := 42;
        ELSIF x =- 7978 THEN
            exp_f := 42;
        ELSIF x =- 7977 THEN
            exp_f := 42;
        ELSIF x =- 7976 THEN
            exp_f := 42;
        ELSIF x =- 7975 THEN
            exp_f := 42;
        ELSIF x =- 7974 THEN
            exp_f := 42;
        ELSIF x =- 7973 THEN
            exp_f := 42;
        ELSIF x =- 7972 THEN
            exp_f := 42;
        ELSIF x =- 7971 THEN
            exp_f := 42;
        ELSIF x =- 7970 THEN
            exp_f := 42;
        ELSIF x =- 7969 THEN
            exp_f := 42;
        ELSIF x =- 7968 THEN
            exp_f := 42;
        ELSIF x =- 7967 THEN
            exp_f := 42;
        ELSIF x =- 7966 THEN
            exp_f := 42;
        ELSIF x =- 7965 THEN
            exp_f := 42;
        ELSIF x =- 7964 THEN
            exp_f := 42;
        ELSIF x =- 7963 THEN
            exp_f := 42;
        ELSIF x =- 7962 THEN
            exp_f := 42;
        ELSIF x =- 7961 THEN
            exp_f := 42;
        ELSIF x =- 7960 THEN
            exp_f := 42;
        ELSIF x =- 7959 THEN
            exp_f := 42;
        ELSIF x =- 7958 THEN
            exp_f := 42;
        ELSIF x =- 7957 THEN
            exp_f := 42;
        ELSIF x =- 7956 THEN
            exp_f := 42;
        ELSIF x =- 7955 THEN
            exp_f := 42;
        ELSIF x =- 7954 THEN
            exp_f := 42;
        ELSIF x =- 7953 THEN
            exp_f := 42;
        ELSIF x =- 7952 THEN
            exp_f := 42;
        ELSIF x =- 7951 THEN
            exp_f := 42;
        ELSIF x =- 7950 THEN
            exp_f := 42;
        ELSIF x =- 7949 THEN
            exp_f := 42;
        ELSIF x =- 7948 THEN
            exp_f := 42;
        ELSIF x =- 7947 THEN
            exp_f := 42;
        ELSIF x =- 7946 THEN
            exp_f := 42;
        ELSIF x =- 7945 THEN
            exp_f := 42;
        ELSIF x =- 7944 THEN
            exp_f := 42;
        ELSIF x =- 7943 THEN
            exp_f := 42;
        ELSIF x =- 7942 THEN
            exp_f := 42;
        ELSIF x =- 7941 THEN
            exp_f := 42;
        ELSIF x =- 7940 THEN
            exp_f := 42;
        ELSIF x =- 7939 THEN
            exp_f := 42;
        ELSIF x =- 7938 THEN
            exp_f := 42;
        ELSIF x =- 7937 THEN
            exp_f := 42;
        ELSIF x =- 7936 THEN
            exp_f := 42;
        ELSIF x =- 7935 THEN
            exp_f := 42;
        ELSIF x =- 7934 THEN
            exp_f := 42;
        ELSIF x =- 7933 THEN
            exp_f := 42;
        ELSIF x =- 7932 THEN
            exp_f := 42;
        ELSIF x =- 7931 THEN
            exp_f := 42;
        ELSIF x =- 7930 THEN
            exp_f := 42;
        ELSIF x =- 7929 THEN
            exp_f := 43;
        ELSIF x =- 7928 THEN
            exp_f := 43;
        ELSIF x =- 7927 THEN
            exp_f := 43;
        ELSIF x =- 7926 THEN
            exp_f := 43;
        ELSIF x =- 7925 THEN
            exp_f := 43;
        ELSIF x =- 7924 THEN
            exp_f := 43;
        ELSIF x =- 7923 THEN
            exp_f := 43;
        ELSIF x =- 7922 THEN
            exp_f := 43;
        ELSIF x =- 7921 THEN
            exp_f := 43;
        ELSIF x =- 7920 THEN
            exp_f := 43;
        ELSIF x =- 7919 THEN
            exp_f := 43;
        ELSIF x =- 7918 THEN
            exp_f := 43;
        ELSIF x =- 7917 THEN
            exp_f := 43;
        ELSIF x =- 7916 THEN
            exp_f := 43;
        ELSIF x =- 7915 THEN
            exp_f := 43;
        ELSIF x =- 7914 THEN
            exp_f := 43;
        ELSIF x =- 7913 THEN
            exp_f := 43;
        ELSIF x =- 7912 THEN
            exp_f := 43;
        ELSIF x =- 7911 THEN
            exp_f := 43;
        ELSIF x =- 7910 THEN
            exp_f := 43;
        ELSIF x =- 7909 THEN
            exp_f := 43;
        ELSIF x =- 7908 THEN
            exp_f := 43;
        ELSIF x =- 7907 THEN
            exp_f := 43;
        ELSIF x =- 7906 THEN
            exp_f := 43;
        ELSIF x =- 7905 THEN
            exp_f := 43;
        ELSIF x =- 7904 THEN
            exp_f := 43;
        ELSIF x =- 7903 THEN
            exp_f := 43;
        ELSIF x =- 7902 THEN
            exp_f := 43;
        ELSIF x =- 7901 THEN
            exp_f := 43;
        ELSIF x =- 7900 THEN
            exp_f := 43;
        ELSIF x =- 7899 THEN
            exp_f := 43;
        ELSIF x =- 7898 THEN
            exp_f := 43;
        ELSIF x =- 7897 THEN
            exp_f := 43;
        ELSIF x =- 7896 THEN
            exp_f := 43;
        ELSIF x =- 7895 THEN
            exp_f := 43;
        ELSIF x =- 7894 THEN
            exp_f := 43;
        ELSIF x =- 7893 THEN
            exp_f := 43;
        ELSIF x =- 7892 THEN
            exp_f := 43;
        ELSIF x =- 7891 THEN
            exp_f := 43;
        ELSIF x =- 7890 THEN
            exp_f := 43;
        ELSIF x =- 7889 THEN
            exp_f := 43;
        ELSIF x =- 7888 THEN
            exp_f := 43;
        ELSIF x =- 7887 THEN
            exp_f := 43;
        ELSIF x =- 7886 THEN
            exp_f := 43;
        ELSIF x =- 7885 THEN
            exp_f := 43;
        ELSIF x =- 7884 THEN
            exp_f := 43;
        ELSIF x =- 7883 THEN
            exp_f := 43;
        ELSIF x =- 7882 THEN
            exp_f := 43;
        ELSIF x =- 7881 THEN
            exp_f := 43;
        ELSIF x =- 7880 THEN
            exp_f := 43;
        ELSIF x =- 7879 THEN
            exp_f := 43;
        ELSIF x =- 7878 THEN
            exp_f := 43;
        ELSIF x =- 7877 THEN
            exp_f := 43;
        ELSIF x =- 7876 THEN
            exp_f := 44;
        ELSIF x =- 7875 THEN
            exp_f := 44;
        ELSIF x =- 7874 THEN
            exp_f := 44;
        ELSIF x =- 7873 THEN
            exp_f := 44;
        ELSIF x =- 7872 THEN
            exp_f := 44;
        ELSIF x =- 7871 THEN
            exp_f := 44;
        ELSIF x =- 7870 THEN
            exp_f := 44;
        ELSIF x =- 7869 THEN
            exp_f := 44;
        ELSIF x =- 7868 THEN
            exp_f := 44;
        ELSIF x =- 7867 THEN
            exp_f := 44;
        ELSIF x =- 7866 THEN
            exp_f := 44;
        ELSIF x =- 7865 THEN
            exp_f := 44;
        ELSIF x =- 7864 THEN
            exp_f := 44;
        ELSIF x =- 7863 THEN
            exp_f := 44;
        ELSIF x =- 7862 THEN
            exp_f := 44;
        ELSIF x =- 7861 THEN
            exp_f := 44;
        ELSIF x =- 7860 THEN
            exp_f := 44;
        ELSIF x =- 7859 THEN
            exp_f := 44;
        ELSIF x =- 7858 THEN
            exp_f := 44;
        ELSIF x =- 7857 THEN
            exp_f := 44;
        ELSIF x =- 7856 THEN
            exp_f := 44;
        ELSIF x =- 7855 THEN
            exp_f := 44;
        ELSIF x =- 7854 THEN
            exp_f := 44;
        ELSIF x =- 7853 THEN
            exp_f := 44;
        ELSIF x =- 7852 THEN
            exp_f := 44;
        ELSIF x =- 7851 THEN
            exp_f := 44;
        ELSIF x =- 7850 THEN
            exp_f := 44;
        ELSIF x =- 7849 THEN
            exp_f := 44;
        ELSIF x =- 7848 THEN
            exp_f := 44;
        ELSIF x =- 7847 THEN
            exp_f := 44;
        ELSIF x =- 7846 THEN
            exp_f := 44;
        ELSIF x =- 7845 THEN
            exp_f := 44;
        ELSIF x =- 7844 THEN
            exp_f := 44;
        ELSIF x =- 7843 THEN
            exp_f := 44;
        ELSIF x =- 7842 THEN
            exp_f := 44;
        ELSIF x =- 7841 THEN
            exp_f := 44;
        ELSIF x =- 7840 THEN
            exp_f := 44;
        ELSIF x =- 7839 THEN
            exp_f := 44;
        ELSIF x =- 7838 THEN
            exp_f := 44;
        ELSIF x =- 7837 THEN
            exp_f := 44;
        ELSIF x =- 7836 THEN
            exp_f := 44;
        ELSIF x =- 7835 THEN
            exp_f := 44;
        ELSIF x =- 7834 THEN
            exp_f := 44;
        ELSIF x =- 7833 THEN
            exp_f := 44;
        ELSIF x =- 7832 THEN
            exp_f := 44;
        ELSIF x =- 7831 THEN
            exp_f := 44;
        ELSIF x =- 7830 THEN
            exp_f := 44;
        ELSIF x =- 7829 THEN
            exp_f := 44;
        ELSIF x =- 7828 THEN
            exp_f := 44;
        ELSIF x =- 7827 THEN
            exp_f := 44;
        ELSIF x =- 7826 THEN
            exp_f := 44;
        ELSIF x =- 7825 THEN
            exp_f := 44;
        ELSIF x =- 7824 THEN
            exp_f := 46;
        ELSIF x =- 7823 THEN
            exp_f := 46;
        ELSIF x =- 7822 THEN
            exp_f := 46;
        ELSIF x =- 7821 THEN
            exp_f := 46;
        ELSIF x =- 7820 THEN
            exp_f := 46;
        ELSIF x =- 7819 THEN
            exp_f := 46;
        ELSIF x =- 7818 THEN
            exp_f := 46;
        ELSIF x =- 7817 THEN
            exp_f := 46;
        ELSIF x =- 7816 THEN
            exp_f := 46;
        ELSIF x =- 7815 THEN
            exp_f := 46;
        ELSIF x =- 7814 THEN
            exp_f := 46;
        ELSIF x =- 7813 THEN
            exp_f := 46;
        ELSIF x =- 7812 THEN
            exp_f := 46;
        ELSIF x =- 7811 THEN
            exp_f := 46;
        ELSIF x =- 7810 THEN
            exp_f := 46;
        ELSIF x =- 7809 THEN
            exp_f := 46;
        ELSIF x =- 7808 THEN
            exp_f := 46;
        ELSIF x =- 7807 THEN
            exp_f := 46;
        ELSIF x =- 7806 THEN
            exp_f := 46;
        ELSIF x =- 7805 THEN
            exp_f := 46;
        ELSIF x =- 7804 THEN
            exp_f := 46;
        ELSIF x =- 7803 THEN
            exp_f := 46;
        ELSIF x =- 7802 THEN
            exp_f := 46;
        ELSIF x =- 7801 THEN
            exp_f := 46;
        ELSIF x =- 7800 THEN
            exp_f := 46;
        ELSIF x =- 7799 THEN
            exp_f := 46;
        ELSIF x =- 7798 THEN
            exp_f := 46;
        ELSIF x =- 7797 THEN
            exp_f := 46;
        ELSIF x =- 7796 THEN
            exp_f := 46;
        ELSIF x =- 7795 THEN
            exp_f := 46;
        ELSIF x =- 7794 THEN
            exp_f := 46;
        ELSIF x =- 7793 THEN
            exp_f := 46;
        ELSIF x =- 7792 THEN
            exp_f := 46;
        ELSIF x =- 7791 THEN
            exp_f := 46;
        ELSIF x =- 7790 THEN
            exp_f := 46;
        ELSIF x =- 7789 THEN
            exp_f := 46;
        ELSIF x =- 7788 THEN
            exp_f := 46;
        ELSIF x =- 7787 THEN
            exp_f := 46;
        ELSIF x =- 7786 THEN
            exp_f := 46;
        ELSIF x =- 7785 THEN
            exp_f := 46;
        ELSIF x =- 7784 THEN
            exp_f := 46;
        ELSIF x =- 7783 THEN
            exp_f := 46;
        ELSIF x =- 7782 THEN
            exp_f := 46;
        ELSIF x =- 7781 THEN
            exp_f := 46;
        ELSIF x =- 7780 THEN
            exp_f := 46;
        ELSIF x =- 7779 THEN
            exp_f := 46;
        ELSIF x =- 7778 THEN
            exp_f := 46;
        ELSIF x =- 7777 THEN
            exp_f := 46;
        ELSIF x =- 7776 THEN
            exp_f := 46;
        ELSIF x =- 7775 THEN
            exp_f := 46;
        ELSIF x =- 7774 THEN
            exp_f := 46;
        ELSIF x =- 7773 THEN
            exp_f := 46;
        ELSIF x =- 7772 THEN
            exp_f := 46;
        ELSIF x =- 7771 THEN
            exp_f := 47;
        ELSIF x =- 7770 THEN
            exp_f := 47;
        ELSIF x =- 7769 THEN
            exp_f := 47;
        ELSIF x =- 7768 THEN
            exp_f := 47;
        ELSIF x =- 7767 THEN
            exp_f := 47;
        ELSIF x =- 7766 THEN
            exp_f := 47;
        ELSIF x =- 7765 THEN
            exp_f := 47;
        ELSIF x =- 7764 THEN
            exp_f := 47;
        ELSIF x =- 7763 THEN
            exp_f := 47;
        ELSIF x =- 7762 THEN
            exp_f := 47;
        ELSIF x =- 7761 THEN
            exp_f := 47;
        ELSIF x =- 7760 THEN
            exp_f := 47;
        ELSIF x =- 7759 THEN
            exp_f := 47;
        ELSIF x =- 7758 THEN
            exp_f := 47;
        ELSIF x =- 7757 THEN
            exp_f := 47;
        ELSIF x =- 7756 THEN
            exp_f := 47;
        ELSIF x =- 7755 THEN
            exp_f := 47;
        ELSIF x =- 7754 THEN
            exp_f := 47;
        ELSIF x =- 7753 THEN
            exp_f := 47;
        ELSIF x =- 7752 THEN
            exp_f := 47;
        ELSIF x =- 7751 THEN
            exp_f := 47;
        ELSIF x =- 7750 THEN
            exp_f := 47;
        ELSIF x =- 7749 THEN
            exp_f := 47;
        ELSIF x =- 7748 THEN
            exp_f := 47;
        ELSIF x =- 7747 THEN
            exp_f := 47;
        ELSIF x =- 7746 THEN
            exp_f := 47;
        ELSIF x =- 7745 THEN
            exp_f := 47;
        ELSIF x =- 7744 THEN
            exp_f := 47;
        ELSIF x =- 7743 THEN
            exp_f := 47;
        ELSIF x =- 7742 THEN
            exp_f := 47;
        ELSIF x =- 7741 THEN
            exp_f := 47;
        ELSIF x =- 7740 THEN
            exp_f := 47;
        ELSIF x =- 7739 THEN
            exp_f := 47;
        ELSIF x =- 7738 THEN
            exp_f := 47;
        ELSIF x =- 7737 THEN
            exp_f := 47;
        ELSIF x =- 7736 THEN
            exp_f := 47;
        ELSIF x =- 7735 THEN
            exp_f := 47;
        ELSIF x =- 7734 THEN
            exp_f := 47;
        ELSIF x =- 7733 THEN
            exp_f := 47;
        ELSIF x =- 7732 THEN
            exp_f := 47;
        ELSIF x =- 7731 THEN
            exp_f := 47;
        ELSIF x =- 7730 THEN
            exp_f := 47;
        ELSIF x =- 7729 THEN
            exp_f := 47;
        ELSIF x =- 7728 THEN
            exp_f := 47;
        ELSIF x =- 7727 THEN
            exp_f := 47;
        ELSIF x =- 7726 THEN
            exp_f := 47;
        ELSIF x =- 7725 THEN
            exp_f := 47;
        ELSIF x =- 7724 THEN
            exp_f := 47;
        ELSIF x =- 7723 THEN
            exp_f := 47;
        ELSIF x =- 7722 THEN
            exp_f := 47;
        ELSIF x =- 7721 THEN
            exp_f := 47;
        ELSIF x =- 7720 THEN
            exp_f := 47;
        ELSIF x =- 7719 THEN
            exp_f := 48;
        ELSIF x =- 7718 THEN
            exp_f := 48;
        ELSIF x =- 7717 THEN
            exp_f := 48;
        ELSIF x =- 7716 THEN
            exp_f := 48;
        ELSIF x =- 7715 THEN
            exp_f := 48;
        ELSIF x =- 7714 THEN
            exp_f := 48;
        ELSIF x =- 7713 THEN
            exp_f := 48;
        ELSIF x =- 7712 THEN
            exp_f := 48;
        ELSIF x =- 7711 THEN
            exp_f := 48;
        ELSIF x =- 7710 THEN
            exp_f := 48;
        ELSIF x =- 7709 THEN
            exp_f := 48;
        ELSIF x =- 7708 THEN
            exp_f := 48;
        ELSIF x =- 7707 THEN
            exp_f := 48;
        ELSIF x =- 7706 THEN
            exp_f := 48;
        ELSIF x =- 7705 THEN
            exp_f := 48;
        ELSIF x =- 7704 THEN
            exp_f := 48;
        ELSIF x =- 7703 THEN
            exp_f := 48;
        ELSIF x =- 7702 THEN
            exp_f := 48;
        ELSIF x =- 7701 THEN
            exp_f := 48;
        ELSIF x =- 7700 THEN
            exp_f := 48;
        ELSIF x =- 7699 THEN
            exp_f := 48;
        ELSIF x =- 7698 THEN
            exp_f := 48;
        ELSIF x =- 7697 THEN
            exp_f := 48;
        ELSIF x =- 7696 THEN
            exp_f := 48;
        ELSIF x =- 7695 THEN
            exp_f := 48;
        ELSIF x =- 7694 THEN
            exp_f := 48;
        ELSIF x =- 7693 THEN
            exp_f := 48;
        ELSIF x =- 7692 THEN
            exp_f := 48;
        ELSIF x =- 7691 THEN
            exp_f := 48;
        ELSIF x =- 7690 THEN
            exp_f := 48;
        ELSIF x =- 7689 THEN
            exp_f := 48;
        ELSIF x =- 7688 THEN
            exp_f := 48;
        ELSIF x =- 7687 THEN
            exp_f := 48;
        ELSIF x =- 7686 THEN
            exp_f := 48;
        ELSIF x =- 7685 THEN
            exp_f := 48;
        ELSIF x =- 7684 THEN
            exp_f := 48;
        ELSIF x =- 7683 THEN
            exp_f := 48;
        ELSIF x =- 7682 THEN
            exp_f := 48;
        ELSIF x =- 7681 THEN
            exp_f := 48;
        ELSIF x =- 7680 THEN
            exp_f := 48;
        ELSIF x =- 7679 THEN
            exp_f := 48;
        ELSIF x =- 7678 THEN
            exp_f := 48;
        ELSIF x =- 7677 THEN
            exp_f := 48;
        ELSIF x =- 7676 THEN
            exp_f := 48;
        ELSIF x =- 7675 THEN
            exp_f := 48;
        ELSIF x =- 7674 THEN
            exp_f := 48;
        ELSIF x =- 7673 THEN
            exp_f := 48;
        ELSIF x =- 7672 THEN
            exp_f := 48;
        ELSIF x =- 7671 THEN
            exp_f := 48;
        ELSIF x =- 7670 THEN
            exp_f := 48;
        ELSIF x =- 7669 THEN
            exp_f := 48;
        ELSIF x =- 7668 THEN
            exp_f := 48;
        ELSIF x =- 7667 THEN
            exp_f := 48;
        ELSIF x =- 7666 THEN
            exp_f := 48;
        ELSIF x =- 7665 THEN
            exp_f := 48;
        ELSIF x =- 7664 THEN
            exp_f := 48;
        ELSIF x =- 7663 THEN
            exp_f := 48;
        ELSIF x =- 7662 THEN
            exp_f := 48;
        ELSIF x =- 7661 THEN
            exp_f := 49;
        ELSIF x =- 7660 THEN
            exp_f := 49;
        ELSIF x =- 7659 THEN
            exp_f := 49;
        ELSIF x =- 7658 THEN
            exp_f := 49;
        ELSIF x =- 7657 THEN
            exp_f := 49;
        ELSIF x =- 7656 THEN
            exp_f := 49;
        ELSIF x =- 7655 THEN
            exp_f := 49;
        ELSIF x =- 7654 THEN
            exp_f := 49;
        ELSIF x =- 7653 THEN
            exp_f := 49;
        ELSIF x =- 7652 THEN
            exp_f := 49;
        ELSIF x =- 7651 THEN
            exp_f := 49;
        ELSIF x =- 7650 THEN
            exp_f := 49;
        ELSIF x =- 7649 THEN
            exp_f := 49;
        ELSIF x =- 7648 THEN
            exp_f := 49;
        ELSIF x =- 7647 THEN
            exp_f := 49;
        ELSIF x =- 7646 THEN
            exp_f := 49;
        ELSIF x =- 7645 THEN
            exp_f := 49;
        ELSIF x =- 7644 THEN
            exp_f := 49;
        ELSIF x =- 7643 THEN
            exp_f := 49;
        ELSIF x =- 7642 THEN
            exp_f := 49;
        ELSIF x =- 7641 THEN
            exp_f := 49;
        ELSIF x =- 7640 THEN
            exp_f := 49;
        ELSIF x =- 7639 THEN
            exp_f := 49;
        ELSIF x =- 7638 THEN
            exp_f := 49;
        ELSIF x =- 7637 THEN
            exp_f := 49;
        ELSIF x =- 7636 THEN
            exp_f := 49;
        ELSIF x =- 7635 THEN
            exp_f := 49;
        ELSIF x =- 7634 THEN
            exp_f := 49;
        ELSIF x =- 7633 THEN
            exp_f := 49;
        ELSIF x =- 7632 THEN
            exp_f := 49;
        ELSIF x =- 7631 THEN
            exp_f := 49;
        ELSIF x =- 7630 THEN
            exp_f := 49;
        ELSIF x =- 7629 THEN
            exp_f := 49;
        ELSIF x =- 7628 THEN
            exp_f := 49;
        ELSIF x =- 7627 THEN
            exp_f := 49;
        ELSIF x =- 7626 THEN
            exp_f := 49;
        ELSIF x =- 7625 THEN
            exp_f := 49;
        ELSIF x =- 7624 THEN
            exp_f := 49;
        ELSIF x =- 7623 THEN
            exp_f := 50;
        ELSIF x =- 7622 THEN
            exp_f := 50;
        ELSIF x =- 7621 THEN
            exp_f := 50;
        ELSIF x =- 7620 THEN
            exp_f := 50;
        ELSIF x =- 7619 THEN
            exp_f := 50;
        ELSIF x =- 7618 THEN
            exp_f := 50;
        ELSIF x =- 7617 THEN
            exp_f := 50;
        ELSIF x =- 7616 THEN
            exp_f := 50;
        ELSIF x =- 7615 THEN
            exp_f := 50;
        ELSIF x =- 7614 THEN
            exp_f := 50;
        ELSIF x =- 7613 THEN
            exp_f := 50;
        ELSIF x =- 7612 THEN
            exp_f := 50;
        ELSIF x =- 7611 THEN
            exp_f := 50;
        ELSIF x =- 7610 THEN
            exp_f := 50;
        ELSIF x =- 7609 THEN
            exp_f := 50;
        ELSIF x =- 7608 THEN
            exp_f := 50;
        ELSIF x =- 7607 THEN
            exp_f := 50;
        ELSIF x =- 7606 THEN
            exp_f := 50;
        ELSIF x =- 7605 THEN
            exp_f := 50;
        ELSIF x =- 7604 THEN
            exp_f := 50;
        ELSIF x =- 7603 THEN
            exp_f := 50;
        ELSIF x =- 7602 THEN
            exp_f := 50;
        ELSIF x =- 7601 THEN
            exp_f := 50;
        ELSIF x =- 7600 THEN
            exp_f := 50;
        ELSIF x =- 7599 THEN
            exp_f := 50;
        ELSIF x =- 7598 THEN
            exp_f := 50;
        ELSIF x =- 7597 THEN
            exp_f := 50;
        ELSIF x =- 7596 THEN
            exp_f := 50;
        ELSIF x =- 7595 THEN
            exp_f := 50;
        ELSIF x =- 7594 THEN
            exp_f := 50;
        ELSIF x =- 7593 THEN
            exp_f := 50;
        ELSIF x =- 7592 THEN
            exp_f := 50;
        ELSIF x =- 7591 THEN
            exp_f := 50;
        ELSIF x =- 7590 THEN
            exp_f := 50;
        ELSIF x =- 7589 THEN
            exp_f := 50;
        ELSIF x =- 7588 THEN
            exp_f := 50;
        ELSIF x =- 7587 THEN
            exp_f := 50;
        ELSIF x =- 7586 THEN
            exp_f := 50;
        ELSIF x =- 7585 THEN
            exp_f := 51;
        ELSIF x =- 7584 THEN
            exp_f := 51;
        ELSIF x =- 7583 THEN
            exp_f := 51;
        ELSIF x =- 7582 THEN
            exp_f := 51;
        ELSIF x =- 7581 THEN
            exp_f := 51;
        ELSIF x =- 7580 THEN
            exp_f := 51;
        ELSIF x =- 7579 THEN
            exp_f := 51;
        ELSIF x =- 7578 THEN
            exp_f := 51;
        ELSIF x =- 7577 THEN
            exp_f := 51;
        ELSIF x =- 7576 THEN
            exp_f := 51;
        ELSIF x =- 7575 THEN
            exp_f := 51;
        ELSIF x =- 7574 THEN
            exp_f := 51;
        ELSIF x =- 7573 THEN
            exp_f := 51;
        ELSIF x =- 7572 THEN
            exp_f := 51;
        ELSIF x =- 7571 THEN
            exp_f := 51;
        ELSIF x =- 7570 THEN
            exp_f := 51;
        ELSIF x =- 7569 THEN
            exp_f := 51;
        ELSIF x =- 7568 THEN
            exp_f := 51;
        ELSIF x =- 7567 THEN
            exp_f := 51;
        ELSIF x =- 7566 THEN
            exp_f := 51;
        ELSIF x =- 7565 THEN
            exp_f := 51;
        ELSIF x =- 7564 THEN
            exp_f := 51;
        ELSIF x =- 7563 THEN
            exp_f := 51;
        ELSIF x =- 7562 THEN
            exp_f := 51;
        ELSIF x =- 7561 THEN
            exp_f := 51;
        ELSIF x =- 7560 THEN
            exp_f := 51;
        ELSIF x =- 7559 THEN
            exp_f := 51;
        ELSIF x =- 7558 THEN
            exp_f := 51;
        ELSIF x =- 7557 THEN
            exp_f := 51;
        ELSIF x =- 7556 THEN
            exp_f := 51;
        ELSIF x =- 7555 THEN
            exp_f := 51;
        ELSIF x =- 7554 THEN
            exp_f := 51;
        ELSIF x =- 7553 THEN
            exp_f := 51;
        ELSIF x =- 7552 THEN
            exp_f := 51;
        ELSIF x =- 7551 THEN
            exp_f := 51;
        ELSIF x =- 7550 THEN
            exp_f := 51;
        ELSIF x =- 7549 THEN
            exp_f := 51;
        ELSIF x =- 7548 THEN
            exp_f := 51;
        ELSIF x =- 7547 THEN
            exp_f := 52;
        ELSIF x =- 7546 THEN
            exp_f := 52;
        ELSIF x =- 7545 THEN
            exp_f := 52;
        ELSIF x =- 7544 THEN
            exp_f := 52;
        ELSIF x =- 7543 THEN
            exp_f := 52;
        ELSIF x =- 7542 THEN
            exp_f := 52;
        ELSIF x =- 7541 THEN
            exp_f := 52;
        ELSIF x =- 7540 THEN
            exp_f := 52;
        ELSIF x =- 7539 THEN
            exp_f := 52;
        ELSIF x =- 7538 THEN
            exp_f := 52;
        ELSIF x =- 7537 THEN
            exp_f := 52;
        ELSIF x =- 7536 THEN
            exp_f := 52;
        ELSIF x =- 7535 THEN
            exp_f := 52;
        ELSIF x =- 7534 THEN
            exp_f := 52;
        ELSIF x =- 7533 THEN
            exp_f := 52;
        ELSIF x =- 7532 THEN
            exp_f := 52;
        ELSIF x =- 7531 THEN
            exp_f := 52;
        ELSIF x =- 7530 THEN
            exp_f := 52;
        ELSIF x =- 7529 THEN
            exp_f := 52;
        ELSIF x =- 7528 THEN
            exp_f := 52;
        ELSIF x =- 7527 THEN
            exp_f := 52;
        ELSIF x =- 7526 THEN
            exp_f := 52;
        ELSIF x =- 7525 THEN
            exp_f := 52;
        ELSIF x =- 7524 THEN
            exp_f := 52;
        ELSIF x =- 7523 THEN
            exp_f := 52;
        ELSIF x =- 7522 THEN
            exp_f := 52;
        ELSIF x =- 7521 THEN
            exp_f := 52;
        ELSIF x =- 7520 THEN
            exp_f := 52;
        ELSIF x =- 7519 THEN
            exp_f := 52;
        ELSIF x =- 7518 THEN
            exp_f := 52;
        ELSIF x =- 7517 THEN
            exp_f := 52;
        ELSIF x =- 7516 THEN
            exp_f := 52;
        ELSIF x =- 7515 THEN
            exp_f := 52;
        ELSIF x =- 7514 THEN
            exp_f := 52;
        ELSIF x =- 7513 THEN
            exp_f := 52;
        ELSIF x =- 7512 THEN
            exp_f := 52;
        ELSIF x =- 7511 THEN
            exp_f := 52;
        ELSIF x =- 7510 THEN
            exp_f := 52;
        ELSIF x =- 7509 THEN
            exp_f := 53;
        ELSIF x =- 7508 THEN
            exp_f := 53;
        ELSIF x =- 7507 THEN
            exp_f := 53;
        ELSIF x =- 7506 THEN
            exp_f := 53;
        ELSIF x =- 7505 THEN
            exp_f := 53;
        ELSIF x =- 7504 THEN
            exp_f := 53;
        ELSIF x =- 7503 THEN
            exp_f := 53;
        ELSIF x =- 7502 THEN
            exp_f := 53;
        ELSIF x =- 7501 THEN
            exp_f := 53;
        ELSIF x =- 7500 THEN
            exp_f := 53;
        ELSIF x =- 7499 THEN
            exp_f := 53;
        ELSIF x =- 7498 THEN
            exp_f := 53;
        ELSIF x =- 7497 THEN
            exp_f := 53;
        ELSIF x =- 7496 THEN
            exp_f := 53;
        ELSIF x =- 7495 THEN
            exp_f := 53;
        ELSIF x =- 7494 THEN
            exp_f := 53;
        ELSIF x =- 7493 THEN
            exp_f := 53;
        ELSIF x =- 7492 THEN
            exp_f := 53;
        ELSIF x =- 7491 THEN
            exp_f := 53;
        ELSIF x =- 7490 THEN
            exp_f := 53;
        ELSIF x =- 7489 THEN
            exp_f := 53;
        ELSIF x =- 7488 THEN
            exp_f := 53;
        ELSIF x =- 7487 THEN
            exp_f := 53;
        ELSIF x =- 7486 THEN
            exp_f := 53;
        ELSIF x =- 7485 THEN
            exp_f := 53;
        ELSIF x =- 7484 THEN
            exp_f := 53;
        ELSIF x =- 7483 THEN
            exp_f := 53;
        ELSIF x =- 7482 THEN
            exp_f := 53;
        ELSIF x =- 7481 THEN
            exp_f := 53;
        ELSIF x =- 7480 THEN
            exp_f := 53;
        ELSIF x =- 7479 THEN
            exp_f := 53;
        ELSIF x =- 7478 THEN
            exp_f := 53;
        ELSIF x =- 7477 THEN
            exp_f := 53;
        ELSIF x =- 7476 THEN
            exp_f := 53;
        ELSIF x =- 7475 THEN
            exp_f := 53;
        ELSIF x =- 7474 THEN
            exp_f := 53;
        ELSIF x =- 7473 THEN
            exp_f := 53;
        ELSIF x =- 7472 THEN
            exp_f := 53;
        ELSIF x =- 7471 THEN
            exp_f := 54;
        ELSIF x =- 7470 THEN
            exp_f := 54;
        ELSIF x =- 7469 THEN
            exp_f := 54;
        ELSIF x =- 7468 THEN
            exp_f := 54;
        ELSIF x =- 7467 THEN
            exp_f := 54;
        ELSIF x =- 7466 THEN
            exp_f := 54;
        ELSIF x =- 7465 THEN
            exp_f := 54;
        ELSIF x =- 7464 THEN
            exp_f := 54;
        ELSIF x =- 7463 THEN
            exp_f := 54;
        ELSIF x =- 7462 THEN
            exp_f := 54;
        ELSIF x =- 7461 THEN
            exp_f := 54;
        ELSIF x =- 7460 THEN
            exp_f := 54;
        ELSIF x =- 7459 THEN
            exp_f := 54;
        ELSIF x =- 7458 THEN
            exp_f := 54;
        ELSIF x =- 7457 THEN
            exp_f := 54;
        ELSIF x =- 7456 THEN
            exp_f := 54;
        ELSIF x =- 7455 THEN
            exp_f := 54;
        ELSIF x =- 7454 THEN
            exp_f := 54;
        ELSIF x =- 7453 THEN
            exp_f := 54;
        ELSIF x =- 7452 THEN
            exp_f := 54;
        ELSIF x =- 7451 THEN
            exp_f := 54;
        ELSIF x =- 7450 THEN
            exp_f := 54;
        ELSIF x =- 7449 THEN
            exp_f := 54;
        ELSIF x =- 7448 THEN
            exp_f := 54;
        ELSIF x =- 7447 THEN
            exp_f := 54;
        ELSIF x =- 7446 THEN
            exp_f := 54;
        ELSIF x =- 7445 THEN
            exp_f := 54;
        ELSIF x =- 7444 THEN
            exp_f := 54;
        ELSIF x =- 7443 THEN
            exp_f := 54;
        ELSIF x =- 7442 THEN
            exp_f := 54;
        ELSIF x =- 7441 THEN
            exp_f := 54;
        ELSIF x =- 7440 THEN
            exp_f := 54;
        ELSIF x =- 7439 THEN
            exp_f := 54;
        ELSIF x =- 7438 THEN
            exp_f := 54;
        ELSIF x =- 7437 THEN
            exp_f := 54;
        ELSIF x =- 7436 THEN
            exp_f := 54;
        ELSIF x =- 7435 THEN
            exp_f := 54;
        ELSIF x =- 7434 THEN
            exp_f := 54;
        ELSIF x =- 7433 THEN
            exp_f := 55;
        ELSIF x =- 7432 THEN
            exp_f := 55;
        ELSIF x =- 7431 THEN
            exp_f := 55;
        ELSIF x =- 7430 THEN
            exp_f := 55;
        ELSIF x =- 7429 THEN
            exp_f := 55;
        ELSIF x =- 7428 THEN
            exp_f := 55;
        ELSIF x =- 7427 THEN
            exp_f := 55;
        ELSIF x =- 7426 THEN
            exp_f := 55;
        ELSIF x =- 7425 THEN
            exp_f := 55;
        ELSIF x =- 7424 THEN
            exp_f := 55;
        ELSIF x =- 7423 THEN
            exp_f := 55;
        ELSIF x =- 7422 THEN
            exp_f := 55;
        ELSIF x =- 7421 THEN
            exp_f := 55;
        ELSIF x =- 7420 THEN
            exp_f := 55;
        ELSIF x =- 7419 THEN
            exp_f := 55;
        ELSIF x =- 7418 THEN
            exp_f := 55;
        ELSIF x =- 7417 THEN
            exp_f := 55;
        ELSIF x =- 7416 THEN
            exp_f := 55;
        ELSIF x =- 7415 THEN
            exp_f := 55;
        ELSIF x =- 7414 THEN
            exp_f := 55;
        ELSIF x =- 7413 THEN
            exp_f := 55;
        ELSIF x =- 7412 THEN
            exp_f := 55;
        ELSIF x =- 7411 THEN
            exp_f := 55;
        ELSIF x =- 7410 THEN
            exp_f := 55;
        ELSIF x =- 7409 THEN
            exp_f := 55;
        ELSIF x =- 7408 THEN
            exp_f := 55;
        ELSIF x =- 7407 THEN
            exp_f := 55;
        ELSIF x =- 7406 THEN
            exp_f := 55;
        ELSIF x =- 7405 THEN
            exp_f := 55;
        ELSIF x =- 7404 THEN
            exp_f := 55;
        ELSIF x =- 7403 THEN
            exp_f := 55;
        ELSIF x =- 7402 THEN
            exp_f := 55;
        ELSIF x =- 7401 THEN
            exp_f := 55;
        ELSIF x =- 7400 THEN
            exp_f := 55;
        ELSIF x =- 7399 THEN
            exp_f := 55;
        ELSIF x =- 7398 THEN
            exp_f := 55;
        ELSIF x =- 7397 THEN
            exp_f := 55;
        ELSIF x =- 7396 THEN
            exp_f := 55;
        ELSIF x =- 7395 THEN
            exp_f := 56;
        ELSIF x =- 7394 THEN
            exp_f := 56;
        ELSIF x =- 7393 THEN
            exp_f := 56;
        ELSIF x =- 7392 THEN
            exp_f := 56;
        ELSIF x =- 7391 THEN
            exp_f := 56;
        ELSIF x =- 7390 THEN
            exp_f := 56;
        ELSIF x =- 7389 THEN
            exp_f := 56;
        ELSIF x =- 7388 THEN
            exp_f := 56;
        ELSIF x =- 7387 THEN
            exp_f := 56;
        ELSIF x =- 7386 THEN
            exp_f := 56;
        ELSIF x =- 7385 THEN
            exp_f := 56;
        ELSIF x =- 7384 THEN
            exp_f := 56;
        ELSIF x =- 7383 THEN
            exp_f := 56;
        ELSIF x =- 7382 THEN
            exp_f := 56;
        ELSIF x =- 7381 THEN
            exp_f := 56;
        ELSIF x =- 7380 THEN
            exp_f := 56;
        ELSIF x =- 7379 THEN
            exp_f := 56;
        ELSIF x =- 7378 THEN
            exp_f := 56;
        ELSIF x =- 7377 THEN
            exp_f := 56;
        ELSIF x =- 7376 THEN
            exp_f := 56;
        ELSIF x =- 7375 THEN
            exp_f := 56;
        ELSIF x =- 7374 THEN
            exp_f := 56;
        ELSIF x =- 7373 THEN
            exp_f := 56;
        ELSIF x =- 7372 THEN
            exp_f := 56;
        ELSIF x =- 7371 THEN
            exp_f := 56;
        ELSIF x =- 7370 THEN
            exp_f := 56;
        ELSIF x =- 7369 THEN
            exp_f := 56;
        ELSIF x =- 7368 THEN
            exp_f := 56;
        ELSIF x =- 7367 THEN
            exp_f := 56;
        ELSIF x =- 7366 THEN
            exp_f := 56;
        ELSIF x =- 7365 THEN
            exp_f := 56;
        ELSIF x =- 7364 THEN
            exp_f := 56;
        ELSIF x =- 7363 THEN
            exp_f := 56;
        ELSIF x =- 7362 THEN
            exp_f := 56;
        ELSIF x =- 7361 THEN
            exp_f := 56;
        ELSIF x =- 7360 THEN
            exp_f := 56;
        ELSIF x =- 7359 THEN
            exp_f := 56;
        ELSIF x =- 7358 THEN
            exp_f := 56;
        ELSIF x =- 7357 THEN
            exp_f := 57;
        ELSIF x =- 7356 THEN
            exp_f := 57;
        ELSIF x =- 7355 THEN
            exp_f := 57;
        ELSIF x =- 7354 THEN
            exp_f := 57;
        ELSIF x =- 7353 THEN
            exp_f := 57;
        ELSIF x =- 7352 THEN
            exp_f := 57;
        ELSIF x =- 7351 THEN
            exp_f := 57;
        ELSIF x =- 7350 THEN
            exp_f := 57;
        ELSIF x =- 7349 THEN
            exp_f := 57;
        ELSIF x =- 7348 THEN
            exp_f := 57;
        ELSIF x =- 7347 THEN
            exp_f := 57;
        ELSIF x =- 7346 THEN
            exp_f := 57;
        ELSIF x =- 7345 THEN
            exp_f := 57;
        ELSIF x =- 7344 THEN
            exp_f := 57;
        ELSIF x =- 7343 THEN
            exp_f := 57;
        ELSIF x =- 7342 THEN
            exp_f := 57;
        ELSIF x =- 7341 THEN
            exp_f := 57;
        ELSIF x =- 7340 THEN
            exp_f := 57;
        ELSIF x =- 7339 THEN
            exp_f := 57;
        ELSIF x =- 7338 THEN
            exp_f := 57;
        ELSIF x =- 7337 THEN
            exp_f := 57;
        ELSIF x =- 7336 THEN
            exp_f := 57;
        ELSIF x =- 7335 THEN
            exp_f := 57;
        ELSIF x =- 7334 THEN
            exp_f := 57;
        ELSIF x =- 7333 THEN
            exp_f := 57;
        ELSIF x =- 7332 THEN
            exp_f := 57;
        ELSIF x =- 7331 THEN
            exp_f := 57;
        ELSIF x =- 7330 THEN
            exp_f := 57;
        ELSIF x =- 7329 THEN
            exp_f := 57;
        ELSIF x =- 7328 THEN
            exp_f := 57;
        ELSIF x =- 7327 THEN
            exp_f := 57;
        ELSIF x =- 7326 THEN
            exp_f := 57;
        ELSIF x =- 7325 THEN
            exp_f := 57;
        ELSIF x =- 7324 THEN
            exp_f := 57;
        ELSIF x =- 7323 THEN
            exp_f := 57;
        ELSIF x =- 7322 THEN
            exp_f := 57;
        ELSIF x =- 7321 THEN
            exp_f := 57;
        ELSIF x =- 7320 THEN
            exp_f := 57;
        ELSIF x =- 7319 THEN
            exp_f := 58;
        ELSIF x =- 7318 THEN
            exp_f := 58;
        ELSIF x =- 7317 THEN
            exp_f := 58;
        ELSIF x =- 7316 THEN
            exp_f := 58;
        ELSIF x =- 7315 THEN
            exp_f := 58;
        ELSIF x =- 7314 THEN
            exp_f := 58;
        ELSIF x =- 7313 THEN
            exp_f := 58;
        ELSIF x =- 7312 THEN
            exp_f := 58;
        ELSIF x =- 7311 THEN
            exp_f := 58;
        ELSIF x =- 7310 THEN
            exp_f := 58;
        ELSIF x =- 7309 THEN
            exp_f := 58;
        ELSIF x =- 7308 THEN
            exp_f := 58;
        ELSIF x =- 7307 THEN
            exp_f := 58;
        ELSIF x =- 7306 THEN
            exp_f := 58;
        ELSIF x =- 7305 THEN
            exp_f := 58;
        ELSIF x =- 7304 THEN
            exp_f := 58;
        ELSIF x =- 7303 THEN
            exp_f := 58;
        ELSIF x =- 7302 THEN
            exp_f := 58;
        ELSIF x =- 7301 THEN
            exp_f := 58;
        ELSIF x =- 7300 THEN
            exp_f := 58;
        ELSIF x =- 7299 THEN
            exp_f := 58;
        ELSIF x =- 7298 THEN
            exp_f := 58;
        ELSIF x =- 7297 THEN
            exp_f := 58;
        ELSIF x =- 7296 THEN
            exp_f := 58;
        ELSIF x =- 7295 THEN
            exp_f := 58;
        ELSIF x =- 7294 THEN
            exp_f := 58;
        ELSIF x =- 7293 THEN
            exp_f := 58;
        ELSIF x =- 7292 THEN
            exp_f := 58;
        ELSIF x =- 7291 THEN
            exp_f := 58;
        ELSIF x =- 7290 THEN
            exp_f := 58;
        ELSIF x =- 7289 THEN
            exp_f := 58;
        ELSIF x =- 7288 THEN
            exp_f := 58;
        ELSIF x =- 7287 THEN
            exp_f := 58;
        ELSIF x =- 7286 THEN
            exp_f := 58;
        ELSIF x =- 7285 THEN
            exp_f := 58;
        ELSIF x =- 7284 THEN
            exp_f := 58;
        ELSIF x =- 7283 THEN
            exp_f := 58;
        ELSIF x =- 7282 THEN
            exp_f := 58;
        ELSIF x =- 7281 THEN
            exp_f := 59;
        ELSIF x =- 7280 THEN
            exp_f := 59;
        ELSIF x =- 7279 THEN
            exp_f := 59;
        ELSIF x =- 7278 THEN
            exp_f := 59;
        ELSIF x =- 7277 THEN
            exp_f := 59;
        ELSIF x =- 7276 THEN
            exp_f := 59;
        ELSIF x =- 7275 THEN
            exp_f := 59;
        ELSIF x =- 7274 THEN
            exp_f := 59;
        ELSIF x =- 7273 THEN
            exp_f := 59;
        ELSIF x =- 7272 THEN
            exp_f := 59;
        ELSIF x =- 7271 THEN
            exp_f := 59;
        ELSIF x =- 7270 THEN
            exp_f := 59;
        ELSIF x =- 7269 THEN
            exp_f := 59;
        ELSIF x =- 7268 THEN
            exp_f := 59;
        ELSIF x =- 7267 THEN
            exp_f := 59;
        ELSIF x =- 7266 THEN
            exp_f := 59;
        ELSIF x =- 7265 THEN
            exp_f := 59;
        ELSIF x =- 7264 THEN
            exp_f := 59;
        ELSIF x =- 7263 THEN
            exp_f := 59;
        ELSIF x =- 7262 THEN
            exp_f := 59;
        ELSIF x =- 7261 THEN
            exp_f := 59;
        ELSIF x =- 7260 THEN
            exp_f := 59;
        ELSIF x =- 7259 THEN
            exp_f := 59;
        ELSIF x =- 7258 THEN
            exp_f := 59;
        ELSIF x =- 7257 THEN
            exp_f := 59;
        ELSIF x =- 7256 THEN
            exp_f := 59;
        ELSIF x =- 7255 THEN
            exp_f := 59;
        ELSIF x =- 7254 THEN
            exp_f := 59;
        ELSIF x =- 7253 THEN
            exp_f := 59;
        ELSIF x =- 7252 THEN
            exp_f := 59;
        ELSIF x =- 7251 THEN
            exp_f := 59;
        ELSIF x =- 7250 THEN
            exp_f := 59;
        ELSIF x =- 7249 THEN
            exp_f := 59;
        ELSIF x =- 7248 THEN
            exp_f := 59;
        ELSIF x =- 7247 THEN
            exp_f := 59;
        ELSIF x =- 7246 THEN
            exp_f := 59;
        ELSIF x =- 7245 THEN
            exp_f := 59;
        ELSIF x =- 7244 THEN
            exp_f := 59;
        ELSIF x =- 7243 THEN
            exp_f := 60;
        ELSIF x =- 7242 THEN
            exp_f := 60;
        ELSIF x =- 7241 THEN
            exp_f := 60;
        ELSIF x =- 7240 THEN
            exp_f := 60;
        ELSIF x =- 7239 THEN
            exp_f := 60;
        ELSIF x =- 7238 THEN
            exp_f := 60;
        ELSIF x =- 7237 THEN
            exp_f := 60;
        ELSIF x =- 7236 THEN
            exp_f := 60;
        ELSIF x =- 7235 THEN
            exp_f := 60;
        ELSIF x =- 7234 THEN
            exp_f := 60;
        ELSIF x =- 7233 THEN
            exp_f := 60;
        ELSIF x =- 7232 THEN
            exp_f := 60;
        ELSIF x =- 7231 THEN
            exp_f := 60;
        ELSIF x =- 7230 THEN
            exp_f := 60;
        ELSIF x =- 7229 THEN
            exp_f := 60;
        ELSIF x =- 7228 THEN
            exp_f := 60;
        ELSIF x =- 7227 THEN
            exp_f := 60;
        ELSIF x =- 7226 THEN
            exp_f := 60;
        ELSIF x =- 7225 THEN
            exp_f := 60;
        ELSIF x =- 7224 THEN
            exp_f := 60;
        ELSIF x =- 7223 THEN
            exp_f := 60;
        ELSIF x =- 7222 THEN
            exp_f := 60;
        ELSIF x =- 7221 THEN
            exp_f := 60;
        ELSIF x =- 7220 THEN
            exp_f := 60;
        ELSIF x =- 7219 THEN
            exp_f := 60;
        ELSIF x =- 7218 THEN
            exp_f := 60;
        ELSIF x =- 7217 THEN
            exp_f := 60;
        ELSIF x =- 7216 THEN
            exp_f := 60;
        ELSIF x =- 7215 THEN
            exp_f := 60;
        ELSIF x =- 7214 THEN
            exp_f := 60;
        ELSIF x =- 7213 THEN
            exp_f := 60;
        ELSIF x =- 7212 THEN
            exp_f := 60;
        ELSIF x =- 7211 THEN
            exp_f := 60;
        ELSIF x =- 7210 THEN
            exp_f := 60;
        ELSIF x =- 7209 THEN
            exp_f := 60;
        ELSIF x =- 7208 THEN
            exp_f := 60;
        ELSIF x =- 7207 THEN
            exp_f := 60;
        ELSIF x =- 7206 THEN
            exp_f := 60;
        ELSIF x =- 7205 THEN
            exp_f := 61;
        ELSIF x =- 7204 THEN
            exp_f := 61;
        ELSIF x =- 7203 THEN
            exp_f := 61;
        ELSIF x =- 7202 THEN
            exp_f := 61;
        ELSIF x =- 7201 THEN
            exp_f := 61;
        ELSIF x =- 7200 THEN
            exp_f := 61;
        ELSIF x =- 7199 THEN
            exp_f := 61;
        ELSIF x =- 7198 THEN
            exp_f := 61;
        ELSIF x =- 7197 THEN
            exp_f := 61;
        ELSIF x =- 7196 THEN
            exp_f := 61;
        ELSIF x =- 7195 THEN
            exp_f := 61;
        ELSIF x =- 7194 THEN
            exp_f := 61;
        ELSIF x =- 7193 THEN
            exp_f := 61;
        ELSIF x =- 7192 THEN
            exp_f := 61;
        ELSIF x =- 7191 THEN
            exp_f := 61;
        ELSIF x =- 7190 THEN
            exp_f := 61;
        ELSIF x =- 7189 THEN
            exp_f := 61;
        ELSIF x =- 7188 THEN
            exp_f := 61;
        ELSIF x =- 7187 THEN
            exp_f := 61;
        ELSIF x =- 7186 THEN
            exp_f := 61;
        ELSIF x =- 7185 THEN
            exp_f := 61;
        ELSIF x =- 7184 THEN
            exp_f := 61;
        ELSIF x =- 7183 THEN
            exp_f := 61;
        ELSIF x =- 7182 THEN
            exp_f := 61;
        ELSIF x =- 7181 THEN
            exp_f := 61;
        ELSIF x =- 7180 THEN
            exp_f := 61;
        ELSIF x =- 7179 THEN
            exp_f := 61;
        ELSIF x =- 7178 THEN
            exp_f := 61;
        ELSIF x =- 7177 THEN
            exp_f := 61;
        ELSIF x =- 7176 THEN
            exp_f := 61;
        ELSIF x =- 7175 THEN
            exp_f := 61;
        ELSIF x =- 7174 THEN
            exp_f := 61;
        ELSIF x =- 7173 THEN
            exp_f := 61;
        ELSIF x =- 7172 THEN
            exp_f := 61;
        ELSIF x =- 7171 THEN
            exp_f := 61;
        ELSIF x =- 7170 THEN
            exp_f := 61;
        ELSIF x =- 7169 THEN
            exp_f := 61;
        ELSIF x =- 7168 THEN
            exp_f := 61;
        ELSIF x =- 7167 THEN
            exp_f := 62;
        ELSIF x =- 7166 THEN
            exp_f := 62;
        ELSIF x =- 7165 THEN
            exp_f := 62;
        ELSIF x =- 7164 THEN
            exp_f := 62;
        ELSIF x =- 7163 THEN
            exp_f := 62;
        ELSIF x =- 7162 THEN
            exp_f := 62;
        ELSIF x =- 7161 THEN
            exp_f := 62;
        ELSIF x =- 7160 THEN
            exp_f := 62;
        ELSIF x =- 7159 THEN
            exp_f := 62;
        ELSIF x =- 7158 THEN
            exp_f := 62;
        ELSIF x =- 7157 THEN
            exp_f := 62;
        ELSIF x =- 7156 THEN
            exp_f := 62;
        ELSIF x =- 7155 THEN
            exp_f := 62;
        ELSIF x =- 7154 THEN
            exp_f := 62;
        ELSIF x =- 7153 THEN
            exp_f := 62;
        ELSIF x =- 7152 THEN
            exp_f := 62;
        ELSIF x =- 7151 THEN
            exp_f := 62;
        ELSIF x =- 7150 THEN
            exp_f := 62;
        ELSIF x =- 7149 THEN
            exp_f := 62;
        ELSIF x =- 7148 THEN
            exp_f := 62;
        ELSIF x =- 7147 THEN
            exp_f := 62;
        ELSIF x =- 7146 THEN
            exp_f := 62;
        ELSIF x =- 7145 THEN
            exp_f := 62;
        ELSIF x =- 7144 THEN
            exp_f := 62;
        ELSIF x =- 7143 THEN
            exp_f := 62;
        ELSIF x =- 7142 THEN
            exp_f := 62;
        ELSIF x =- 7141 THEN
            exp_f := 62;
        ELSIF x =- 7140 THEN
            exp_f := 62;
        ELSIF x =- 7139 THEN
            exp_f := 62;
        ELSIF x =- 7138 THEN
            exp_f := 62;
        ELSIF x =- 7137 THEN
            exp_f := 62;
        ELSIF x =- 7136 THEN
            exp_f := 62;
        ELSIF x =- 7135 THEN
            exp_f := 63;
        ELSIF x =- 7134 THEN
            exp_f := 63;
        ELSIF x =- 7133 THEN
            exp_f := 63;
        ELSIF x =- 7132 THEN
            exp_f := 63;
        ELSIF x =- 7131 THEN
            exp_f := 63;
        ELSIF x =- 7130 THEN
            exp_f := 63;
        ELSIF x =- 7129 THEN
            exp_f := 63;
        ELSIF x =- 7128 THEN
            exp_f := 63;
        ELSIF x =- 7127 THEN
            exp_f := 63;
        ELSIF x =- 7126 THEN
            exp_f := 63;
        ELSIF x =- 7125 THEN
            exp_f := 63;
        ELSIF x =- 7124 THEN
            exp_f := 63;
        ELSIF x =- 7123 THEN
            exp_f := 63;
        ELSIF x =- 7122 THEN
            exp_f := 63;
        ELSIF x =- 7121 THEN
            exp_f := 63;
        ELSIF x =- 7120 THEN
            exp_f := 63;
        ELSIF x =- 7119 THEN
            exp_f := 63;
        ELSIF x =- 7118 THEN
            exp_f := 63;
        ELSIF x =- 7117 THEN
            exp_f := 63;
        ELSIF x =- 7116 THEN
            exp_f := 63;
        ELSIF x =- 7115 THEN
            exp_f := 63;
        ELSIF x =- 7114 THEN
            exp_f := 63;
        ELSIF x =- 7113 THEN
            exp_f := 63;
        ELSIF x =- 7112 THEN
            exp_f := 63;
        ELSIF x =- 7111 THEN
            exp_f := 63;
        ELSIF x =- 7110 THEN
            exp_f := 63;
        ELSIF x =- 7109 THEN
            exp_f := 63;
        ELSIF x =- 7108 THEN
            exp_f := 63;
        ELSIF x =- 7107 THEN
            exp_f := 63;
        ELSIF x =- 7106 THEN
            exp_f := 63;
        ELSIF x =- 7105 THEN
            exp_f := 63;
        ELSIF x =- 7104 THEN
            exp_f := 63;
        ELSIF x =- 7103 THEN
            exp_f := 64;
        ELSIF x =- 7102 THEN
            exp_f := 64;
        ELSIF x =- 7101 THEN
            exp_f := 64;
        ELSIF x =- 7100 THEN
            exp_f := 64;
        ELSIF x =- 7099 THEN
            exp_f := 64;
        ELSIF x =- 7098 THEN
            exp_f := 64;
        ELSIF x =- 7097 THEN
            exp_f := 64;
        ELSIF x =- 7096 THEN
            exp_f := 64;
        ELSIF x =- 7095 THEN
            exp_f := 64;
        ELSIF x =- 7094 THEN
            exp_f := 64;
        ELSIF x =- 7093 THEN
            exp_f := 64;
        ELSIF x =- 7092 THEN
            exp_f := 64;
        ELSIF x =- 7091 THEN
            exp_f := 64;
        ELSIF x =- 7090 THEN
            exp_f := 64;
        ELSIF x =- 7089 THEN
            exp_f := 64;
        ELSIF x =- 7088 THEN
            exp_f := 64;
        ELSIF x =- 7087 THEN
            exp_f := 64;
        ELSIF x =- 7086 THEN
            exp_f := 64;
        ELSIF x =- 7085 THEN
            exp_f := 64;
        ELSIF x =- 7084 THEN
            exp_f := 64;
        ELSIF x =- 7083 THEN
            exp_f := 64;
        ELSIF x =- 7082 THEN
            exp_f := 64;
        ELSIF x =- 7081 THEN
            exp_f := 64;
        ELSIF x =- 7080 THEN
            exp_f := 64;
        ELSIF x =- 7079 THEN
            exp_f := 64;
        ELSIF x =- 7078 THEN
            exp_f := 64;
        ELSIF x =- 7077 THEN
            exp_f := 64;
        ELSIF x =- 7076 THEN
            exp_f := 64;
        ELSIF x =- 7075 THEN
            exp_f := 64;
        ELSIF x =- 7074 THEN
            exp_f := 64;
        ELSIF x =- 7073 THEN
            exp_f := 64;
        ELSIF x =- 7072 THEN
            exp_f := 64;
        ELSIF x =- 7071 THEN
            exp_f := 66;
        ELSIF x =- 7070 THEN
            exp_f := 66;
        ELSIF x =- 7069 THEN
            exp_f := 66;
        ELSIF x =- 7068 THEN
            exp_f := 66;
        ELSIF x =- 7067 THEN
            exp_f := 66;
        ELSIF x =- 7066 THEN
            exp_f := 66;
        ELSIF x =- 7065 THEN
            exp_f := 66;
        ELSIF x =- 7064 THEN
            exp_f := 66;
        ELSIF x =- 7063 THEN
            exp_f := 66;
        ELSIF x =- 7062 THEN
            exp_f := 66;
        ELSIF x =- 7061 THEN
            exp_f := 66;
        ELSIF x =- 7060 THEN
            exp_f := 66;
        ELSIF x =- 7059 THEN
            exp_f := 66;
        ELSIF x =- 7058 THEN
            exp_f := 66;
        ELSIF x =- 7057 THEN
            exp_f := 66;
        ELSIF x =- 7056 THEN
            exp_f := 66;
        ELSIF x =- 7055 THEN
            exp_f := 66;
        ELSIF x =- 7054 THEN
            exp_f := 66;
        ELSIF x =- 7053 THEN
            exp_f := 66;
        ELSIF x =- 7052 THEN
            exp_f := 66;
        ELSIF x =- 7051 THEN
            exp_f := 66;
        ELSIF x =- 7050 THEN
            exp_f := 66;
        ELSIF x =- 7049 THEN
            exp_f := 66;
        ELSIF x =- 7048 THEN
            exp_f := 66;
        ELSIF x =- 7047 THEN
            exp_f := 66;
        ELSIF x =- 7046 THEN
            exp_f := 66;
        ELSIF x =- 7045 THEN
            exp_f := 66;
        ELSIF x =- 7044 THEN
            exp_f := 66;
        ELSIF x =- 7043 THEN
            exp_f := 66;
        ELSIF x =- 7042 THEN
            exp_f := 66;
        ELSIF x =- 7041 THEN
            exp_f := 66;
        ELSIF x =- 7040 THEN
            exp_f := 66;
        ELSIF x =- 7039 THEN
            exp_f := 67;
        ELSIF x =- 7038 THEN
            exp_f := 67;
        ELSIF x =- 7037 THEN
            exp_f := 67;
        ELSIF x =- 7036 THEN
            exp_f := 67;
        ELSIF x =- 7035 THEN
            exp_f := 67;
        ELSIF x =- 7034 THEN
            exp_f := 67;
        ELSIF x =- 7033 THEN
            exp_f := 67;
        ELSIF x =- 7032 THEN
            exp_f := 67;
        ELSIF x =- 7031 THEN
            exp_f := 67;
        ELSIF x =- 7030 THEN
            exp_f := 67;
        ELSIF x =- 7029 THEN
            exp_f := 67;
        ELSIF x =- 7028 THEN
            exp_f := 67;
        ELSIF x =- 7027 THEN
            exp_f := 67;
        ELSIF x =- 7026 THEN
            exp_f := 67;
        ELSIF x =- 7025 THEN
            exp_f := 67;
        ELSIF x =- 7024 THEN
            exp_f := 67;
        ELSIF x =- 7023 THEN
            exp_f := 67;
        ELSIF x =- 7022 THEN
            exp_f := 67;
        ELSIF x =- 7021 THEN
            exp_f := 67;
        ELSIF x =- 7020 THEN
            exp_f := 67;
        ELSIF x =- 7019 THEN
            exp_f := 67;
        ELSIF x =- 7018 THEN
            exp_f := 67;
        ELSIF x =- 7017 THEN
            exp_f := 67;
        ELSIF x =- 7016 THEN
            exp_f := 67;
        ELSIF x =- 7015 THEN
            exp_f := 67;
        ELSIF x =- 7014 THEN
            exp_f := 67;
        ELSIF x =- 7013 THEN
            exp_f := 67;
        ELSIF x =- 7012 THEN
            exp_f := 67;
        ELSIF x =- 7011 THEN
            exp_f := 67;
        ELSIF x =- 7010 THEN
            exp_f := 67;
        ELSIF x =- 7009 THEN
            exp_f := 67;
        ELSIF x =- 7008 THEN
            exp_f := 67;
        ELSIF x =- 7007 THEN
            exp_f := 68;
        ELSIF x =- 7006 THEN
            exp_f := 68;
        ELSIF x =- 7005 THEN
            exp_f := 68;
        ELSIF x =- 7004 THEN
            exp_f := 68;
        ELSIF x =- 7003 THEN
            exp_f := 68;
        ELSIF x =- 7002 THEN
            exp_f := 68;
        ELSIF x =- 7001 THEN
            exp_f := 68;
        ELSIF x =- 7000 THEN
            exp_f := 68;
        ELSIF x =- 6999 THEN
            exp_f := 68;
        ELSIF x =- 6998 THEN
            exp_f := 68;
        ELSIF x =- 6997 THEN
            exp_f := 68;
        ELSIF x =- 6996 THEN
            exp_f := 68;
        ELSIF x =- 6995 THEN
            exp_f := 68;
        ELSIF x =- 6994 THEN
            exp_f := 68;
        ELSIF x =- 6993 THEN
            exp_f := 68;
        ELSIF x =- 6992 THEN
            exp_f := 68;
        ELSIF x =- 6991 THEN
            exp_f := 68;
        ELSIF x =- 6990 THEN
            exp_f := 68;
        ELSIF x =- 6989 THEN
            exp_f := 68;
        ELSIF x =- 6988 THEN
            exp_f := 68;
        ELSIF x =- 6987 THEN
            exp_f := 68;
        ELSIF x =- 6986 THEN
            exp_f := 68;
        ELSIF x =- 6985 THEN
            exp_f := 68;
        ELSIF x =- 6984 THEN
            exp_f := 68;
        ELSIF x =- 6983 THEN
            exp_f := 68;
        ELSIF x =- 6982 THEN
            exp_f := 68;
        ELSIF x =- 6981 THEN
            exp_f := 68;
        ELSIF x =- 6980 THEN
            exp_f := 68;
        ELSIF x =- 6979 THEN
            exp_f := 68;
        ELSIF x =- 6978 THEN
            exp_f := 68;
        ELSIF x =- 6977 THEN
            exp_f := 68;
        ELSIF x =- 6976 THEN
            exp_f := 68;
        ELSIF x =- 6975 THEN
            exp_f := 69;
        ELSIF x =- 6974 THEN
            exp_f := 69;
        ELSIF x =- 6973 THEN
            exp_f := 69;
        ELSIF x =- 6972 THEN
            exp_f := 69;
        ELSIF x =- 6971 THEN
            exp_f := 69;
        ELSIF x =- 6970 THEN
            exp_f := 69;
        ELSIF x =- 6969 THEN
            exp_f := 69;
        ELSIF x =- 6968 THEN
            exp_f := 69;
        ELSIF x =- 6967 THEN
            exp_f := 69;
        ELSIF x =- 6966 THEN
            exp_f := 69;
        ELSIF x =- 6965 THEN
            exp_f := 69;
        ELSIF x =- 6964 THEN
            exp_f := 69;
        ELSIF x =- 6963 THEN
            exp_f := 69;
        ELSIF x =- 6962 THEN
            exp_f := 69;
        ELSIF x =- 6961 THEN
            exp_f := 69;
        ELSIF x =- 6960 THEN
            exp_f := 69;
        ELSIF x =- 6959 THEN
            exp_f := 69;
        ELSIF x =- 6958 THEN
            exp_f := 69;
        ELSIF x =- 6957 THEN
            exp_f := 69;
        ELSIF x =- 6956 THEN
            exp_f := 69;
        ELSIF x =- 6955 THEN
            exp_f := 69;
        ELSIF x =- 6954 THEN
            exp_f := 69;
        ELSIF x =- 6953 THEN
            exp_f := 69;
        ELSIF x =- 6952 THEN
            exp_f := 69;
        ELSIF x =- 6951 THEN
            exp_f := 69;
        ELSIF x =- 6950 THEN
            exp_f := 69;
        ELSIF x =- 6949 THEN
            exp_f := 69;
        ELSIF x =- 6948 THEN
            exp_f := 69;
        ELSIF x =- 6947 THEN
            exp_f := 69;
        ELSIF x =- 6946 THEN
            exp_f := 69;
        ELSIF x =- 6945 THEN
            exp_f := 69;
        ELSIF x =- 6944 THEN
            exp_f := 69;
        ELSIF x =- 6943 THEN
            exp_f := 70;
        ELSIF x =- 6942 THEN
            exp_f := 70;
        ELSIF x =- 6941 THEN
            exp_f := 70;
        ELSIF x =- 6940 THEN
            exp_f := 70;
        ELSIF x =- 6939 THEN
            exp_f := 70;
        ELSIF x =- 6938 THEN
            exp_f := 70;
        ELSIF x =- 6937 THEN
            exp_f := 70;
        ELSIF x =- 6936 THEN
            exp_f := 70;
        ELSIF x =- 6935 THEN
            exp_f := 70;
        ELSIF x =- 6934 THEN
            exp_f := 70;
        ELSIF x =- 6933 THEN
            exp_f := 70;
        ELSIF x =- 6932 THEN
            exp_f := 70;
        ELSIF x =- 6931 THEN
            exp_f := 70;
        ELSIF x =- 6930 THEN
            exp_f := 70;
        ELSIF x =- 6929 THEN
            exp_f := 70;
        ELSIF x =- 6928 THEN
            exp_f := 70;
        ELSIF x =- 6927 THEN
            exp_f := 70;
        ELSIF x =- 6926 THEN
            exp_f := 70;
        ELSIF x =- 6925 THEN
            exp_f := 70;
        ELSIF x =- 6924 THEN
            exp_f := 70;
        ELSIF x =- 6923 THEN
            exp_f := 70;
        ELSIF x =- 6922 THEN
            exp_f := 70;
        ELSIF x =- 6921 THEN
            exp_f := 70;
        ELSIF x =- 6920 THEN
            exp_f := 70;
        ELSIF x =- 6919 THEN
            exp_f := 70;
        ELSIF x =- 6918 THEN
            exp_f := 70;
        ELSIF x =- 6917 THEN
            exp_f := 70;
        ELSIF x =- 6916 THEN
            exp_f := 70;
        ELSIF x =- 6915 THEN
            exp_f := 70;
        ELSIF x =- 6914 THEN
            exp_f := 70;
        ELSIF x =- 6913 THEN
            exp_f := 70;
        ELSIF x =- 6912 THEN
            exp_f := 70;
        ELSIF x =- 6911 THEN
            exp_f := 71;
        ELSIF x =- 6910 THEN
            exp_f := 71;
        ELSIF x =- 6909 THEN
            exp_f := 71;
        ELSIF x =- 6908 THEN
            exp_f := 71;
        ELSIF x =- 6907 THEN
            exp_f := 71;
        ELSIF x =- 6906 THEN
            exp_f := 71;
        ELSIF x =- 6905 THEN
            exp_f := 71;
        ELSIF x =- 6904 THEN
            exp_f := 71;
        ELSIF x =- 6903 THEN
            exp_f := 71;
        ELSIF x =- 6902 THEN
            exp_f := 71;
        ELSIF x =- 6901 THEN
            exp_f := 71;
        ELSIF x =- 6900 THEN
            exp_f := 71;
        ELSIF x =- 6899 THEN
            exp_f := 71;
        ELSIF x =- 6898 THEN
            exp_f := 71;
        ELSIF x =- 6897 THEN
            exp_f := 71;
        ELSIF x =- 6896 THEN
            exp_f := 71;
        ELSIF x =- 6895 THEN
            exp_f := 71;
        ELSIF x =- 6894 THEN
            exp_f := 71;
        ELSIF x =- 6893 THEN
            exp_f := 71;
        ELSIF x =- 6892 THEN
            exp_f := 71;
        ELSIF x =- 6891 THEN
            exp_f := 71;
        ELSIF x =- 6890 THEN
            exp_f := 71;
        ELSIF x =- 6889 THEN
            exp_f := 71;
        ELSIF x =- 6888 THEN
            exp_f := 71;
        ELSIF x =- 6887 THEN
            exp_f := 71;
        ELSIF x =- 6886 THEN
            exp_f := 71;
        ELSIF x =- 6885 THEN
            exp_f := 71;
        ELSIF x =- 6884 THEN
            exp_f := 71;
        ELSIF x =- 6883 THEN
            exp_f := 71;
        ELSIF x =- 6882 THEN
            exp_f := 71;
        ELSIF x =- 6881 THEN
            exp_f := 71;
        ELSIF x =- 6880 THEN
            exp_f := 71;
        ELSIF x =- 6879 THEN
            exp_f := 72;
        ELSIF x =- 6878 THEN
            exp_f := 72;
        ELSIF x =- 6877 THEN
            exp_f := 72;
        ELSIF x =- 6876 THEN
            exp_f := 72;
        ELSIF x =- 6875 THEN
            exp_f := 72;
        ELSIF x =- 6874 THEN
            exp_f := 72;
        ELSIF x =- 6873 THEN
            exp_f := 72;
        ELSIF x =- 6872 THEN
            exp_f := 72;
        ELSIF x =- 6871 THEN
            exp_f := 72;
        ELSIF x =- 6870 THEN
            exp_f := 72;
        ELSIF x =- 6869 THEN
            exp_f := 72;
        ELSIF x =- 6868 THEN
            exp_f := 72;
        ELSIF x =- 6867 THEN
            exp_f := 72;
        ELSIF x =- 6866 THEN
            exp_f := 72;
        ELSIF x =- 6865 THEN
            exp_f := 72;
        ELSIF x =- 6864 THEN
            exp_f := 72;
        ELSIF x =- 6863 THEN
            exp_f := 72;
        ELSIF x =- 6862 THEN
            exp_f := 72;
        ELSIF x =- 6861 THEN
            exp_f := 72;
        ELSIF x =- 6860 THEN
            exp_f := 72;
        ELSIF x =- 6859 THEN
            exp_f := 72;
        ELSIF x =- 6858 THEN
            exp_f := 72;
        ELSIF x =- 6857 THEN
            exp_f := 72;
        ELSIF x =- 6856 THEN
            exp_f := 72;
        ELSIF x =- 6855 THEN
            exp_f := 72;
        ELSIF x =- 6854 THEN
            exp_f := 72;
        ELSIF x =- 6853 THEN
            exp_f := 72;
        ELSIF x =- 6852 THEN
            exp_f := 72;
        ELSIF x =- 6851 THEN
            exp_f := 72;
        ELSIF x =- 6850 THEN
            exp_f := 72;
        ELSIF x =- 6849 THEN
            exp_f := 72;
        ELSIF x =- 6848 THEN
            exp_f := 72;
        ELSIF x =- 6847 THEN
            exp_f := 73;
        ELSIF x =- 6846 THEN
            exp_f := 73;
        ELSIF x =- 6845 THEN
            exp_f := 73;
        ELSIF x =- 6844 THEN
            exp_f := 73;
        ELSIF x =- 6843 THEN
            exp_f := 73;
        ELSIF x =- 6842 THEN
            exp_f := 73;
        ELSIF x =- 6841 THEN
            exp_f := 73;
        ELSIF x =- 6840 THEN
            exp_f := 73;
        ELSIF x =- 6839 THEN
            exp_f := 73;
        ELSIF x =- 6838 THEN
            exp_f := 73;
        ELSIF x =- 6837 THEN
            exp_f := 73;
        ELSIF x =- 6836 THEN
            exp_f := 73;
        ELSIF x =- 6835 THEN
            exp_f := 73;
        ELSIF x =- 6834 THEN
            exp_f := 73;
        ELSIF x =- 6833 THEN
            exp_f := 73;
        ELSIF x =- 6832 THEN
            exp_f := 73;
        ELSIF x =- 6831 THEN
            exp_f := 73;
        ELSIF x =- 6830 THEN
            exp_f := 73;
        ELSIF x =- 6829 THEN
            exp_f := 73;
        ELSIF x =- 6828 THEN
            exp_f := 73;
        ELSIF x =- 6827 THEN
            exp_f := 73;
        ELSIF x =- 6826 THEN
            exp_f := 73;
        ELSIF x =- 6825 THEN
            exp_f := 73;
        ELSIF x =- 6824 THEN
            exp_f := 73;
        ELSIF x =- 6823 THEN
            exp_f := 73;
        ELSIF x =- 6822 THEN
            exp_f := 73;
        ELSIF x =- 6821 THEN
            exp_f := 73;
        ELSIF x =- 6820 THEN
            exp_f := 73;
        ELSIF x =- 6819 THEN
            exp_f := 73;
        ELSIF x =- 6818 THEN
            exp_f := 73;
        ELSIF x =- 6817 THEN
            exp_f := 73;
        ELSIF x =- 6816 THEN
            exp_f := 73;
        ELSIF x =- 6815 THEN
            exp_f := 74;
        ELSIF x =- 6814 THEN
            exp_f := 74;
        ELSIF x =- 6813 THEN
            exp_f := 74;
        ELSIF x =- 6812 THEN
            exp_f := 74;
        ELSIF x =- 6811 THEN
            exp_f := 74;
        ELSIF x =- 6810 THEN
            exp_f := 74;
        ELSIF x =- 6809 THEN
            exp_f := 74;
        ELSIF x =- 6808 THEN
            exp_f := 74;
        ELSIF x =- 6807 THEN
            exp_f := 74;
        ELSIF x =- 6806 THEN
            exp_f := 74;
        ELSIF x =- 6805 THEN
            exp_f := 74;
        ELSIF x =- 6804 THEN
            exp_f := 74;
        ELSIF x =- 6803 THEN
            exp_f := 74;
        ELSIF x =- 6802 THEN
            exp_f := 74;
        ELSIF x =- 6801 THEN
            exp_f := 74;
        ELSIF x =- 6800 THEN
            exp_f := 74;
        ELSIF x =- 6799 THEN
            exp_f := 74;
        ELSIF x =- 6798 THEN
            exp_f := 74;
        ELSIF x =- 6797 THEN
            exp_f := 74;
        ELSIF x =- 6796 THEN
            exp_f := 74;
        ELSIF x =- 6795 THEN
            exp_f := 74;
        ELSIF x =- 6794 THEN
            exp_f := 74;
        ELSIF x =- 6793 THEN
            exp_f := 74;
        ELSIF x =- 6792 THEN
            exp_f := 74;
        ELSIF x =- 6791 THEN
            exp_f := 74;
        ELSIF x =- 6790 THEN
            exp_f := 74;
        ELSIF x =- 6789 THEN
            exp_f := 74;
        ELSIF x =- 6788 THEN
            exp_f := 74;
        ELSIF x =- 6787 THEN
            exp_f := 74;
        ELSIF x =- 6786 THEN
            exp_f := 74;
        ELSIF x =- 6785 THEN
            exp_f := 74;
        ELSIF x =- 6784 THEN
            exp_f := 74;
        ELSIF x =- 6783 THEN
            exp_f := 75;
        ELSIF x =- 6782 THEN
            exp_f := 75;
        ELSIF x =- 6781 THEN
            exp_f := 75;
        ELSIF x =- 6780 THEN
            exp_f := 75;
        ELSIF x =- 6779 THEN
            exp_f := 75;
        ELSIF x =- 6778 THEN
            exp_f := 75;
        ELSIF x =- 6777 THEN
            exp_f := 75;
        ELSIF x =- 6776 THEN
            exp_f := 75;
        ELSIF x =- 6775 THEN
            exp_f := 75;
        ELSIF x =- 6774 THEN
            exp_f := 75;
        ELSIF x =- 6773 THEN
            exp_f := 75;
        ELSIF x =- 6772 THEN
            exp_f := 75;
        ELSIF x =- 6771 THEN
            exp_f := 75;
        ELSIF x =- 6770 THEN
            exp_f := 75;
        ELSIF x =- 6769 THEN
            exp_f := 75;
        ELSIF x =- 6768 THEN
            exp_f := 75;
        ELSIF x =- 6767 THEN
            exp_f := 75;
        ELSIF x =- 6766 THEN
            exp_f := 75;
        ELSIF x =- 6765 THEN
            exp_f := 75;
        ELSIF x =- 6764 THEN
            exp_f := 75;
        ELSIF x =- 6763 THEN
            exp_f := 75;
        ELSIF x =- 6762 THEN
            exp_f := 75;
        ELSIF x =- 6761 THEN
            exp_f := 75;
        ELSIF x =- 6760 THEN
            exp_f := 75;
        ELSIF x =- 6759 THEN
            exp_f := 75;
        ELSIF x =- 6758 THEN
            exp_f := 75;
        ELSIF x =- 6757 THEN
            exp_f := 75;
        ELSIF x =- 6756 THEN
            exp_f := 75;
        ELSIF x =- 6755 THEN
            exp_f := 75;
        ELSIF x =- 6754 THEN
            exp_f := 75;
        ELSIF x =- 6753 THEN
            exp_f := 75;
        ELSIF x =- 6752 THEN
            exp_f := 75;
        ELSIF x =- 6751 THEN
            exp_f := 76;
        ELSIF x =- 6750 THEN
            exp_f := 76;
        ELSIF x =- 6749 THEN
            exp_f := 76;
        ELSIF x =- 6748 THEN
            exp_f := 76;
        ELSIF x =- 6747 THEN
            exp_f := 76;
        ELSIF x =- 6746 THEN
            exp_f := 76;
        ELSIF x =- 6745 THEN
            exp_f := 76;
        ELSIF x =- 6744 THEN
            exp_f := 76;
        ELSIF x =- 6743 THEN
            exp_f := 76;
        ELSIF x =- 6742 THEN
            exp_f := 76;
        ELSIF x =- 6741 THEN
            exp_f := 76;
        ELSIF x =- 6740 THEN
            exp_f := 76;
        ELSIF x =- 6739 THEN
            exp_f := 76;
        ELSIF x =- 6738 THEN
            exp_f := 76;
        ELSIF x =- 6737 THEN
            exp_f := 76;
        ELSIF x =- 6736 THEN
            exp_f := 76;
        ELSIF x =- 6735 THEN
            exp_f := 76;
        ELSIF x =- 6734 THEN
            exp_f := 76;
        ELSIF x =- 6733 THEN
            exp_f := 76;
        ELSIF x =- 6732 THEN
            exp_f := 76;
        ELSIF x =- 6731 THEN
            exp_f := 76;
        ELSIF x =- 6730 THEN
            exp_f := 76;
        ELSIF x =- 6729 THEN
            exp_f := 76;
        ELSIF x =- 6728 THEN
            exp_f := 76;
        ELSIF x =- 6727 THEN
            exp_f := 76;
        ELSIF x =- 6726 THEN
            exp_f := 76;
        ELSIF x =- 6725 THEN
            exp_f := 76;
        ELSIF x =- 6724 THEN
            exp_f := 76;
        ELSIF x =- 6723 THEN
            exp_f := 76;
        ELSIF x =- 6722 THEN
            exp_f := 76;
        ELSIF x =- 6721 THEN
            exp_f := 76;
        ELSIF x =- 6720 THEN
            exp_f := 76;
        ELSIF x =- 6719 THEN
            exp_f := 77;
        ELSIF x =- 6718 THEN
            exp_f := 77;
        ELSIF x =- 6717 THEN
            exp_f := 77;
        ELSIF x =- 6716 THEN
            exp_f := 77;
        ELSIF x =- 6715 THEN
            exp_f := 77;
        ELSIF x =- 6714 THEN
            exp_f := 77;
        ELSIF x =- 6713 THEN
            exp_f := 77;
        ELSIF x =- 6712 THEN
            exp_f := 77;
        ELSIF x =- 6711 THEN
            exp_f := 77;
        ELSIF x =- 6710 THEN
            exp_f := 77;
        ELSIF x =- 6709 THEN
            exp_f := 77;
        ELSIF x =- 6708 THEN
            exp_f := 77;
        ELSIF x =- 6707 THEN
            exp_f := 77;
        ELSIF x =- 6706 THEN
            exp_f := 77;
        ELSIF x =- 6705 THEN
            exp_f := 77;
        ELSIF x =- 6704 THEN
            exp_f := 77;
        ELSIF x =- 6703 THEN
            exp_f := 77;
        ELSIF x =- 6702 THEN
            exp_f := 77;
        ELSIF x =- 6701 THEN
            exp_f := 77;
        ELSIF x =- 6700 THEN
            exp_f := 77;
        ELSIF x =- 6699 THEN
            exp_f := 77;
        ELSIF x =- 6698 THEN
            exp_f := 77;
        ELSIF x =- 6697 THEN
            exp_f := 77;
        ELSIF x =- 6696 THEN
            exp_f := 77;
        ELSIF x =- 6695 THEN
            exp_f := 77;
        ELSIF x =- 6694 THEN
            exp_f := 77;
        ELSIF x =- 6693 THEN
            exp_f := 77;
        ELSIF x =- 6692 THEN
            exp_f := 77;
        ELSIF x =- 6691 THEN
            exp_f := 77;
        ELSIF x =- 6690 THEN
            exp_f := 77;
        ELSIF x =- 6689 THEN
            exp_f := 77;
        ELSIF x =- 6688 THEN
            exp_f := 77;
        ELSIF x =- 6687 THEN
            exp_f := 78;
        ELSIF x =- 6686 THEN
            exp_f := 78;
        ELSIF x =- 6685 THEN
            exp_f := 78;
        ELSIF x =- 6684 THEN
            exp_f := 78;
        ELSIF x =- 6683 THEN
            exp_f := 78;
        ELSIF x =- 6682 THEN
            exp_f := 78;
        ELSIF x =- 6681 THEN
            exp_f := 78;
        ELSIF x =- 6680 THEN
            exp_f := 78;
        ELSIF x =- 6679 THEN
            exp_f := 78;
        ELSIF x =- 6678 THEN
            exp_f := 78;
        ELSIF x =- 6677 THEN
            exp_f := 78;
        ELSIF x =- 6676 THEN
            exp_f := 78;
        ELSIF x =- 6675 THEN
            exp_f := 78;
        ELSIF x =- 6674 THEN
            exp_f := 78;
        ELSIF x =- 6673 THEN
            exp_f := 78;
        ELSIF x =- 6672 THEN
            exp_f := 78;
        ELSIF x =- 6671 THEN
            exp_f := 78;
        ELSIF x =- 6670 THEN
            exp_f := 78;
        ELSIF x =- 6669 THEN
            exp_f := 78;
        ELSIF x =- 6668 THEN
            exp_f := 78;
        ELSIF x =- 6667 THEN
            exp_f := 78;
        ELSIF x =- 6666 THEN
            exp_f := 78;
        ELSIF x =- 6665 THEN
            exp_f := 78;
        ELSIF x =- 6664 THEN
            exp_f := 78;
        ELSIF x =- 6663 THEN
            exp_f := 78;
        ELSIF x =- 6662 THEN
            exp_f := 78;
        ELSIF x =- 6661 THEN
            exp_f := 78;
        ELSIF x =- 6660 THEN
            exp_f := 78;
        ELSIF x =- 6659 THEN
            exp_f := 78;
        ELSIF x =- 6658 THEN
            exp_f := 78;
        ELSIF x =- 6657 THEN
            exp_f := 78;
        ELSIF x =- 6656 THEN
            exp_f := 78;
        ELSIF x =- 6655 THEN
            exp_f := 80;
        ELSIF x =- 6654 THEN
            exp_f := 80;
        ELSIF x =- 6653 THEN
            exp_f := 80;
        ELSIF x =- 6652 THEN
            exp_f := 80;
        ELSIF x =- 6651 THEN
            exp_f := 80;
        ELSIF x =- 6650 THEN
            exp_f := 80;
        ELSIF x =- 6649 THEN
            exp_f := 80;
        ELSIF x =- 6648 THEN
            exp_f := 80;
        ELSIF x =- 6647 THEN
            exp_f := 80;
        ELSIF x =- 6646 THEN
            exp_f := 80;
        ELSIF x =- 6645 THEN
            exp_f := 80;
        ELSIF x =- 6644 THEN
            exp_f := 80;
        ELSIF x =- 6643 THEN
            exp_f := 80;
        ELSIF x =- 6642 THEN
            exp_f := 80;
        ELSIF x =- 6641 THEN
            exp_f := 80;
        ELSIF x =- 6640 THEN
            exp_f := 80;
        ELSIF x =- 6639 THEN
            exp_f := 80;
        ELSIF x =- 6638 THEN
            exp_f := 80;
        ELSIF x =- 6637 THEN
            exp_f := 80;
        ELSIF x =- 6636 THEN
            exp_f := 80;
        ELSIF x =- 6635 THEN
            exp_f := 80;
        ELSIF x =- 6634 THEN
            exp_f := 80;
        ELSIF x =- 6633 THEN
            exp_f := 80;
        ELSIF x =- 6632 THEN
            exp_f := 80;
        ELSIF x =- 6631 THEN
            exp_f := 81;
        ELSIF x =- 6630 THEN
            exp_f := 81;
        ELSIF x =- 6629 THEN
            exp_f := 81;
        ELSIF x =- 6628 THEN
            exp_f := 81;
        ELSIF x =- 6627 THEN
            exp_f := 81;
        ELSIF x =- 6626 THEN
            exp_f := 81;
        ELSIF x =- 6625 THEN
            exp_f := 81;
        ELSIF x =- 6624 THEN
            exp_f := 81;
        ELSIF x =- 6623 THEN
            exp_f := 81;
        ELSIF x =- 6622 THEN
            exp_f := 81;
        ELSIF x =- 6621 THEN
            exp_f := 81;
        ELSIF x =- 6620 THEN
            exp_f := 81;
        ELSIF x =- 6619 THEN
            exp_f := 81;
        ELSIF x =- 6618 THEN
            exp_f := 81;
        ELSIF x =- 6617 THEN
            exp_f := 81;
        ELSIF x =- 6616 THEN
            exp_f := 81;
        ELSIF x =- 6615 THEN
            exp_f := 81;
        ELSIF x =- 6614 THEN
            exp_f := 81;
        ELSIF x =- 6613 THEN
            exp_f := 81;
        ELSIF x =- 6612 THEN
            exp_f := 81;
        ELSIF x =- 6611 THEN
            exp_f := 81;
        ELSIF x =- 6610 THEN
            exp_f := 81;
        ELSIF x =- 6609 THEN
            exp_f := 81;
        ELSIF x =- 6608 THEN
            exp_f := 81;
        ELSIF x =- 6607 THEN
            exp_f := 82;
        ELSIF x =- 6606 THEN
            exp_f := 82;
        ELSIF x =- 6605 THEN
            exp_f := 82;
        ELSIF x =- 6604 THEN
            exp_f := 82;
        ELSIF x =- 6603 THEN
            exp_f := 82;
        ELSIF x =- 6602 THEN
            exp_f := 82;
        ELSIF x =- 6601 THEN
            exp_f := 82;
        ELSIF x =- 6600 THEN
            exp_f := 82;
        ELSIF x =- 6599 THEN
            exp_f := 82;
        ELSIF x =- 6598 THEN
            exp_f := 82;
        ELSIF x =- 6597 THEN
            exp_f := 82;
        ELSIF x =- 6596 THEN
            exp_f := 82;
        ELSIF x =- 6595 THEN
            exp_f := 82;
        ELSIF x =- 6594 THEN
            exp_f := 82;
        ELSIF x =- 6593 THEN
            exp_f := 82;
        ELSIF x =- 6592 THEN
            exp_f := 82;
        ELSIF x =- 6591 THEN
            exp_f := 82;
        ELSIF x =- 6590 THEN
            exp_f := 82;
        ELSIF x =- 6589 THEN
            exp_f := 82;
        ELSIF x =- 6588 THEN
            exp_f := 82;
        ELSIF x =- 6587 THEN
            exp_f := 82;
        ELSIF x =- 6586 THEN
            exp_f := 82;
        ELSIF x =- 6585 THEN
            exp_f := 82;
        ELSIF x =- 6584 THEN
            exp_f := 82;
        ELSIF x =- 6583 THEN
            exp_f := 82;
        ELSIF x =- 6582 THEN
            exp_f := 83;
        ELSIF x =- 6581 THEN
            exp_f := 83;
        ELSIF x =- 6580 THEN
            exp_f := 83;
        ELSIF x =- 6579 THEN
            exp_f := 83;
        ELSIF x =- 6578 THEN
            exp_f := 83;
        ELSIF x =- 6577 THEN
            exp_f := 83;
        ELSIF x =- 6576 THEN
            exp_f := 83;
        ELSIF x =- 6575 THEN
            exp_f := 83;
        ELSIF x =- 6574 THEN
            exp_f := 83;
        ELSIF x =- 6573 THEN
            exp_f := 83;
        ELSIF x =- 6572 THEN
            exp_f := 83;
        ELSIF x =- 6571 THEN
            exp_f := 83;
        ELSIF x =- 6570 THEN
            exp_f := 83;
        ELSIF x =- 6569 THEN
            exp_f := 83;
        ELSIF x =- 6568 THEN
            exp_f := 83;
        ELSIF x =- 6567 THEN
            exp_f := 83;
        ELSIF x =- 6566 THEN
            exp_f := 83;
        ELSIF x =- 6565 THEN
            exp_f := 83;
        ELSIF x =- 6564 THEN
            exp_f := 83;
        ELSIF x =- 6563 THEN
            exp_f := 83;
        ELSIF x =- 6562 THEN
            exp_f := 83;
        ELSIF x =- 6561 THEN
            exp_f := 83;
        ELSIF x =- 6560 THEN
            exp_f := 83;
        ELSIF x =- 6559 THEN
            exp_f := 83;
        ELSIF x =- 6558 THEN
            exp_f := 84;
        ELSIF x =- 6557 THEN
            exp_f := 84;
        ELSIF x =- 6556 THEN
            exp_f := 84;
        ELSIF x =- 6555 THEN
            exp_f := 84;
        ELSIF x =- 6554 THEN
            exp_f := 84;
        ELSIF x =- 6553 THEN
            exp_f := 84;
        ELSIF x =- 6552 THEN
            exp_f := 84;
        ELSIF x =- 6551 THEN
            exp_f := 84;
        ELSIF x =- 6550 THEN
            exp_f := 84;
        ELSIF x =- 6549 THEN
            exp_f := 84;
        ELSIF x =- 6548 THEN
            exp_f := 84;
        ELSIF x =- 6547 THEN
            exp_f := 84;
        ELSIF x =- 6546 THEN
            exp_f := 84;
        ELSIF x =- 6545 THEN
            exp_f := 84;
        ELSIF x =- 6544 THEN
            exp_f := 84;
        ELSIF x =- 6543 THEN
            exp_f := 84;
        ELSIF x =- 6542 THEN
            exp_f := 84;
        ELSIF x =- 6541 THEN
            exp_f := 84;
        ELSIF x =- 6540 THEN
            exp_f := 84;
        ELSIF x =- 6539 THEN
            exp_f := 84;
        ELSIF x =- 6538 THEN
            exp_f := 84;
        ELSIF x =- 6537 THEN
            exp_f := 84;
        ELSIF x =- 6536 THEN
            exp_f := 84;
        ELSIF x =- 6535 THEN
            exp_f := 84;
        ELSIF x =- 6534 THEN
            exp_f := 85;
        ELSIF x =- 6533 THEN
            exp_f := 85;
        ELSIF x =- 6532 THEN
            exp_f := 85;
        ELSIF x =- 6531 THEN
            exp_f := 85;
        ELSIF x =- 6530 THEN
            exp_f := 85;
        ELSIF x =- 6529 THEN
            exp_f := 85;
        ELSIF x =- 6528 THEN
            exp_f := 85;
        ELSIF x =- 6527 THEN
            exp_f := 85;
        ELSIF x =- 6526 THEN
            exp_f := 85;
        ELSIF x =- 6525 THEN
            exp_f := 85;
        ELSIF x =- 6524 THEN
            exp_f := 85;
        ELSIF x =- 6523 THEN
            exp_f := 85;
        ELSIF x =- 6522 THEN
            exp_f := 85;
        ELSIF x =- 6521 THEN
            exp_f := 85;
        ELSIF x =- 6520 THEN
            exp_f := 85;
        ELSIF x =- 6519 THEN
            exp_f := 85;
        ELSIF x =- 6518 THEN
            exp_f := 85;
        ELSIF x =- 6517 THEN
            exp_f := 85;
        ELSIF x =- 6516 THEN
            exp_f := 85;
        ELSIF x =- 6515 THEN
            exp_f := 85;
        ELSIF x =- 6514 THEN
            exp_f := 85;
        ELSIF x =- 6513 THEN
            exp_f := 85;
        ELSIF x =- 6512 THEN
            exp_f := 85;
        ELSIF x =- 6511 THEN
            exp_f := 85;
        ELSIF x =- 6510 THEN
            exp_f := 85;
        ELSIF x =- 6509 THEN
            exp_f := 86;
        ELSIF x =- 6508 THEN
            exp_f := 86;
        ELSIF x =- 6507 THEN
            exp_f := 86;
        ELSIF x =- 6506 THEN
            exp_f := 86;
        ELSIF x =- 6505 THEN
            exp_f := 86;
        ELSIF x =- 6504 THEN
            exp_f := 86;
        ELSIF x =- 6503 THEN
            exp_f := 86;
        ELSIF x =- 6502 THEN
            exp_f := 86;
        ELSIF x =- 6501 THEN
            exp_f := 86;
        ELSIF x =- 6500 THEN
            exp_f := 86;
        ELSIF x =- 6499 THEN
            exp_f := 86;
        ELSIF x =- 6498 THEN
            exp_f := 86;
        ELSIF x =- 6497 THEN
            exp_f := 86;
        ELSIF x =- 6496 THEN
            exp_f := 86;
        ELSIF x =- 6495 THEN
            exp_f := 86;
        ELSIF x =- 6494 THEN
            exp_f := 86;
        ELSIF x =- 6493 THEN
            exp_f := 86;
        ELSIF x =- 6492 THEN
            exp_f := 86;
        ELSIF x =- 6491 THEN
            exp_f := 86;
        ELSIF x =- 6490 THEN
            exp_f := 86;
        ELSIF x =- 6489 THEN
            exp_f := 86;
        ELSIF x =- 6488 THEN
            exp_f := 86;
        ELSIF x =- 6487 THEN
            exp_f := 86;
        ELSIF x =- 6486 THEN
            exp_f := 86;
        ELSIF x =- 6485 THEN
            exp_f := 87;
        ELSIF x =- 6484 THEN
            exp_f := 87;
        ELSIF x =- 6483 THEN
            exp_f := 87;
        ELSIF x =- 6482 THEN
            exp_f := 87;
        ELSIF x =- 6481 THEN
            exp_f := 87;
        ELSIF x =- 6480 THEN
            exp_f := 87;
        ELSIF x =- 6479 THEN
            exp_f := 87;
        ELSIF x =- 6478 THEN
            exp_f := 87;
        ELSIF x =- 6477 THEN
            exp_f := 87;
        ELSIF x =- 6476 THEN
            exp_f := 87;
        ELSIF x =- 6475 THEN
            exp_f := 87;
        ELSIF x =- 6474 THEN
            exp_f := 87;
        ELSIF x =- 6473 THEN
            exp_f := 87;
        ELSIF x =- 6472 THEN
            exp_f := 87;
        ELSIF x =- 6471 THEN
            exp_f := 87;
        ELSIF x =- 6470 THEN
            exp_f := 87;
        ELSIF x =- 6469 THEN
            exp_f := 87;
        ELSIF x =- 6468 THEN
            exp_f := 87;
        ELSIF x =- 6467 THEN
            exp_f := 87;
        ELSIF x =- 6466 THEN
            exp_f := 87;
        ELSIF x =- 6465 THEN
            exp_f := 87;
        ELSIF x =- 6464 THEN
            exp_f := 87;
        ELSIF x =- 6463 THEN
            exp_f := 87;
        ELSIF x =- 6462 THEN
            exp_f := 87;
        ELSIF x =- 6461 THEN
            exp_f := 87;
        ELSIF x =- 6460 THEN
            exp_f := 88;
        ELSIF x =- 6459 THEN
            exp_f := 88;
        ELSIF x =- 6458 THEN
            exp_f := 88;
        ELSIF x =- 6457 THEN
            exp_f := 88;
        ELSIF x =- 6456 THEN
            exp_f := 88;
        ELSIF x =- 6455 THEN
            exp_f := 88;
        ELSIF x =- 6454 THEN
            exp_f := 88;
        ELSIF x =- 6453 THEN
            exp_f := 88;
        ELSIF x =- 6452 THEN
            exp_f := 88;
        ELSIF x =- 6451 THEN
            exp_f := 88;
        ELSIF x =- 6450 THEN
            exp_f := 88;
        ELSIF x =- 6449 THEN
            exp_f := 88;
        ELSIF x =- 6448 THEN
            exp_f := 88;
        ELSIF x =- 6447 THEN
            exp_f := 88;
        ELSIF x =- 6446 THEN
            exp_f := 88;
        ELSIF x =- 6445 THEN
            exp_f := 88;
        ELSIF x =- 6444 THEN
            exp_f := 88;
        ELSIF x =- 6443 THEN
            exp_f := 88;
        ELSIF x =- 6442 THEN
            exp_f := 88;
        ELSIF x =- 6441 THEN
            exp_f := 88;
        ELSIF x =- 6440 THEN
            exp_f := 88;
        ELSIF x =- 6439 THEN
            exp_f := 88;
        ELSIF x =- 6438 THEN
            exp_f := 88;
        ELSIF x =- 6437 THEN
            exp_f := 88;
        ELSIF x =- 6436 THEN
            exp_f := 89;
        ELSIF x =- 6435 THEN
            exp_f := 89;
        ELSIF x =- 6434 THEN
            exp_f := 89;
        ELSIF x =- 6433 THEN
            exp_f := 89;
        ELSIF x =- 6432 THEN
            exp_f := 89;
        ELSIF x =- 6431 THEN
            exp_f := 89;
        ELSIF x =- 6430 THEN
            exp_f := 89;
        ELSIF x =- 6429 THEN
            exp_f := 89;
        ELSIF x =- 6428 THEN
            exp_f := 89;
        ELSIF x =- 6427 THEN
            exp_f := 89;
        ELSIF x =- 6426 THEN
            exp_f := 89;
        ELSIF x =- 6425 THEN
            exp_f := 89;
        ELSIF x =- 6424 THEN
            exp_f := 89;
        ELSIF x =- 6423 THEN
            exp_f := 89;
        ELSIF x =- 6422 THEN
            exp_f := 89;
        ELSIF x =- 6421 THEN
            exp_f := 89;
        ELSIF x =- 6420 THEN
            exp_f := 89;
        ELSIF x =- 6419 THEN
            exp_f := 89;
        ELSIF x =- 6418 THEN
            exp_f := 89;
        ELSIF x =- 6417 THEN
            exp_f := 89;
        ELSIF x =- 6416 THEN
            exp_f := 89;
        ELSIF x =- 6415 THEN
            exp_f := 89;
        ELSIF x =- 6414 THEN
            exp_f := 89;
        ELSIF x =- 6413 THEN
            exp_f := 89;
        ELSIF x =- 6412 THEN
            exp_f := 90;
        ELSIF x =- 6411 THEN
            exp_f := 90;
        ELSIF x =- 6410 THEN
            exp_f := 90;
        ELSIF x =- 6409 THEN
            exp_f := 90;
        ELSIF x =- 6408 THEN
            exp_f := 90;
        ELSIF x =- 6407 THEN
            exp_f := 90;
        ELSIF x =- 6406 THEN
            exp_f := 90;
        ELSIF x =- 6405 THEN
            exp_f := 90;
        ELSIF x =- 6404 THEN
            exp_f := 90;
        ELSIF x =- 6403 THEN
            exp_f := 90;
        ELSIF x =- 6402 THEN
            exp_f := 90;
        ELSIF x =- 6401 THEN
            exp_f := 90;
        ELSIF x =- 6400 THEN
            exp_f := 90;
        ELSIF x =- 6399 THEN
            exp_f := 90;
        ELSIF x =- 6398 THEN
            exp_f := 90;
        ELSIF x =- 6397 THEN
            exp_f := 90;
        ELSIF x =- 6396 THEN
            exp_f := 90;
        ELSIF x =- 6395 THEN
            exp_f := 90;
        ELSIF x =- 6394 THEN
            exp_f := 90;
        ELSIF x =- 6393 THEN
            exp_f := 90;
        ELSIF x =- 6392 THEN
            exp_f := 90;
        ELSIF x =- 6391 THEN
            exp_f := 90;
        ELSIF x =- 6390 THEN
            exp_f := 90;
        ELSIF x =- 6389 THEN
            exp_f := 90;
        ELSIF x =- 6388 THEN
            exp_f := 90;
        ELSIF x =- 6387 THEN
            exp_f := 91;
        ELSIF x =- 6386 THEN
            exp_f := 91;
        ELSIF x =- 6385 THEN
            exp_f := 91;
        ELSIF x =- 6384 THEN
            exp_f := 91;
        ELSIF x =- 6383 THEN
            exp_f := 91;
        ELSIF x =- 6382 THEN
            exp_f := 91;
        ELSIF x =- 6381 THEN
            exp_f := 91;
        ELSIF x =- 6380 THEN
            exp_f := 91;
        ELSIF x =- 6379 THEN
            exp_f := 91;
        ELSIF x =- 6378 THEN
            exp_f := 91;
        ELSIF x =- 6377 THEN
            exp_f := 91;
        ELSIF x =- 6376 THEN
            exp_f := 91;
        ELSIF x =- 6375 THEN
            exp_f := 91;
        ELSIF x =- 6374 THEN
            exp_f := 91;
        ELSIF x =- 6373 THEN
            exp_f := 91;
        ELSIF x =- 6372 THEN
            exp_f := 91;
        ELSIF x =- 6371 THEN
            exp_f := 91;
        ELSIF x =- 6370 THEN
            exp_f := 91;
        ELSIF x =- 6369 THEN
            exp_f := 91;
        ELSIF x =- 6368 THEN
            exp_f := 91;
        ELSIF x =- 6367 THEN
            exp_f := 91;
        ELSIF x =- 6366 THEN
            exp_f := 91;
        ELSIF x =- 6365 THEN
            exp_f := 91;
        ELSIF x =- 6364 THEN
            exp_f := 91;
        ELSIF x =- 6363 THEN
            exp_f := 93;
        ELSIF x =- 6362 THEN
            exp_f := 93;
        ELSIF x =- 6361 THEN
            exp_f := 93;
        ELSIF x =- 6360 THEN
            exp_f := 93;
        ELSIF x =- 6359 THEN
            exp_f := 93;
        ELSIF x =- 6358 THEN
            exp_f := 93;
        ELSIF x =- 6357 THEN
            exp_f := 93;
        ELSIF x =- 6356 THEN
            exp_f := 93;
        ELSIF x =- 6355 THEN
            exp_f := 93;
        ELSIF x =- 6354 THEN
            exp_f := 93;
        ELSIF x =- 6353 THEN
            exp_f := 93;
        ELSIF x =- 6352 THEN
            exp_f := 93;
        ELSIF x =- 6351 THEN
            exp_f := 93;
        ELSIF x =- 6350 THEN
            exp_f := 93;
        ELSIF x =- 6349 THEN
            exp_f := 93;
        ELSIF x =- 6348 THEN
            exp_f := 93;
        ELSIF x =- 6347 THEN
            exp_f := 93;
        ELSIF x =- 6346 THEN
            exp_f := 93;
        ELSIF x =- 6345 THEN
            exp_f := 93;
        ELSIF x =- 6344 THEN
            exp_f := 93;
        ELSIF x =- 6343 THEN
            exp_f := 93;
        ELSIF x =- 6342 THEN
            exp_f := 93;
        ELSIF x =- 6341 THEN
            exp_f := 93;
        ELSIF x =- 6340 THEN
            exp_f := 93;
        ELSIF x =- 6339 THEN
            exp_f := 94;
        ELSIF x =- 6338 THEN
            exp_f := 94;
        ELSIF x =- 6337 THEN
            exp_f := 94;
        ELSIF x =- 6336 THEN
            exp_f := 94;
        ELSIF x =- 6335 THEN
            exp_f := 94;
        ELSIF x =- 6334 THEN
            exp_f := 94;
        ELSIF x =- 6333 THEN
            exp_f := 94;
        ELSIF x =- 6332 THEN
            exp_f := 94;
        ELSIF x =- 6331 THEN
            exp_f := 94;
        ELSIF x =- 6330 THEN
            exp_f := 94;
        ELSIF x =- 6329 THEN
            exp_f := 94;
        ELSIF x =- 6328 THEN
            exp_f := 94;
        ELSIF x =- 6327 THEN
            exp_f := 94;
        ELSIF x =- 6326 THEN
            exp_f := 94;
        ELSIF x =- 6325 THEN
            exp_f := 94;
        ELSIF x =- 6324 THEN
            exp_f := 94;
        ELSIF x =- 6323 THEN
            exp_f := 94;
        ELSIF x =- 6322 THEN
            exp_f := 94;
        ELSIF x =- 6321 THEN
            exp_f := 94;
        ELSIF x =- 6320 THEN
            exp_f := 94;
        ELSIF x =- 6319 THEN
            exp_f := 94;
        ELSIF x =- 6318 THEN
            exp_f := 94;
        ELSIF x =- 6317 THEN
            exp_f := 94;
        ELSIF x =- 6316 THEN
            exp_f := 94;
        ELSIF x =- 6315 THEN
            exp_f := 94;
        ELSIF x =- 6314 THEN
            exp_f := 95;
        ELSIF x =- 6313 THEN
            exp_f := 95;
        ELSIF x =- 6312 THEN
            exp_f := 95;
        ELSIF x =- 6311 THEN
            exp_f := 95;
        ELSIF x =- 6310 THEN
            exp_f := 95;
        ELSIF x =- 6309 THEN
            exp_f := 95;
        ELSIF x =- 6308 THEN
            exp_f := 95;
        ELSIF x =- 6307 THEN
            exp_f := 95;
        ELSIF x =- 6306 THEN
            exp_f := 95;
        ELSIF x =- 6305 THEN
            exp_f := 95;
        ELSIF x =- 6304 THEN
            exp_f := 95;
        ELSIF x =- 6303 THEN
            exp_f := 95;
        ELSIF x =- 6302 THEN
            exp_f := 95;
        ELSIF x =- 6301 THEN
            exp_f := 95;
        ELSIF x =- 6300 THEN
            exp_f := 95;
        ELSIF x =- 6299 THEN
            exp_f := 95;
        ELSIF x =- 6298 THEN
            exp_f := 95;
        ELSIF x =- 6297 THEN
            exp_f := 95;
        ELSIF x =- 6296 THEN
            exp_f := 95;
        ELSIF x =- 6295 THEN
            exp_f := 95;
        ELSIF x =- 6294 THEN
            exp_f := 95;
        ELSIF x =- 6293 THEN
            exp_f := 95;
        ELSIF x =- 6292 THEN
            exp_f := 95;
        ELSIF x =- 6291 THEN
            exp_f := 95;
        ELSIF x =- 6290 THEN
            exp_f := 96;
        ELSIF x =- 6289 THEN
            exp_f := 96;
        ELSIF x =- 6288 THEN
            exp_f := 96;
        ELSIF x =- 6287 THEN
            exp_f := 96;
        ELSIF x =- 6286 THEN
            exp_f := 96;
        ELSIF x =- 6285 THEN
            exp_f := 96;
        ELSIF x =- 6284 THEN
            exp_f := 96;
        ELSIF x =- 6283 THEN
            exp_f := 96;
        ELSIF x =- 6282 THEN
            exp_f := 96;
        ELSIF x =- 6281 THEN
            exp_f := 96;
        ELSIF x =- 6280 THEN
            exp_f := 96;
        ELSIF x =- 6279 THEN
            exp_f := 96;
        ELSIF x =- 6278 THEN
            exp_f := 96;
        ELSIF x =- 6277 THEN
            exp_f := 96;
        ELSIF x =- 6276 THEN
            exp_f := 96;
        ELSIF x =- 6275 THEN
            exp_f := 96;
        ELSIF x =- 6274 THEN
            exp_f := 96;
        ELSIF x =- 6273 THEN
            exp_f := 96;
        ELSIF x =- 6272 THEN
            exp_f := 96;
        ELSIF x =- 6271 THEN
            exp_f := 96;
        ELSIF x =- 6270 THEN
            exp_f := 96;
        ELSIF x =- 6269 THEN
            exp_f := 96;
        ELSIF x =- 6268 THEN
            exp_f := 96;
        ELSIF x =- 6267 THEN
            exp_f := 96;
        ELSIF x =- 6266 THEN
            exp_f := 96;
        ELSIF x =- 6265 THEN
            exp_f := 97;
        ELSIF x =- 6264 THEN
            exp_f := 97;
        ELSIF x =- 6263 THEN
            exp_f := 97;
        ELSIF x =- 6262 THEN
            exp_f := 97;
        ELSIF x =- 6261 THEN
            exp_f := 97;
        ELSIF x =- 6260 THEN
            exp_f := 97;
        ELSIF x =- 6259 THEN
            exp_f := 97;
        ELSIF x =- 6258 THEN
            exp_f := 97;
        ELSIF x =- 6257 THEN
            exp_f := 97;
        ELSIF x =- 6256 THEN
            exp_f := 97;
        ELSIF x =- 6255 THEN
            exp_f := 97;
        ELSIF x =- 6254 THEN
            exp_f := 97;
        ELSIF x =- 6253 THEN
            exp_f := 97;
        ELSIF x =- 6252 THEN
            exp_f := 97;
        ELSIF x =- 6251 THEN
            exp_f := 97;
        ELSIF x =- 6250 THEN
            exp_f := 97;
        ELSIF x =- 6249 THEN
            exp_f := 97;
        ELSIF x =- 6248 THEN
            exp_f := 97;
        ELSIF x =- 6247 THEN
            exp_f := 97;
        ELSIF x =- 6246 THEN
            exp_f := 97;
        ELSIF x =- 6245 THEN
            exp_f := 97;
        ELSIF x =- 6244 THEN
            exp_f := 97;
        ELSIF x =- 6243 THEN
            exp_f := 97;
        ELSIF x =- 6242 THEN
            exp_f := 97;
        ELSIF x =- 6241 THEN
            exp_f := 98;
        ELSIF x =- 6240 THEN
            exp_f := 98;
        ELSIF x =- 6239 THEN
            exp_f := 98;
        ELSIF x =- 6238 THEN
            exp_f := 98;
        ELSIF x =- 6237 THEN
            exp_f := 98;
        ELSIF x =- 6236 THEN
            exp_f := 98;
        ELSIF x =- 6235 THEN
            exp_f := 98;
        ELSIF x =- 6234 THEN
            exp_f := 98;
        ELSIF x =- 6233 THEN
            exp_f := 98;
        ELSIF x =- 6232 THEN
            exp_f := 98;
        ELSIF x =- 6231 THEN
            exp_f := 98;
        ELSIF x =- 6230 THEN
            exp_f := 98;
        ELSIF x =- 6229 THEN
            exp_f := 98;
        ELSIF x =- 6228 THEN
            exp_f := 98;
        ELSIF x =- 6227 THEN
            exp_f := 98;
        ELSIF x =- 6226 THEN
            exp_f := 98;
        ELSIF x =- 6225 THEN
            exp_f := 98;
        ELSIF x =- 6224 THEN
            exp_f := 98;
        ELSIF x =- 6223 THEN
            exp_f := 98;
        ELSIF x =- 6222 THEN
            exp_f := 98;
        ELSIF x =- 6221 THEN
            exp_f := 98;
        ELSIF x =- 6220 THEN
            exp_f := 98;
        ELSIF x =- 6219 THEN
            exp_f := 98;
        ELSIF x =- 6218 THEN
            exp_f := 98;
        ELSIF x =- 6217 THEN
            exp_f := 99;
        ELSIF x =- 6216 THEN
            exp_f := 99;
        ELSIF x =- 6215 THEN
            exp_f := 99;
        ELSIF x =- 6214 THEN
            exp_f := 99;
        ELSIF x =- 6213 THEN
            exp_f := 99;
        ELSIF x =- 6212 THEN
            exp_f := 99;
        ELSIF x =- 6211 THEN
            exp_f := 99;
        ELSIF x =- 6210 THEN
            exp_f := 99;
        ELSIF x =- 6209 THEN
            exp_f := 99;
        ELSIF x =- 6208 THEN
            exp_f := 99;
        ELSIF x =- 6207 THEN
            exp_f := 99;
        ELSIF x =- 6206 THEN
            exp_f := 99;
        ELSIF x =- 6205 THEN
            exp_f := 99;
        ELSIF x =- 6204 THEN
            exp_f := 99;
        ELSIF x =- 6203 THEN
            exp_f := 99;
        ELSIF x =- 6202 THEN
            exp_f := 99;
        ELSIF x =- 6201 THEN
            exp_f := 99;
        ELSIF x =- 6200 THEN
            exp_f := 99;
        ELSIF x =- 6199 THEN
            exp_f := 99;
        ELSIF x =- 6198 THEN
            exp_f := 99;
        ELSIF x =- 6197 THEN
            exp_f := 99;
        ELSIF x =- 6196 THEN
            exp_f := 99;
        ELSIF x =- 6195 THEN
            exp_f := 99;
        ELSIF x =- 6194 THEN
            exp_f := 99;
        ELSIF x =- 6193 THEN
            exp_f := 99;
        ELSIF x =- 6192 THEN
            exp_f := 100;
        ELSIF x =- 6191 THEN
            exp_f := 100;
        ELSIF x =- 6190 THEN
            exp_f := 100;
        ELSIF x =- 6189 THEN
            exp_f := 100;
        ELSIF x =- 6188 THEN
            exp_f := 100;
        ELSIF x =- 6187 THEN
            exp_f := 100;
        ELSIF x =- 6186 THEN
            exp_f := 100;
        ELSIF x =- 6185 THEN
            exp_f := 100;
        ELSIF x =- 6184 THEN
            exp_f := 100;
        ELSIF x =- 6183 THEN
            exp_f := 100;
        ELSIF x =- 6182 THEN
            exp_f := 100;
        ELSIF x =- 6181 THEN
            exp_f := 100;
        ELSIF x =- 6180 THEN
            exp_f := 100;
        ELSIF x =- 6179 THEN
            exp_f := 100;
        ELSIF x =- 6178 THEN
            exp_f := 100;
        ELSIF x =- 6177 THEN
            exp_f := 100;
        ELSIF x =- 6176 THEN
            exp_f := 100;
        ELSIF x =- 6175 THEN
            exp_f := 100;
        ELSIF x =- 6174 THEN
            exp_f := 100;
        ELSIF x =- 6173 THEN
            exp_f := 100;
        ELSIF x =- 6172 THEN
            exp_f := 100;
        ELSIF x =- 6171 THEN
            exp_f := 100;
        ELSIF x =- 6170 THEN
            exp_f := 100;
        ELSIF x =- 6169 THEN
            exp_f := 100;
        ELSIF x =- 6168 THEN
            exp_f := 101;
        ELSIF x =- 6167 THEN
            exp_f := 101;
        ELSIF x =- 6166 THEN
            exp_f := 101;
        ELSIF x =- 6165 THEN
            exp_f := 101;
        ELSIF x =- 6164 THEN
            exp_f := 101;
        ELSIF x =- 6163 THEN
            exp_f := 101;
        ELSIF x =- 6162 THEN
            exp_f := 101;
        ELSIF x =- 6161 THEN
            exp_f := 101;
        ELSIF x =- 6160 THEN
            exp_f := 101;
        ELSIF x =- 6159 THEN
            exp_f := 101;
        ELSIF x =- 6158 THEN
            exp_f := 101;
        ELSIF x =- 6157 THEN
            exp_f := 101;
        ELSIF x =- 6156 THEN
            exp_f := 101;
        ELSIF x =- 6155 THEN
            exp_f := 101;
        ELSIF x =- 6154 THEN
            exp_f := 101;
        ELSIF x =- 6153 THEN
            exp_f := 101;
        ELSIF x =- 6152 THEN
            exp_f := 101;
        ELSIF x =- 6151 THEN
            exp_f := 101;
        ELSIF x =- 6150 THEN
            exp_f := 101;
        ELSIF x =- 6149 THEN
            exp_f := 101;
        ELSIF x =- 6148 THEN
            exp_f := 101;
        ELSIF x =- 6147 THEN
            exp_f := 101;
        ELSIF x =- 6146 THEN
            exp_f := 101;
        ELSIF x =- 6145 THEN
            exp_f := 101;
        ELSIF x =- 6144 THEN
            exp_f := 101;
        ELSIF x =- 6143 THEN
            exp_f := 102;
        ELSIF x =- 6142 THEN
            exp_f := 102;
        ELSIF x =- 6141 THEN
            exp_f := 102;
        ELSIF x =- 6140 THEN
            exp_f := 102;
        ELSIF x =- 6139 THEN
            exp_f := 102;
        ELSIF x =- 6138 THEN
            exp_f := 102;
        ELSIF x =- 6137 THEN
            exp_f := 102;
        ELSIF x =- 6136 THEN
            exp_f := 102;
        ELSIF x =- 6135 THEN
            exp_f := 102;
        ELSIF x =- 6134 THEN
            exp_f := 102;
        ELSIF x =- 6133 THEN
            exp_f := 102;
        ELSIF x =- 6132 THEN
            exp_f := 102;
        ELSIF x =- 6131 THEN
            exp_f := 102;
        ELSIF x =- 6130 THEN
            exp_f := 102;
        ELSIF x =- 6129 THEN
            exp_f := 102;
        ELSIF x =- 6128 THEN
            exp_f := 102;
        ELSIF x =- 6127 THEN
            exp_f := 102;
        ELSIF x =- 6126 THEN
            exp_f := 102;
        ELSIF x =- 6125 THEN
            exp_f := 102;
        ELSIF x =- 6124 THEN
            exp_f := 102;
        ELSIF x =- 6123 THEN
            exp_f := 104;
        ELSIF x =- 6122 THEN
            exp_f := 104;
        ELSIF x =- 6121 THEN
            exp_f := 104;
        ELSIF x =- 6120 THEN
            exp_f := 104;
        ELSIF x =- 6119 THEN
            exp_f := 104;
        ELSIF x =- 6118 THEN
            exp_f := 104;
        ELSIF x =- 6117 THEN
            exp_f := 104;
        ELSIF x =- 6116 THEN
            exp_f := 104;
        ELSIF x =- 6115 THEN
            exp_f := 104;
        ELSIF x =- 6114 THEN
            exp_f := 104;
        ELSIF x =- 6113 THEN
            exp_f := 104;
        ELSIF x =- 6112 THEN
            exp_f := 104;
        ELSIF x =- 6111 THEN
            exp_f := 104;
        ELSIF x =- 6110 THEN
            exp_f := 104;
        ELSIF x =- 6109 THEN
            exp_f := 104;
        ELSIF x =- 6108 THEN
            exp_f := 104;
        ELSIF x =- 6107 THEN
            exp_f := 104;
        ELSIF x =- 6106 THEN
            exp_f := 104;
        ELSIF x =- 6105 THEN
            exp_f := 104;
        ELSIF x =- 6104 THEN
            exp_f := 104;
        ELSIF x =- 6103 THEN
            exp_f := 105;
        ELSIF x =- 6102 THEN
            exp_f := 105;
        ELSIF x =- 6101 THEN
            exp_f := 105;
        ELSIF x =- 6100 THEN
            exp_f := 105;
        ELSIF x =- 6099 THEN
            exp_f := 105;
        ELSIF x =- 6098 THEN
            exp_f := 105;
        ELSIF x =- 6097 THEN
            exp_f := 105;
        ELSIF x =- 6096 THEN
            exp_f := 105;
        ELSIF x =- 6095 THEN
            exp_f := 105;
        ELSIF x =- 6094 THEN
            exp_f := 105;
        ELSIF x =- 6093 THEN
            exp_f := 105;
        ELSIF x =- 6092 THEN
            exp_f := 105;
        ELSIF x =- 6091 THEN
            exp_f := 105;
        ELSIF x =- 6090 THEN
            exp_f := 105;
        ELSIF x =- 6089 THEN
            exp_f := 105;
        ELSIF x =- 6088 THEN
            exp_f := 105;
        ELSIF x =- 6087 THEN
            exp_f := 105;
        ELSIF x =- 6086 THEN
            exp_f := 105;
        ELSIF x =- 6085 THEN
            exp_f := 105;
        ELSIF x =- 6084 THEN
            exp_f := 105;
        ELSIF x =- 6083 THEN
            exp_f := 106;
        ELSIF x =- 6082 THEN
            exp_f := 106;
        ELSIF x =- 6081 THEN
            exp_f := 106;
        ELSIF x =- 6080 THEN
            exp_f := 106;
        ELSIF x =- 6079 THEN
            exp_f := 106;
        ELSIF x =- 6078 THEN
            exp_f := 106;
        ELSIF x =- 6077 THEN
            exp_f := 106;
        ELSIF x =- 6076 THEN
            exp_f := 106;
        ELSIF x =- 6075 THEN
            exp_f := 106;
        ELSIF x =- 6074 THEN
            exp_f := 106;
        ELSIF x =- 6073 THEN
            exp_f := 106;
        ELSIF x =- 6072 THEN
            exp_f := 106;
        ELSIF x =- 6071 THEN
            exp_f := 106;
        ELSIF x =- 6070 THEN
            exp_f := 106;
        ELSIF x =- 6069 THEN
            exp_f := 106;
        ELSIF x =- 6068 THEN
            exp_f := 106;
        ELSIF x =- 6067 THEN
            exp_f := 106;
        ELSIF x =- 6066 THEN
            exp_f := 106;
        ELSIF x =- 6065 THEN
            exp_f := 106;
        ELSIF x =- 6064 THEN
            exp_f := 106;
        ELSIF x =- 6063 THEN
            exp_f := 107;
        ELSIF x =- 6062 THEN
            exp_f := 107;
        ELSIF x =- 6061 THEN
            exp_f := 107;
        ELSIF x =- 6060 THEN
            exp_f := 107;
        ELSIF x =- 6059 THEN
            exp_f := 107;
        ELSIF x =- 6058 THEN
            exp_f := 107;
        ELSIF x =- 6057 THEN
            exp_f := 107;
        ELSIF x =- 6056 THEN
            exp_f := 107;
        ELSIF x =- 6055 THEN
            exp_f := 107;
        ELSIF x =- 6054 THEN
            exp_f := 107;
        ELSIF x =- 6053 THEN
            exp_f := 107;
        ELSIF x =- 6052 THEN
            exp_f := 107;
        ELSIF x =- 6051 THEN
            exp_f := 107;
        ELSIF x =- 6050 THEN
            exp_f := 107;
        ELSIF x =- 6049 THEN
            exp_f := 107;
        ELSIF x =- 6048 THEN
            exp_f := 107;
        ELSIF x =- 6047 THEN
            exp_f := 107;
        ELSIF x =- 6046 THEN
            exp_f := 107;
        ELSIF x =- 6045 THEN
            exp_f := 107;
        ELSIF x =- 6044 THEN
            exp_f := 107;
        ELSIF x =- 6043 THEN
            exp_f := 108;
        ELSIF x =- 6042 THEN
            exp_f := 108;
        ELSIF x =- 6041 THEN
            exp_f := 108;
        ELSIF x =- 6040 THEN
            exp_f := 108;
        ELSIF x =- 6039 THEN
            exp_f := 108;
        ELSIF x =- 6038 THEN
            exp_f := 108;
        ELSIF x =- 6037 THEN
            exp_f := 108;
        ELSIF x =- 6036 THEN
            exp_f := 108;
        ELSIF x =- 6035 THEN
            exp_f := 108;
        ELSIF x =- 6034 THEN
            exp_f := 108;
        ELSIF x =- 6033 THEN
            exp_f := 108;
        ELSIF x =- 6032 THEN
            exp_f := 108;
        ELSIF x =- 6031 THEN
            exp_f := 108;
        ELSIF x =- 6030 THEN
            exp_f := 108;
        ELSIF x =- 6029 THEN
            exp_f := 108;
        ELSIF x =- 6028 THEN
            exp_f := 108;
        ELSIF x =- 6027 THEN
            exp_f := 108;
        ELSIF x =- 6026 THEN
            exp_f := 108;
        ELSIF x =- 6025 THEN
            exp_f := 108;
        ELSIF x =- 6024 THEN
            exp_f := 108;
        ELSIF x =- 6023 THEN
            exp_f := 109;
        ELSIF x =- 6022 THEN
            exp_f := 109;
        ELSIF x =- 6021 THEN
            exp_f := 109;
        ELSIF x =- 6020 THEN
            exp_f := 109;
        ELSIF x =- 6019 THEN
            exp_f := 109;
        ELSIF x =- 6018 THEN
            exp_f := 109;
        ELSIF x =- 6017 THEN
            exp_f := 109;
        ELSIF x =- 6016 THEN
            exp_f := 109;
        ELSIF x =- 6015 THEN
            exp_f := 109;
        ELSIF x =- 6014 THEN
            exp_f := 109;
        ELSIF x =- 6013 THEN
            exp_f := 109;
        ELSIF x =- 6012 THEN
            exp_f := 109;
        ELSIF x =- 6011 THEN
            exp_f := 109;
        ELSIF x =- 6010 THEN
            exp_f := 109;
        ELSIF x =- 6009 THEN
            exp_f := 109;
        ELSIF x =- 6008 THEN
            exp_f := 109;
        ELSIF x =- 6007 THEN
            exp_f := 109;
        ELSIF x =- 6006 THEN
            exp_f := 109;
        ELSIF x =- 6005 THEN
            exp_f := 109;
        ELSIF x =- 6004 THEN
            exp_f := 109;
        ELSIF x =- 6003 THEN
            exp_f := 110;
        ELSIF x =- 6002 THEN
            exp_f := 110;
        ELSIF x =- 6001 THEN
            exp_f := 110;
        ELSIF x =- 6000 THEN
            exp_f := 110;
        ELSIF x =- 5999 THEN
            exp_f := 110;
        ELSIF x =- 5998 THEN
            exp_f := 110;
        ELSIF x =- 5997 THEN
            exp_f := 110;
        ELSIF x =- 5996 THEN
            exp_f := 110;
        ELSIF x =- 5995 THEN
            exp_f := 110;
        ELSIF x =- 5994 THEN
            exp_f := 110;
        ELSIF x =- 5993 THEN
            exp_f := 110;
        ELSIF x =- 5992 THEN
            exp_f := 110;
        ELSIF x =- 5991 THEN
            exp_f := 110;
        ELSIF x =- 5990 THEN
            exp_f := 110;
        ELSIF x =- 5989 THEN
            exp_f := 110;
        ELSIF x =- 5988 THEN
            exp_f := 110;
        ELSIF x =- 5987 THEN
            exp_f := 110;
        ELSIF x =- 5986 THEN
            exp_f := 110;
        ELSIF x =- 5985 THEN
            exp_f := 110;
        ELSIF x =- 5984 THEN
            exp_f := 110;
        ELSIF x =- 5983 THEN
            exp_f := 111;
        ELSIF x =- 5982 THEN
            exp_f := 111;
        ELSIF x =- 5981 THEN
            exp_f := 111;
        ELSIF x =- 5980 THEN
            exp_f := 111;
        ELSIF x =- 5979 THEN
            exp_f := 111;
        ELSIF x =- 5978 THEN
            exp_f := 111;
        ELSIF x =- 5977 THEN
            exp_f := 111;
        ELSIF x =- 5976 THEN
            exp_f := 111;
        ELSIF x =- 5975 THEN
            exp_f := 111;
        ELSIF x =- 5974 THEN
            exp_f := 111;
        ELSIF x =- 5973 THEN
            exp_f := 111;
        ELSIF x =- 5972 THEN
            exp_f := 111;
        ELSIF x =- 5971 THEN
            exp_f := 111;
        ELSIF x =- 5970 THEN
            exp_f := 111;
        ELSIF x =- 5969 THEN
            exp_f := 111;
        ELSIF x =- 5968 THEN
            exp_f := 111;
        ELSIF x =- 5967 THEN
            exp_f := 111;
        ELSIF x =- 5966 THEN
            exp_f := 111;
        ELSIF x =- 5965 THEN
            exp_f := 111;
        ELSIF x =- 5964 THEN
            exp_f := 111;
        ELSIF x =- 5963 THEN
            exp_f := 112;
        ELSIF x =- 5962 THEN
            exp_f := 112;
        ELSIF x =- 5961 THEN
            exp_f := 112;
        ELSIF x =- 5960 THEN
            exp_f := 112;
        ELSIF x =- 5959 THEN
            exp_f := 112;
        ELSIF x =- 5958 THEN
            exp_f := 112;
        ELSIF x =- 5957 THEN
            exp_f := 112;
        ELSIF x =- 5956 THEN
            exp_f := 112;
        ELSIF x =- 5955 THEN
            exp_f := 112;
        ELSIF x =- 5954 THEN
            exp_f := 112;
        ELSIF x =- 5953 THEN
            exp_f := 112;
        ELSIF x =- 5952 THEN
            exp_f := 112;
        ELSIF x =- 5951 THEN
            exp_f := 112;
        ELSIF x =- 5950 THEN
            exp_f := 112;
        ELSIF x =- 5949 THEN
            exp_f := 112;
        ELSIF x =- 5948 THEN
            exp_f := 112;
        ELSIF x =- 5947 THEN
            exp_f := 112;
        ELSIF x =- 5946 THEN
            exp_f := 112;
        ELSIF x =- 5945 THEN
            exp_f := 112;
        ELSIF x =- 5944 THEN
            exp_f := 112;
        ELSIF x =- 5943 THEN
            exp_f := 114;
        ELSIF x =- 5942 THEN
            exp_f := 114;
        ELSIF x =- 5941 THEN
            exp_f := 114;
        ELSIF x =- 5940 THEN
            exp_f := 114;
        ELSIF x =- 5939 THEN
            exp_f := 114;
        ELSIF x =- 5938 THEN
            exp_f := 114;
        ELSIF x =- 5937 THEN
            exp_f := 114;
        ELSIF x =- 5936 THEN
            exp_f := 114;
        ELSIF x =- 5935 THEN
            exp_f := 114;
        ELSIF x =- 5934 THEN
            exp_f := 114;
        ELSIF x =- 5933 THEN
            exp_f := 114;
        ELSIF x =- 5932 THEN
            exp_f := 114;
        ELSIF x =- 5931 THEN
            exp_f := 114;
        ELSIF x =- 5930 THEN
            exp_f := 114;
        ELSIF x =- 5929 THEN
            exp_f := 114;
        ELSIF x =- 5928 THEN
            exp_f := 114;
        ELSIF x =- 5927 THEN
            exp_f := 114;
        ELSIF x =- 5926 THEN
            exp_f := 114;
        ELSIF x =- 5925 THEN
            exp_f := 114;
        ELSIF x =- 5924 THEN
            exp_f := 114;
        ELSIF x =- 5923 THEN
            exp_f := 115;
        ELSIF x =- 5922 THEN
            exp_f := 115;
        ELSIF x =- 5921 THEN
            exp_f := 115;
        ELSIF x =- 5920 THEN
            exp_f := 115;
        ELSIF x =- 5919 THEN
            exp_f := 115;
        ELSIF x =- 5918 THEN
            exp_f := 115;
        ELSIF x =- 5917 THEN
            exp_f := 115;
        ELSIF x =- 5916 THEN
            exp_f := 115;
        ELSIF x =- 5915 THEN
            exp_f := 115;
        ELSIF x =- 5914 THEN
            exp_f := 115;
        ELSIF x =- 5913 THEN
            exp_f := 115;
        ELSIF x =- 5912 THEN
            exp_f := 115;
        ELSIF x =- 5911 THEN
            exp_f := 115;
        ELSIF x =- 5910 THEN
            exp_f := 115;
        ELSIF x =- 5909 THEN
            exp_f := 115;
        ELSIF x =- 5908 THEN
            exp_f := 115;
        ELSIF x =- 5907 THEN
            exp_f := 115;
        ELSIF x =- 5906 THEN
            exp_f := 115;
        ELSIF x =- 5905 THEN
            exp_f := 115;
        ELSIF x =- 5904 THEN
            exp_f := 115;
        ELSIF x =- 5903 THEN
            exp_f := 116;
        ELSIF x =- 5902 THEN
            exp_f := 116;
        ELSIF x =- 5901 THEN
            exp_f := 116;
        ELSIF x =- 5900 THEN
            exp_f := 116;
        ELSIF x =- 5899 THEN
            exp_f := 116;
        ELSIF x =- 5898 THEN
            exp_f := 116;
        ELSIF x =- 5897 THEN
            exp_f := 116;
        ELSIF x =- 5896 THEN
            exp_f := 116;
        ELSIF x =- 5895 THEN
            exp_f := 116;
        ELSIF x =- 5894 THEN
            exp_f := 116;
        ELSIF x =- 5893 THEN
            exp_f := 116;
        ELSIF x =- 5892 THEN
            exp_f := 116;
        ELSIF x =- 5891 THEN
            exp_f := 116;
        ELSIF x =- 5890 THEN
            exp_f := 116;
        ELSIF x =- 5889 THEN
            exp_f := 116;
        ELSIF x =- 5888 THEN
            exp_f := 116;
        ELSIF x =- 5887 THEN
            exp_f := 116;
        ELSIF x =- 5886 THEN
            exp_f := 116;
        ELSIF x =- 5885 THEN
            exp_f := 116;
        ELSIF x =- 5884 THEN
            exp_f := 116;
        ELSIF x =- 5883 THEN
            exp_f := 116;
        ELSIF x =- 5882 THEN
            exp_f := 117;
        ELSIF x =- 5881 THEN
            exp_f := 117;
        ELSIF x =- 5880 THEN
            exp_f := 117;
        ELSIF x =- 5879 THEN
            exp_f := 117;
        ELSIF x =- 5878 THEN
            exp_f := 117;
        ELSIF x =- 5877 THEN
            exp_f := 117;
        ELSIF x =- 5876 THEN
            exp_f := 117;
        ELSIF x =- 5875 THEN
            exp_f := 117;
        ELSIF x =- 5874 THEN
            exp_f := 117;
        ELSIF x =- 5873 THEN
            exp_f := 117;
        ELSIF x =- 5872 THEN
            exp_f := 117;
        ELSIF x =- 5871 THEN
            exp_f := 117;
        ELSIF x =- 5870 THEN
            exp_f := 117;
        ELSIF x =- 5869 THEN
            exp_f := 117;
        ELSIF x =- 5868 THEN
            exp_f := 117;
        ELSIF x =- 5867 THEN
            exp_f := 117;
        ELSIF x =- 5866 THEN
            exp_f := 117;
        ELSIF x =- 5865 THEN
            exp_f := 117;
        ELSIF x =- 5864 THEN
            exp_f := 117;
        ELSIF x =- 5863 THEN
            exp_f := 117;
        ELSIF x =- 5862 THEN
            exp_f := 118;
        ELSIF x =- 5861 THEN
            exp_f := 118;
        ELSIF x =- 5860 THEN
            exp_f := 118;
        ELSIF x =- 5859 THEN
            exp_f := 118;
        ELSIF x =- 5858 THEN
            exp_f := 118;
        ELSIF x =- 5857 THEN
            exp_f := 118;
        ELSIF x =- 5856 THEN
            exp_f := 118;
        ELSIF x =- 5855 THEN
            exp_f := 118;
        ELSIF x =- 5854 THEN
            exp_f := 118;
        ELSIF x =- 5853 THEN
            exp_f := 118;
        ELSIF x =- 5852 THEN
            exp_f := 118;
        ELSIF x =- 5851 THEN
            exp_f := 118;
        ELSIF x =- 5850 THEN
            exp_f := 118;
        ELSIF x =- 5849 THEN
            exp_f := 118;
        ELSIF x =- 5848 THEN
            exp_f := 118;
        ELSIF x =- 5847 THEN
            exp_f := 118;
        ELSIF x =- 5846 THEN
            exp_f := 118;
        ELSIF x =- 5845 THEN
            exp_f := 118;
        ELSIF x =- 5844 THEN
            exp_f := 118;
        ELSIF x =- 5843 THEN
            exp_f := 118;
        ELSIF x =- 5842 THEN
            exp_f := 119;
        ELSIF x =- 5841 THEN
            exp_f := 119;
        ELSIF x =- 5840 THEN
            exp_f := 119;
        ELSIF x =- 5839 THEN
            exp_f := 119;
        ELSIF x =- 5838 THEN
            exp_f := 119;
        ELSIF x =- 5837 THEN
            exp_f := 119;
        ELSIF x =- 5836 THEN
            exp_f := 119;
        ELSIF x =- 5835 THEN
            exp_f := 119;
        ELSIF x =- 5834 THEN
            exp_f := 119;
        ELSIF x =- 5833 THEN
            exp_f := 119;
        ELSIF x =- 5832 THEN
            exp_f := 119;
        ELSIF x =- 5831 THEN
            exp_f := 119;
        ELSIF x =- 5830 THEN
            exp_f := 119;
        ELSIF x =- 5829 THEN
            exp_f := 119;
        ELSIF x =- 5828 THEN
            exp_f := 119;
        ELSIF x =- 5827 THEN
            exp_f := 119;
        ELSIF x =- 5826 THEN
            exp_f := 119;
        ELSIF x =- 5825 THEN
            exp_f := 119;
        ELSIF x =- 5824 THEN
            exp_f := 119;
        ELSIF x =- 5823 THEN
            exp_f := 119;
        ELSIF x =- 5822 THEN
            exp_f := 120;
        ELSIF x =- 5821 THEN
            exp_f := 120;
        ELSIF x =- 5820 THEN
            exp_f := 120;
        ELSIF x =- 5819 THEN
            exp_f := 120;
        ELSIF x =- 5818 THEN
            exp_f := 120;
        ELSIF x =- 5817 THEN
            exp_f := 120;
        ELSIF x =- 5816 THEN
            exp_f := 120;
        ELSIF x =- 5815 THEN
            exp_f := 120;
        ELSIF x =- 5814 THEN
            exp_f := 120;
        ELSIF x =- 5813 THEN
            exp_f := 120;
        ELSIF x =- 5812 THEN
            exp_f := 120;
        ELSIF x =- 5811 THEN
            exp_f := 120;
        ELSIF x =- 5810 THEN
            exp_f := 120;
        ELSIF x =- 5809 THEN
            exp_f := 120;
        ELSIF x =- 5808 THEN
            exp_f := 120;
        ELSIF x =- 5807 THEN
            exp_f := 120;
        ELSIF x =- 5806 THEN
            exp_f := 120;
        ELSIF x =- 5805 THEN
            exp_f := 120;
        ELSIF x =- 5804 THEN
            exp_f := 120;
        ELSIF x =- 5803 THEN
            exp_f := 120;
        ELSIF x =- 5802 THEN
            exp_f := 121;
        ELSIF x =- 5801 THEN
            exp_f := 121;
        ELSIF x =- 5800 THEN
            exp_f := 121;
        ELSIF x =- 5799 THEN
            exp_f := 121;
        ELSIF x =- 5798 THEN
            exp_f := 121;
        ELSIF x =- 5797 THEN
            exp_f := 121;
        ELSIF x =- 5796 THEN
            exp_f := 121;
        ELSIF x =- 5795 THEN
            exp_f := 121;
        ELSIF x =- 5794 THEN
            exp_f := 121;
        ELSIF x =- 5793 THEN
            exp_f := 121;
        ELSIF x =- 5792 THEN
            exp_f := 121;
        ELSIF x =- 5791 THEN
            exp_f := 121;
        ELSIF x =- 5790 THEN
            exp_f := 121;
        ELSIF x =- 5789 THEN
            exp_f := 121;
        ELSIF x =- 5788 THEN
            exp_f := 121;
        ELSIF x =- 5787 THEN
            exp_f := 121;
        ELSIF x =- 5786 THEN
            exp_f := 121;
        ELSIF x =- 5785 THEN
            exp_f := 121;
        ELSIF x =- 5784 THEN
            exp_f := 121;
        ELSIF x =- 5783 THEN
            exp_f := 121;
        ELSIF x =- 5782 THEN
            exp_f := 122;
        ELSIF x =- 5781 THEN
            exp_f := 122;
        ELSIF x =- 5780 THEN
            exp_f := 122;
        ELSIF x =- 5779 THEN
            exp_f := 122;
        ELSIF x =- 5778 THEN
            exp_f := 122;
        ELSIF x =- 5777 THEN
            exp_f := 122;
        ELSIF x =- 5776 THEN
            exp_f := 122;
        ELSIF x =- 5775 THEN
            exp_f := 122;
        ELSIF x =- 5774 THEN
            exp_f := 122;
        ELSIF x =- 5773 THEN
            exp_f := 122;
        ELSIF x =- 5772 THEN
            exp_f := 122;
        ELSIF x =- 5771 THEN
            exp_f := 122;
        ELSIF x =- 5770 THEN
            exp_f := 122;
        ELSIF x =- 5769 THEN
            exp_f := 122;
        ELSIF x =- 5768 THEN
            exp_f := 122;
        ELSIF x =- 5767 THEN
            exp_f := 122;
        ELSIF x =- 5766 THEN
            exp_f := 122;
        ELSIF x =- 5765 THEN
            exp_f := 122;
        ELSIF x =- 5764 THEN
            exp_f := 122;
        ELSIF x =- 5763 THEN
            exp_f := 122;
        ELSIF x =- 5762 THEN
            exp_f := 124;
        ELSIF x =- 5761 THEN
            exp_f := 124;
        ELSIF x =- 5760 THEN
            exp_f := 124;
        ELSIF x =- 5759 THEN
            exp_f := 124;
        ELSIF x =- 5758 THEN
            exp_f := 124;
        ELSIF x =- 5757 THEN
            exp_f := 124;
        ELSIF x =- 5756 THEN
            exp_f := 124;
        ELSIF x =- 5755 THEN
            exp_f := 124;
        ELSIF x =- 5754 THEN
            exp_f := 124;
        ELSIF x =- 5753 THEN
            exp_f := 124;
        ELSIF x =- 5752 THEN
            exp_f := 124;
        ELSIF x =- 5751 THEN
            exp_f := 124;
        ELSIF x =- 5750 THEN
            exp_f := 124;
        ELSIF x =- 5749 THEN
            exp_f := 124;
        ELSIF x =- 5748 THEN
            exp_f := 124;
        ELSIF x =- 5747 THEN
            exp_f := 124;
        ELSIF x =- 5746 THEN
            exp_f := 124;
        ELSIF x =- 5745 THEN
            exp_f := 124;
        ELSIF x =- 5744 THEN
            exp_f := 124;
        ELSIF x =- 5743 THEN
            exp_f := 124;
        ELSIF x =- 5742 THEN
            exp_f := 125;
        ELSIF x =- 5741 THEN
            exp_f := 125;
        ELSIF x =- 5740 THEN
            exp_f := 125;
        ELSIF x =- 5739 THEN
            exp_f := 125;
        ELSIF x =- 5738 THEN
            exp_f := 125;
        ELSIF x =- 5737 THEN
            exp_f := 125;
        ELSIF x =- 5736 THEN
            exp_f := 125;
        ELSIF x =- 5735 THEN
            exp_f := 125;
        ELSIF x =- 5734 THEN
            exp_f := 125;
        ELSIF x =- 5733 THEN
            exp_f := 125;
        ELSIF x =- 5732 THEN
            exp_f := 125;
        ELSIF x =- 5731 THEN
            exp_f := 125;
        ELSIF x =- 5730 THEN
            exp_f := 125;
        ELSIF x =- 5729 THEN
            exp_f := 125;
        ELSIF x =- 5728 THEN
            exp_f := 125;
        ELSIF x =- 5727 THEN
            exp_f := 125;
        ELSIF x =- 5726 THEN
            exp_f := 125;
        ELSIF x =- 5725 THEN
            exp_f := 125;
        ELSIF x =- 5724 THEN
            exp_f := 125;
        ELSIF x =- 5723 THEN
            exp_f := 125;
        ELSIF x =- 5722 THEN
            exp_f := 126;
        ELSIF x =- 5721 THEN
            exp_f := 126;
        ELSIF x =- 5720 THEN
            exp_f := 126;
        ELSIF x =- 5719 THEN
            exp_f := 126;
        ELSIF x =- 5718 THEN
            exp_f := 126;
        ELSIF x =- 5717 THEN
            exp_f := 126;
        ELSIF x =- 5716 THEN
            exp_f := 126;
        ELSIF x =- 5715 THEN
            exp_f := 126;
        ELSIF x =- 5714 THEN
            exp_f := 126;
        ELSIF x =- 5713 THEN
            exp_f := 126;
        ELSIF x =- 5712 THEN
            exp_f := 126;
        ELSIF x =- 5711 THEN
            exp_f := 126;
        ELSIF x =- 5710 THEN
            exp_f := 126;
        ELSIF x =- 5709 THEN
            exp_f := 126;
        ELSIF x =- 5708 THEN
            exp_f := 126;
        ELSIF x =- 5707 THEN
            exp_f := 126;
        ELSIF x =- 5706 THEN
            exp_f := 126;
        ELSIF x =- 5705 THEN
            exp_f := 126;
        ELSIF x =- 5704 THEN
            exp_f := 126;
        ELSIF x =- 5703 THEN
            exp_f := 126;
        ELSIF x =- 5702 THEN
            exp_f := 127;
        ELSIF x =- 5701 THEN
            exp_f := 127;
        ELSIF x =- 5700 THEN
            exp_f := 127;
        ELSIF x =- 5699 THEN
            exp_f := 127;
        ELSIF x =- 5698 THEN
            exp_f := 127;
        ELSIF x =- 5697 THEN
            exp_f := 127;
        ELSIF x =- 5696 THEN
            exp_f := 127;
        ELSIF x =- 5695 THEN
            exp_f := 127;
        ELSIF x =- 5694 THEN
            exp_f := 127;
        ELSIF x =- 5693 THEN
            exp_f := 127;
        ELSIF x =- 5692 THEN
            exp_f := 127;
        ELSIF x =- 5691 THEN
            exp_f := 127;
        ELSIF x =- 5690 THEN
            exp_f := 127;
        ELSIF x =- 5689 THEN
            exp_f := 127;
        ELSIF x =- 5688 THEN
            exp_f := 127;
        ELSIF x =- 5687 THEN
            exp_f := 127;
        ELSIF x =- 5686 THEN
            exp_f := 127;
        ELSIF x =- 5685 THEN
            exp_f := 127;
        ELSIF x =- 5684 THEN
            exp_f := 127;
        ELSIF x =- 5683 THEN
            exp_f := 127;
        ELSIF x =- 5682 THEN
            exp_f := 128;
        ELSIF x =- 5681 THEN
            exp_f := 128;
        ELSIF x =- 5680 THEN
            exp_f := 128;
        ELSIF x =- 5679 THEN
            exp_f := 128;
        ELSIF x =- 5678 THEN
            exp_f := 128;
        ELSIF x =- 5677 THEN
            exp_f := 128;
        ELSIF x =- 5676 THEN
            exp_f := 128;
        ELSIF x =- 5675 THEN
            exp_f := 128;
        ELSIF x =- 5674 THEN
            exp_f := 128;
        ELSIF x =- 5673 THEN
            exp_f := 128;
        ELSIF x =- 5672 THEN
            exp_f := 128;
        ELSIF x =- 5671 THEN
            exp_f := 128;
        ELSIF x =- 5670 THEN
            exp_f := 128;
        ELSIF x =- 5669 THEN
            exp_f := 128;
        ELSIF x =- 5668 THEN
            exp_f := 128;
        ELSIF x =- 5667 THEN
            exp_f := 128;
        ELSIF x =- 5666 THEN
            exp_f := 128;
        ELSIF x =- 5665 THEN
            exp_f := 128;
        ELSIF x =- 5664 THEN
            exp_f := 128;
        ELSIF x =- 5663 THEN
            exp_f := 128;
        ELSIF x =- 5662 THEN
            exp_f := 129;
        ELSIF x =- 5661 THEN
            exp_f := 129;
        ELSIF x =- 5660 THEN
            exp_f := 129;
        ELSIF x =- 5659 THEN
            exp_f := 129;
        ELSIF x =- 5658 THEN
            exp_f := 129;
        ELSIF x =- 5657 THEN
            exp_f := 129;
        ELSIF x =- 5656 THEN
            exp_f := 129;
        ELSIF x =- 5655 THEN
            exp_f := 129;
        ELSIF x =- 5654 THEN
            exp_f := 129;
        ELSIF x =- 5653 THEN
            exp_f := 129;
        ELSIF x =- 5652 THEN
            exp_f := 129;
        ELSIF x =- 5651 THEN
            exp_f := 129;
        ELSIF x =- 5650 THEN
            exp_f := 129;
        ELSIF x =- 5649 THEN
            exp_f := 129;
        ELSIF x =- 5648 THEN
            exp_f := 129;
        ELSIF x =- 5647 THEN
            exp_f := 129;
        ELSIF x =- 5646 THEN
            exp_f := 129;
        ELSIF x =- 5645 THEN
            exp_f := 129;
        ELSIF x =- 5644 THEN
            exp_f := 129;
        ELSIF x =- 5643 THEN
            exp_f := 129;
        ELSIF x =- 5642 THEN
            exp_f := 130;
        ELSIF x =- 5641 THEN
            exp_f := 130;
        ELSIF x =- 5640 THEN
            exp_f := 130;
        ELSIF x =- 5639 THEN
            exp_f := 130;
        ELSIF x =- 5638 THEN
            exp_f := 130;
        ELSIF x =- 5637 THEN
            exp_f := 130;
        ELSIF x =- 5636 THEN
            exp_f := 130;
        ELSIF x =- 5635 THEN
            exp_f := 130;
        ELSIF x =- 5634 THEN
            exp_f := 130;
        ELSIF x =- 5633 THEN
            exp_f := 130;
        ELSIF x =- 5632 THEN
            exp_f := 130;
        ELSIF x =- 5631 THEN
            exp_f := 130;
        ELSIF x =- 5630 THEN
            exp_f := 130;
        ELSIF x =- 5629 THEN
            exp_f := 130;
        ELSIF x =- 5628 THEN
            exp_f := 130;
        ELSIF x =- 5627 THEN
            exp_f := 131;
        ELSIF x =- 5626 THEN
            exp_f := 131;
        ELSIF x =- 5625 THEN
            exp_f := 131;
        ELSIF x =- 5624 THEN
            exp_f := 131;
        ELSIF x =- 5623 THEN
            exp_f := 131;
        ELSIF x =- 5622 THEN
            exp_f := 131;
        ELSIF x =- 5621 THEN
            exp_f := 131;
        ELSIF x =- 5620 THEN
            exp_f := 131;
        ELSIF x =- 5619 THEN
            exp_f := 131;
        ELSIF x =- 5618 THEN
            exp_f := 131;
        ELSIF x =- 5617 THEN
            exp_f := 131;
        ELSIF x =- 5616 THEN
            exp_f := 131;
        ELSIF x =- 5615 THEN
            exp_f := 131;
        ELSIF x =- 5614 THEN
            exp_f := 131;
        ELSIF x =- 5613 THEN
            exp_f := 131;
        ELSIF x =- 5612 THEN
            exp_f := 131;
        ELSIF x =- 5611 THEN
            exp_f := 133;
        ELSIF x =- 5610 THEN
            exp_f := 133;
        ELSIF x =- 5609 THEN
            exp_f := 133;
        ELSIF x =- 5608 THEN
            exp_f := 133;
        ELSIF x =- 5607 THEN
            exp_f := 133;
        ELSIF x =- 5606 THEN
            exp_f := 133;
        ELSIF x =- 5605 THEN
            exp_f := 133;
        ELSIF x =- 5604 THEN
            exp_f := 133;
        ELSIF x =- 5603 THEN
            exp_f := 133;
        ELSIF x =- 5602 THEN
            exp_f := 133;
        ELSIF x =- 5601 THEN
            exp_f := 133;
        ELSIF x =- 5600 THEN
            exp_f := 133;
        ELSIF x =- 5599 THEN
            exp_f := 133;
        ELSIF x =- 5598 THEN
            exp_f := 133;
        ELSIF x =- 5597 THEN
            exp_f := 133;
        ELSIF x =- 5596 THEN
            exp_f := 133;
        ELSIF x =- 5595 THEN
            exp_f := 134;
        ELSIF x =- 5594 THEN
            exp_f := 134;
        ELSIF x =- 5593 THEN
            exp_f := 134;
        ELSIF x =- 5592 THEN
            exp_f := 134;
        ELSIF x =- 5591 THEN
            exp_f := 134;
        ELSIF x =- 5590 THEN
            exp_f := 134;
        ELSIF x =- 5589 THEN
            exp_f := 134;
        ELSIF x =- 5588 THEN
            exp_f := 134;
        ELSIF x =- 5587 THEN
            exp_f := 134;
        ELSIF x =- 5586 THEN
            exp_f := 134;
        ELSIF x =- 5585 THEN
            exp_f := 134;
        ELSIF x =- 5584 THEN
            exp_f := 134;
        ELSIF x =- 5583 THEN
            exp_f := 134;
        ELSIF x =- 5582 THEN
            exp_f := 134;
        ELSIF x =- 5581 THEN
            exp_f := 134;
        ELSIF x =- 5580 THEN
            exp_f := 134;
        ELSIF x =- 5579 THEN
            exp_f := 135;
        ELSIF x =- 5578 THEN
            exp_f := 135;
        ELSIF x =- 5577 THEN
            exp_f := 135;
        ELSIF x =- 5576 THEN
            exp_f := 135;
        ELSIF x =- 5575 THEN
            exp_f := 135;
        ELSIF x =- 5574 THEN
            exp_f := 135;
        ELSIF x =- 5573 THEN
            exp_f := 135;
        ELSIF x =- 5572 THEN
            exp_f := 135;
        ELSIF x =- 5571 THEN
            exp_f := 135;
        ELSIF x =- 5570 THEN
            exp_f := 135;
        ELSIF x =- 5569 THEN
            exp_f := 135;
        ELSIF x =- 5568 THEN
            exp_f := 135;
        ELSIF x =- 5567 THEN
            exp_f := 135;
        ELSIF x =- 5566 THEN
            exp_f := 135;
        ELSIF x =- 5565 THEN
            exp_f := 135;
        ELSIF x =- 5564 THEN
            exp_f := 135;
        ELSIF x =- 5563 THEN
            exp_f := 136;
        ELSIF x =- 5562 THEN
            exp_f := 136;
        ELSIF x =- 5561 THEN
            exp_f := 136;
        ELSIF x =- 5560 THEN
            exp_f := 136;
        ELSIF x =- 5559 THEN
            exp_f := 136;
        ELSIF x =- 5558 THEN
            exp_f := 136;
        ELSIF x =- 5557 THEN
            exp_f := 136;
        ELSIF x =- 5556 THEN
            exp_f := 136;
        ELSIF x =- 5555 THEN
            exp_f := 136;
        ELSIF x =- 5554 THEN
            exp_f := 136;
        ELSIF x =- 5553 THEN
            exp_f := 136;
        ELSIF x =- 5552 THEN
            exp_f := 136;
        ELSIF x =- 5551 THEN
            exp_f := 136;
        ELSIF x =- 5550 THEN
            exp_f := 136;
        ELSIF x =- 5549 THEN
            exp_f := 136;
        ELSIF x =- 5548 THEN
            exp_f := 136;
        ELSIF x =- 5547 THEN
            exp_f := 137;
        ELSIF x =- 5546 THEN
            exp_f := 137;
        ELSIF x =- 5545 THEN
            exp_f := 137;
        ELSIF x =- 5544 THEN
            exp_f := 137;
        ELSIF x =- 5543 THEN
            exp_f := 137;
        ELSIF x =- 5542 THEN
            exp_f := 137;
        ELSIF x =- 5541 THEN
            exp_f := 137;
        ELSIF x =- 5540 THEN
            exp_f := 137;
        ELSIF x =- 5539 THEN
            exp_f := 137;
        ELSIF x =- 5538 THEN
            exp_f := 137;
        ELSIF x =- 5537 THEN
            exp_f := 137;
        ELSIF x =- 5536 THEN
            exp_f := 137;
        ELSIF x =- 5535 THEN
            exp_f := 137;
        ELSIF x =- 5534 THEN
            exp_f := 137;
        ELSIF x =- 5533 THEN
            exp_f := 137;
        ELSIF x =- 5532 THEN
            exp_f := 137;
        ELSIF x =- 5531 THEN
            exp_f := 138;
        ELSIF x =- 5530 THEN
            exp_f := 138;
        ELSIF x =- 5529 THEN
            exp_f := 138;
        ELSIF x =- 5528 THEN
            exp_f := 138;
        ELSIF x =- 5527 THEN
            exp_f := 138;
        ELSIF x =- 5526 THEN
            exp_f := 138;
        ELSIF x =- 5525 THEN
            exp_f := 138;
        ELSIF x =- 5524 THEN
            exp_f := 138;
        ELSIF x =- 5523 THEN
            exp_f := 138;
        ELSIF x =- 5522 THEN
            exp_f := 138;
        ELSIF x =- 5521 THEN
            exp_f := 138;
        ELSIF x =- 5520 THEN
            exp_f := 138;
        ELSIF x =- 5519 THEN
            exp_f := 138;
        ELSIF x =- 5518 THEN
            exp_f := 138;
        ELSIF x =- 5517 THEN
            exp_f := 138;
        ELSIF x =- 5516 THEN
            exp_f := 138;
        ELSIF x =- 5515 THEN
            exp_f := 139;
        ELSIF x =- 5514 THEN
            exp_f := 139;
        ELSIF x =- 5513 THEN
            exp_f := 139;
        ELSIF x =- 5512 THEN
            exp_f := 139;
        ELSIF x =- 5511 THEN
            exp_f := 139;
        ELSIF x =- 5510 THEN
            exp_f := 139;
        ELSIF x =- 5509 THEN
            exp_f := 139;
        ELSIF x =- 5508 THEN
            exp_f := 139;
        ELSIF x =- 5507 THEN
            exp_f := 139;
        ELSIF x =- 5506 THEN
            exp_f := 139;
        ELSIF x =- 5505 THEN
            exp_f := 139;
        ELSIF x =- 5504 THEN
            exp_f := 139;
        ELSIF x =- 5503 THEN
            exp_f := 139;
        ELSIF x =- 5502 THEN
            exp_f := 139;
        ELSIF x =- 5501 THEN
            exp_f := 139;
        ELSIF x =- 5500 THEN
            exp_f := 139;
        ELSIF x =- 5499 THEN
            exp_f := 139;
        ELSIF x =- 5498 THEN
            exp_f := 141;
        ELSIF x =- 5497 THEN
            exp_f := 141;
        ELSIF x =- 5496 THEN
            exp_f := 141;
        ELSIF x =- 5495 THEN
            exp_f := 141;
        ELSIF x =- 5494 THEN
            exp_f := 141;
        ELSIF x =- 5493 THEN
            exp_f := 141;
        ELSIF x =- 5492 THEN
            exp_f := 141;
        ELSIF x =- 5491 THEN
            exp_f := 141;
        ELSIF x =- 5490 THEN
            exp_f := 141;
        ELSIF x =- 5489 THEN
            exp_f := 141;
        ELSIF x =- 5488 THEN
            exp_f := 141;
        ELSIF x =- 5487 THEN
            exp_f := 141;
        ELSIF x =- 5486 THEN
            exp_f := 141;
        ELSIF x =- 5485 THEN
            exp_f := 141;
        ELSIF x =- 5484 THEN
            exp_f := 141;
        ELSIF x =- 5483 THEN
            exp_f := 141;
        ELSIF x =- 5482 THEN
            exp_f := 142;
        ELSIF x =- 5481 THEN
            exp_f := 142;
        ELSIF x =- 5480 THEN
            exp_f := 142;
        ELSIF x =- 5479 THEN
            exp_f := 142;
        ELSIF x =- 5478 THEN
            exp_f := 142;
        ELSIF x =- 5477 THEN
            exp_f := 142;
        ELSIF x =- 5476 THEN
            exp_f := 142;
        ELSIF x =- 5475 THEN
            exp_f := 142;
        ELSIF x =- 5474 THEN
            exp_f := 142;
        ELSIF x =- 5473 THEN
            exp_f := 142;
        ELSIF x =- 5472 THEN
            exp_f := 142;
        ELSIF x =- 5471 THEN
            exp_f := 142;
        ELSIF x =- 5470 THEN
            exp_f := 142;
        ELSIF x =- 5469 THEN
            exp_f := 142;
        ELSIF x =- 5468 THEN
            exp_f := 142;
        ELSIF x =- 5467 THEN
            exp_f := 142;
        ELSIF x =- 5466 THEN
            exp_f := 143;
        ELSIF x =- 5465 THEN
            exp_f := 143;
        ELSIF x =- 5464 THEN
            exp_f := 143;
        ELSIF x =- 5463 THEN
            exp_f := 143;
        ELSIF x =- 5462 THEN
            exp_f := 143;
        ELSIF x =- 5461 THEN
            exp_f := 143;
        ELSIF x =- 5460 THEN
            exp_f := 143;
        ELSIF x =- 5459 THEN
            exp_f := 143;
        ELSIF x =- 5458 THEN
            exp_f := 143;
        ELSIF x =- 5457 THEN
            exp_f := 143;
        ELSIF x =- 5456 THEN
            exp_f := 143;
        ELSIF x =- 5455 THEN
            exp_f := 143;
        ELSIF x =- 5454 THEN
            exp_f := 143;
        ELSIF x =- 5453 THEN
            exp_f := 143;
        ELSIF x =- 5452 THEN
            exp_f := 143;
        ELSIF x =- 5451 THEN
            exp_f := 143;
        ELSIF x =- 5450 THEN
            exp_f := 144;
        ELSIF x =- 5449 THEN
            exp_f := 144;
        ELSIF x =- 5448 THEN
            exp_f := 144;
        ELSIF x =- 5447 THEN
            exp_f := 144;
        ELSIF x =- 5446 THEN
            exp_f := 144;
        ELSIF x =- 5445 THEN
            exp_f := 144;
        ELSIF x =- 5444 THEN
            exp_f := 144;
        ELSIF x =- 5443 THEN
            exp_f := 144;
        ELSIF x =- 5442 THEN
            exp_f := 144;
        ELSIF x =- 5441 THEN
            exp_f := 144;
        ELSIF x =- 5440 THEN
            exp_f := 144;
        ELSIF x =- 5439 THEN
            exp_f := 144;
        ELSIF x =- 5438 THEN
            exp_f := 144;
        ELSIF x =- 5437 THEN
            exp_f := 144;
        ELSIF x =- 5436 THEN
            exp_f := 144;
        ELSIF x =- 5435 THEN
            exp_f := 144;
        ELSIF x =- 5434 THEN
            exp_f := 145;
        ELSIF x =- 5433 THEN
            exp_f := 145;
        ELSIF x =- 5432 THEN
            exp_f := 145;
        ELSIF x =- 5431 THEN
            exp_f := 145;
        ELSIF x =- 5430 THEN
            exp_f := 145;
        ELSIF x =- 5429 THEN
            exp_f := 145;
        ELSIF x =- 5428 THEN
            exp_f := 145;
        ELSIF x =- 5427 THEN
            exp_f := 145;
        ELSIF x =- 5426 THEN
            exp_f := 145;
        ELSIF x =- 5425 THEN
            exp_f := 145;
        ELSIF x =- 5424 THEN
            exp_f := 145;
        ELSIF x =- 5423 THEN
            exp_f := 145;
        ELSIF x =- 5422 THEN
            exp_f := 145;
        ELSIF x =- 5421 THEN
            exp_f := 145;
        ELSIF x =- 5420 THEN
            exp_f := 145;
        ELSIF x =- 5419 THEN
            exp_f := 145;
        ELSIF x =- 5418 THEN
            exp_f := 146;
        ELSIF x =- 5417 THEN
            exp_f := 146;
        ELSIF x =- 5416 THEN
            exp_f := 146;
        ELSIF x =- 5415 THEN
            exp_f := 146;
        ELSIF x =- 5414 THEN
            exp_f := 146;
        ELSIF x =- 5413 THEN
            exp_f := 146;
        ELSIF x =- 5412 THEN
            exp_f := 146;
        ELSIF x =- 5411 THEN
            exp_f := 146;
        ELSIF x =- 5410 THEN
            exp_f := 146;
        ELSIF x =- 5409 THEN
            exp_f := 146;
        ELSIF x =- 5408 THEN
            exp_f := 146;
        ELSIF x =- 5407 THEN
            exp_f := 146;
        ELSIF x =- 5406 THEN
            exp_f := 146;
        ELSIF x =- 5405 THEN
            exp_f := 146;
        ELSIF x =- 5404 THEN
            exp_f := 146;
        ELSIF x =- 5403 THEN
            exp_f := 146;
        ELSIF x =- 5402 THEN
            exp_f := 147;
        ELSIF x =- 5401 THEN
            exp_f := 147;
        ELSIF x =- 5400 THEN
            exp_f := 147;
        ELSIF x =- 5399 THEN
            exp_f := 147;
        ELSIF x =- 5398 THEN
            exp_f := 147;
        ELSIF x =- 5397 THEN
            exp_f := 147;
        ELSIF x =- 5396 THEN
            exp_f := 147;
        ELSIF x =- 5395 THEN
            exp_f := 147;
        ELSIF x =- 5394 THEN
            exp_f := 147;
        ELSIF x =- 5393 THEN
            exp_f := 147;
        ELSIF x =- 5392 THEN
            exp_f := 147;
        ELSIF x =- 5391 THEN
            exp_f := 147;
        ELSIF x =- 5390 THEN
            exp_f := 147;
        ELSIF x =- 5389 THEN
            exp_f := 147;
        ELSIF x =- 5388 THEN
            exp_f := 147;
        ELSIF x =- 5387 THEN
            exp_f := 147;
        ELSIF x =- 5386 THEN
            exp_f := 149;
        ELSIF x =- 5385 THEN
            exp_f := 149;
        ELSIF x =- 5384 THEN
            exp_f := 149;
        ELSIF x =- 5383 THEN
            exp_f := 149;
        ELSIF x =- 5382 THEN
            exp_f := 149;
        ELSIF x =- 5381 THEN
            exp_f := 149;
        ELSIF x =- 5380 THEN
            exp_f := 149;
        ELSIF x =- 5379 THEN
            exp_f := 149;
        ELSIF x =- 5378 THEN
            exp_f := 149;
        ELSIF x =- 5377 THEN
            exp_f := 149;
        ELSIF x =- 5376 THEN
            exp_f := 149;
        ELSIF x =- 5375 THEN
            exp_f := 149;
        ELSIF x =- 5374 THEN
            exp_f := 149;
        ELSIF x =- 5373 THEN
            exp_f := 149;
        ELSIF x =- 5372 THEN
            exp_f := 149;
        ELSIF x =- 5371 THEN
            exp_f := 149;
        ELSIF x =- 5370 THEN
            exp_f := 149;
        ELSIF x =- 5369 THEN
            exp_f := 150;
        ELSIF x =- 5368 THEN
            exp_f := 150;
        ELSIF x =- 5367 THEN
            exp_f := 150;
        ELSIF x =- 5366 THEN
            exp_f := 150;
        ELSIF x =- 5365 THEN
            exp_f := 150;
        ELSIF x =- 5364 THEN
            exp_f := 150;
        ELSIF x =- 5363 THEN
            exp_f := 150;
        ELSIF x =- 5362 THEN
            exp_f := 150;
        ELSIF x =- 5361 THEN
            exp_f := 150;
        ELSIF x =- 5360 THEN
            exp_f := 150;
        ELSIF x =- 5359 THEN
            exp_f := 150;
        ELSIF x =- 5358 THEN
            exp_f := 150;
        ELSIF x =- 5357 THEN
            exp_f := 150;
        ELSIF x =- 5356 THEN
            exp_f := 150;
        ELSIF x =- 5355 THEN
            exp_f := 150;
        ELSIF x =- 5354 THEN
            exp_f := 150;
        ELSIF x =- 5353 THEN
            exp_f := 151;
        ELSIF x =- 5352 THEN
            exp_f := 151;
        ELSIF x =- 5351 THEN
            exp_f := 151;
        ELSIF x =- 5350 THEN
            exp_f := 151;
        ELSIF x =- 5349 THEN
            exp_f := 151;
        ELSIF x =- 5348 THEN
            exp_f := 151;
        ELSIF x =- 5347 THEN
            exp_f := 151;
        ELSIF x =- 5346 THEN
            exp_f := 151;
        ELSIF x =- 5345 THEN
            exp_f := 151;
        ELSIF x =- 5344 THEN
            exp_f := 151;
        ELSIF x =- 5343 THEN
            exp_f := 151;
        ELSIF x =- 5342 THEN
            exp_f := 151;
        ELSIF x =- 5341 THEN
            exp_f := 151;
        ELSIF x =- 5340 THEN
            exp_f := 151;
        ELSIF x =- 5339 THEN
            exp_f := 151;
        ELSIF x =- 5338 THEN
            exp_f := 151;
        ELSIF x =- 5337 THEN
            exp_f := 152;
        ELSIF x =- 5336 THEN
            exp_f := 152;
        ELSIF x =- 5335 THEN
            exp_f := 152;
        ELSIF x =- 5334 THEN
            exp_f := 152;
        ELSIF x =- 5333 THEN
            exp_f := 152;
        ELSIF x =- 5332 THEN
            exp_f := 152;
        ELSIF x =- 5331 THEN
            exp_f := 152;
        ELSIF x =- 5330 THEN
            exp_f := 152;
        ELSIF x =- 5329 THEN
            exp_f := 152;
        ELSIF x =- 5328 THEN
            exp_f := 152;
        ELSIF x =- 5327 THEN
            exp_f := 152;
        ELSIF x =- 5326 THEN
            exp_f := 152;
        ELSIF x =- 5325 THEN
            exp_f := 152;
        ELSIF x =- 5324 THEN
            exp_f := 152;
        ELSIF x =- 5323 THEN
            exp_f := 152;
        ELSIF x =- 5322 THEN
            exp_f := 152;
        ELSIF x =- 5321 THEN
            exp_f := 153;
        ELSIF x =- 5320 THEN
            exp_f := 153;
        ELSIF x =- 5319 THEN
            exp_f := 153;
        ELSIF x =- 5318 THEN
            exp_f := 153;
        ELSIF x =- 5317 THEN
            exp_f := 153;
        ELSIF x =- 5316 THEN
            exp_f := 153;
        ELSIF x =- 5315 THEN
            exp_f := 153;
        ELSIF x =- 5314 THEN
            exp_f := 153;
        ELSIF x =- 5313 THEN
            exp_f := 153;
        ELSIF x =- 5312 THEN
            exp_f := 153;
        ELSIF x =- 5311 THEN
            exp_f := 153;
        ELSIF x =- 5310 THEN
            exp_f := 153;
        ELSIF x =- 5309 THEN
            exp_f := 153;
        ELSIF x =- 5308 THEN
            exp_f := 153;
        ELSIF x =- 5307 THEN
            exp_f := 153;
        ELSIF x =- 5306 THEN
            exp_f := 153;
        ELSIF x =- 5305 THEN
            exp_f := 154;
        ELSIF x =- 5304 THEN
            exp_f := 154;
        ELSIF x =- 5303 THEN
            exp_f := 154;
        ELSIF x =- 5302 THEN
            exp_f := 154;
        ELSIF x =- 5301 THEN
            exp_f := 154;
        ELSIF x =- 5300 THEN
            exp_f := 154;
        ELSIF x =- 5299 THEN
            exp_f := 154;
        ELSIF x =- 5298 THEN
            exp_f := 154;
        ELSIF x =- 5297 THEN
            exp_f := 154;
        ELSIF x =- 5296 THEN
            exp_f := 154;
        ELSIF x =- 5295 THEN
            exp_f := 154;
        ELSIF x =- 5294 THEN
            exp_f := 154;
        ELSIF x =- 5293 THEN
            exp_f := 154;
        ELSIF x =- 5292 THEN
            exp_f := 154;
        ELSIF x =- 5291 THEN
            exp_f := 154;
        ELSIF x =- 5290 THEN
            exp_f := 154;
        ELSIF x =- 5289 THEN
            exp_f := 156;
        ELSIF x =- 5288 THEN
            exp_f := 156;
        ELSIF x =- 5287 THEN
            exp_f := 156;
        ELSIF x =- 5286 THEN
            exp_f := 156;
        ELSIF x =- 5285 THEN
            exp_f := 156;
        ELSIF x =- 5284 THEN
            exp_f := 156;
        ELSIF x =- 5283 THEN
            exp_f := 156;
        ELSIF x =- 5282 THEN
            exp_f := 156;
        ELSIF x =- 5281 THEN
            exp_f := 156;
        ELSIF x =- 5280 THEN
            exp_f := 156;
        ELSIF x =- 5279 THEN
            exp_f := 156;
        ELSIF x =- 5278 THEN
            exp_f := 156;
        ELSIF x =- 5277 THEN
            exp_f := 156;
        ELSIF x =- 5276 THEN
            exp_f := 156;
        ELSIF x =- 5275 THEN
            exp_f := 156;
        ELSIF x =- 5274 THEN
            exp_f := 156;
        ELSIF x =- 5273 THEN
            exp_f := 157;
        ELSIF x =- 5272 THEN
            exp_f := 157;
        ELSIF x =- 5271 THEN
            exp_f := 157;
        ELSIF x =- 5270 THEN
            exp_f := 157;
        ELSIF x =- 5269 THEN
            exp_f := 157;
        ELSIF x =- 5268 THEN
            exp_f := 157;
        ELSIF x =- 5267 THEN
            exp_f := 157;
        ELSIF x =- 5266 THEN
            exp_f := 157;
        ELSIF x =- 5265 THEN
            exp_f := 157;
        ELSIF x =- 5264 THEN
            exp_f := 157;
        ELSIF x =- 5263 THEN
            exp_f := 157;
        ELSIF x =- 5262 THEN
            exp_f := 157;
        ELSIF x =- 5261 THEN
            exp_f := 157;
        ELSIF x =- 5260 THEN
            exp_f := 157;
        ELSIF x =- 5259 THEN
            exp_f := 157;
        ELSIF x =- 5258 THEN
            exp_f := 157;
        ELSIF x =- 5257 THEN
            exp_f := 158;
        ELSIF x =- 5256 THEN
            exp_f := 158;
        ELSIF x =- 5255 THEN
            exp_f := 158;
        ELSIF x =- 5254 THEN
            exp_f := 158;
        ELSIF x =- 5253 THEN
            exp_f := 158;
        ELSIF x =- 5252 THEN
            exp_f := 158;
        ELSIF x =- 5251 THEN
            exp_f := 158;
        ELSIF x =- 5250 THEN
            exp_f := 158;
        ELSIF x =- 5249 THEN
            exp_f := 158;
        ELSIF x =- 5248 THEN
            exp_f := 158;
        ELSIF x =- 5247 THEN
            exp_f := 158;
        ELSIF x =- 5246 THEN
            exp_f := 158;
        ELSIF x =- 5245 THEN
            exp_f := 158;
        ELSIF x =- 5244 THEN
            exp_f := 158;
        ELSIF x =- 5243 THEN
            exp_f := 158;
        ELSIF x =- 5242 THEN
            exp_f := 158;
        ELSIF x =- 5241 THEN
            exp_f := 158;
        ELSIF x =- 5240 THEN
            exp_f := 159;
        ELSIF x =- 5239 THEN
            exp_f := 159;
        ELSIF x =- 5238 THEN
            exp_f := 159;
        ELSIF x =- 5237 THEN
            exp_f := 159;
        ELSIF x =- 5236 THEN
            exp_f := 159;
        ELSIF x =- 5235 THEN
            exp_f := 159;
        ELSIF x =- 5234 THEN
            exp_f := 159;
        ELSIF x =- 5233 THEN
            exp_f := 159;
        ELSIF x =- 5232 THEN
            exp_f := 159;
        ELSIF x =- 5231 THEN
            exp_f := 159;
        ELSIF x =- 5230 THEN
            exp_f := 159;
        ELSIF x =- 5229 THEN
            exp_f := 159;
        ELSIF x =- 5228 THEN
            exp_f := 159;
        ELSIF x =- 5227 THEN
            exp_f := 159;
        ELSIF x =- 5226 THEN
            exp_f := 159;
        ELSIF x =- 5225 THEN
            exp_f := 159;
        ELSIF x =- 5224 THEN
            exp_f := 160;
        ELSIF x =- 5223 THEN
            exp_f := 160;
        ELSIF x =- 5222 THEN
            exp_f := 160;
        ELSIF x =- 5221 THEN
            exp_f := 160;
        ELSIF x =- 5220 THEN
            exp_f := 160;
        ELSIF x =- 5219 THEN
            exp_f := 160;
        ELSIF x =- 5218 THEN
            exp_f := 160;
        ELSIF x =- 5217 THEN
            exp_f := 160;
        ELSIF x =- 5216 THEN
            exp_f := 160;
        ELSIF x =- 5215 THEN
            exp_f := 160;
        ELSIF x =- 5214 THEN
            exp_f := 160;
        ELSIF x =- 5213 THEN
            exp_f := 160;
        ELSIF x =- 5212 THEN
            exp_f := 160;
        ELSIF x =- 5211 THEN
            exp_f := 160;
        ELSIF x =- 5210 THEN
            exp_f := 160;
        ELSIF x =- 5209 THEN
            exp_f := 160;
        ELSIF x =- 5208 THEN
            exp_f := 161;
        ELSIF x =- 5207 THEN
            exp_f := 161;
        ELSIF x =- 5206 THEN
            exp_f := 161;
        ELSIF x =- 5205 THEN
            exp_f := 161;
        ELSIF x =- 5204 THEN
            exp_f := 161;
        ELSIF x =- 5203 THEN
            exp_f := 161;
        ELSIF x =- 5202 THEN
            exp_f := 161;
        ELSIF x =- 5201 THEN
            exp_f := 161;
        ELSIF x =- 5200 THEN
            exp_f := 161;
        ELSIF x =- 5199 THEN
            exp_f := 161;
        ELSIF x =- 5198 THEN
            exp_f := 161;
        ELSIF x =- 5197 THEN
            exp_f := 161;
        ELSIF x =- 5196 THEN
            exp_f := 161;
        ELSIF x =- 5195 THEN
            exp_f := 161;
        ELSIF x =- 5194 THEN
            exp_f := 161;
        ELSIF x =- 5193 THEN
            exp_f := 161;
        ELSIF x =- 5192 THEN
            exp_f := 163;
        ELSIF x =- 5191 THEN
            exp_f := 163;
        ELSIF x =- 5190 THEN
            exp_f := 163;
        ELSIF x =- 5189 THEN
            exp_f := 163;
        ELSIF x =- 5188 THEN
            exp_f := 163;
        ELSIF x =- 5187 THEN
            exp_f := 163;
        ELSIF x =- 5186 THEN
            exp_f := 163;
        ELSIF x =- 5185 THEN
            exp_f := 163;
        ELSIF x =- 5184 THEN
            exp_f := 163;
        ELSIF x =- 5183 THEN
            exp_f := 163;
        ELSIF x =- 5182 THEN
            exp_f := 163;
        ELSIF x =- 5181 THEN
            exp_f := 163;
        ELSIF x =- 5180 THEN
            exp_f := 163;
        ELSIF x =- 5179 THEN
            exp_f := 163;
        ELSIF x =- 5178 THEN
            exp_f := 163;
        ELSIF x =- 5177 THEN
            exp_f := 163;
        ELSIF x =- 5176 THEN
            exp_f := 164;
        ELSIF x =- 5175 THEN
            exp_f := 164;
        ELSIF x =- 5174 THEN
            exp_f := 164;
        ELSIF x =- 5173 THEN
            exp_f := 164;
        ELSIF x =- 5172 THEN
            exp_f := 164;
        ELSIF x =- 5171 THEN
            exp_f := 164;
        ELSIF x =- 5170 THEN
            exp_f := 164;
        ELSIF x =- 5169 THEN
            exp_f := 164;
        ELSIF x =- 5168 THEN
            exp_f := 164;
        ELSIF x =- 5167 THEN
            exp_f := 164;
        ELSIF x =- 5166 THEN
            exp_f := 164;
        ELSIF x =- 5165 THEN
            exp_f := 164;
        ELSIF x =- 5164 THEN
            exp_f := 164;
        ELSIF x =- 5163 THEN
            exp_f := 164;
        ELSIF x =- 5162 THEN
            exp_f := 164;
        ELSIF x =- 5161 THEN
            exp_f := 164;
        ELSIF x =- 5160 THEN
            exp_f := 165;
        ELSIF x =- 5159 THEN
            exp_f := 165;
        ELSIF x =- 5158 THEN
            exp_f := 165;
        ELSIF x =- 5157 THEN
            exp_f := 165;
        ELSIF x =- 5156 THEN
            exp_f := 165;
        ELSIF x =- 5155 THEN
            exp_f := 165;
        ELSIF x =- 5154 THEN
            exp_f := 165;
        ELSIF x =- 5153 THEN
            exp_f := 165;
        ELSIF x =- 5152 THEN
            exp_f := 165;
        ELSIF x =- 5151 THEN
            exp_f := 165;
        ELSIF x =- 5150 THEN
            exp_f := 165;
        ELSIF x =- 5149 THEN
            exp_f := 165;
        ELSIF x =- 5148 THEN
            exp_f := 165;
        ELSIF x =- 5147 THEN
            exp_f := 165;
        ELSIF x =- 5146 THEN
            exp_f := 165;
        ELSIF x =- 5145 THEN
            exp_f := 165;
        ELSIF x =- 5144 THEN
            exp_f := 166;
        ELSIF x =- 5143 THEN
            exp_f := 166;
        ELSIF x =- 5142 THEN
            exp_f := 166;
        ELSIF x =- 5141 THEN
            exp_f := 166;
        ELSIF x =- 5140 THEN
            exp_f := 166;
        ELSIF x =- 5139 THEN
            exp_f := 166;
        ELSIF x =- 5138 THEN
            exp_f := 166;
        ELSIF x =- 5137 THEN
            exp_f := 166;
        ELSIF x =- 5136 THEN
            exp_f := 166;
        ELSIF x =- 5135 THEN
            exp_f := 166;
        ELSIF x =- 5134 THEN
            exp_f := 166;
        ELSIF x =- 5133 THEN
            exp_f := 166;
        ELSIF x =- 5132 THEN
            exp_f := 166;
        ELSIF x =- 5131 THEN
            exp_f := 166;
        ELSIF x =- 5130 THEN
            exp_f := 166;
        ELSIF x =- 5129 THEN
            exp_f := 166;
        ELSIF x =- 5128 THEN
            exp_f := 167;
        ELSIF x =- 5127 THEN
            exp_f := 167;
        ELSIF x =- 5126 THEN
            exp_f := 167;
        ELSIF x =- 5125 THEN
            exp_f := 167;
        ELSIF x =- 5124 THEN
            exp_f := 167;
        ELSIF x =- 5123 THEN
            exp_f := 167;
        ELSIF x =- 5122 THEN
            exp_f := 167;
        ELSIF x =- 5121 THEN
            exp_f := 167;
        ELSIF x =- 5120 THEN
            exp_f := 167;
        ELSIF x =- 5119 THEN
            exp_f := 167;
        ELSIF x =- 5118 THEN
            exp_f := 167;
        ELSIF x =- 5117 THEN
            exp_f := 167;
        ELSIF x =- 5116 THEN
            exp_f := 167;
        ELSIF x =- 5115 THEN
            exp_f := 167;
        ELSIF x =- 5114 THEN
            exp_f := 167;
        ELSIF x =- 5113 THEN
            exp_f := 168;
        ELSIF x =- 5112 THEN
            exp_f := 168;
        ELSIF x =- 5111 THEN
            exp_f := 168;
        ELSIF x =- 5110 THEN
            exp_f := 168;
        ELSIF x =- 5109 THEN
            exp_f := 168;
        ELSIF x =- 5108 THEN
            exp_f := 168;
        ELSIF x =- 5107 THEN
            exp_f := 168;
        ELSIF x =- 5106 THEN
            exp_f := 168;
        ELSIF x =- 5105 THEN
            exp_f := 168;
        ELSIF x =- 5104 THEN
            exp_f := 168;
        ELSIF x =- 5103 THEN
            exp_f := 168;
        ELSIF x =- 5102 THEN
            exp_f := 168;
        ELSIF x =- 5101 THEN
            exp_f := 168;
        ELSIF x =- 5100 THEN
            exp_f := 170;
        ELSIF x =- 5099 THEN
            exp_f := 170;
        ELSIF x =- 5098 THEN
            exp_f := 170;
        ELSIF x =- 5097 THEN
            exp_f := 170;
        ELSIF x =- 5096 THEN
            exp_f := 170;
        ELSIF x =- 5095 THEN
            exp_f := 170;
        ELSIF x =- 5094 THEN
            exp_f := 170;
        ELSIF x =- 5093 THEN
            exp_f := 170;
        ELSIF x =- 5092 THEN
            exp_f := 170;
        ELSIF x =- 5091 THEN
            exp_f := 170;
        ELSIF x =- 5090 THEN
            exp_f := 170;
        ELSIF x =- 5089 THEN
            exp_f := 170;
        ELSIF x =- 5088 THEN
            exp_f := 171;
        ELSIF x =- 5087 THEN
            exp_f := 171;
        ELSIF x =- 5086 THEN
            exp_f := 171;
        ELSIF x =- 5085 THEN
            exp_f := 171;
        ELSIF x =- 5084 THEN
            exp_f := 171;
        ELSIF x =- 5083 THEN
            exp_f := 171;
        ELSIF x =- 5082 THEN
            exp_f := 171;
        ELSIF x =- 5081 THEN
            exp_f := 171;
        ELSIF x =- 5080 THEN
            exp_f := 171;
        ELSIF x =- 5079 THEN
            exp_f := 171;
        ELSIF x =- 5078 THEN
            exp_f := 171;
        ELSIF x =- 5077 THEN
            exp_f := 171;
        ELSIF x =- 5076 THEN
            exp_f := 171;
        ELSIF x =- 5075 THEN
            exp_f := 172;
        ELSIF x =- 5074 THEN
            exp_f := 172;
        ELSIF x =- 5073 THEN
            exp_f := 172;
        ELSIF x =- 5072 THEN
            exp_f := 172;
        ELSIF x =- 5071 THEN
            exp_f := 172;
        ELSIF x =- 5070 THEN
            exp_f := 172;
        ELSIF x =- 5069 THEN
            exp_f := 172;
        ELSIF x =- 5068 THEN
            exp_f := 172;
        ELSIF x =- 5067 THEN
            exp_f := 172;
        ELSIF x =- 5066 THEN
            exp_f := 172;
        ELSIF x =- 5065 THEN
            exp_f := 172;
        ELSIF x =- 5064 THEN
            exp_f := 172;
        ELSIF x =- 5063 THEN
            exp_f := 172;
        ELSIF x =- 5062 THEN
            exp_f := 173;
        ELSIF x =- 5061 THEN
            exp_f := 173;
        ELSIF x =- 5060 THEN
            exp_f := 173;
        ELSIF x =- 5059 THEN
            exp_f := 173;
        ELSIF x =- 5058 THEN
            exp_f := 173;
        ELSIF x =- 5057 THEN
            exp_f := 173;
        ELSIF x =- 5056 THEN
            exp_f := 173;
        ELSIF x =- 5055 THEN
            exp_f := 173;
        ELSIF x =- 5054 THEN
            exp_f := 173;
        ELSIF x =- 5053 THEN
            exp_f := 173;
        ELSIF x =- 5052 THEN
            exp_f := 173;
        ELSIF x =- 5051 THEN
            exp_f := 173;
        ELSIF x =- 5050 THEN
            exp_f := 174;
        ELSIF x =- 5049 THEN
            exp_f := 174;
        ELSIF x =- 5048 THEN
            exp_f := 174;
        ELSIF x =- 5047 THEN
            exp_f := 174;
        ELSIF x =- 5046 THEN
            exp_f := 174;
        ELSIF x =- 5045 THEN
            exp_f := 174;
        ELSIF x =- 5044 THEN
            exp_f := 174;
        ELSIF x =- 5043 THEN
            exp_f := 174;
        ELSIF x =- 5042 THEN
            exp_f := 174;
        ELSIF x =- 5041 THEN
            exp_f := 174;
        ELSIF x =- 5040 THEN
            exp_f := 174;
        ELSIF x =- 5039 THEN
            exp_f := 174;
        ELSIF x =- 5038 THEN
            exp_f := 174;
        ELSIF x =- 5037 THEN
            exp_f := 175;
        ELSIF x =- 5036 THEN
            exp_f := 175;
        ELSIF x =- 5035 THEN
            exp_f := 175;
        ELSIF x =- 5034 THEN
            exp_f := 175;
        ELSIF x =- 5033 THEN
            exp_f := 175;
        ELSIF x =- 5032 THEN
            exp_f := 175;
        ELSIF x =- 5031 THEN
            exp_f := 175;
        ELSIF x =- 5030 THEN
            exp_f := 175;
        ELSIF x =- 5029 THEN
            exp_f := 175;
        ELSIF x =- 5028 THEN
            exp_f := 175;
        ELSIF x =- 5027 THEN
            exp_f := 175;
        ELSIF x =- 5026 THEN
            exp_f := 175;
        ELSIF x =- 5025 THEN
            exp_f := 175;
        ELSIF x =- 5024 THEN
            exp_f := 177;
        ELSIF x =- 5023 THEN
            exp_f := 177;
        ELSIF x =- 5022 THEN
            exp_f := 177;
        ELSIF x =- 5021 THEN
            exp_f := 177;
        ELSIF x =- 5020 THEN
            exp_f := 177;
        ELSIF x =- 5019 THEN
            exp_f := 177;
        ELSIF x =- 5018 THEN
            exp_f := 177;
        ELSIF x =- 5017 THEN
            exp_f := 177;
        ELSIF x =- 5016 THEN
            exp_f := 177;
        ELSIF x =- 5015 THEN
            exp_f := 177;
        ELSIF x =- 5014 THEN
            exp_f := 177;
        ELSIF x =- 5013 THEN
            exp_f := 177;
        ELSIF x =- 5012 THEN
            exp_f := 177;
        ELSIF x =- 5011 THEN
            exp_f := 178;
        ELSIF x =- 5010 THEN
            exp_f := 178;
        ELSIF x =- 5009 THEN
            exp_f := 178;
        ELSIF x =- 5008 THEN
            exp_f := 178;
        ELSIF x =- 5007 THEN
            exp_f := 178;
        ELSIF x =- 5006 THEN
            exp_f := 178;
        ELSIF x =- 5005 THEN
            exp_f := 178;
        ELSIF x =- 5004 THEN
            exp_f := 178;
        ELSIF x =- 5003 THEN
            exp_f := 178;
        ELSIF x =- 5002 THEN
            exp_f := 178;
        ELSIF x =- 5001 THEN
            exp_f := 178;
        ELSIF x =- 5000 THEN
            exp_f := 178;
        ELSIF x =- 4999 THEN
            exp_f := 179;
        ELSIF x =- 4998 THEN
            exp_f := 179;
        ELSIF x =- 4997 THEN
            exp_f := 179;
        ELSIF x =- 4996 THEN
            exp_f := 179;
        ELSIF x =- 4995 THEN
            exp_f := 179;
        ELSIF x =- 4994 THEN
            exp_f := 179;
        ELSIF x =- 4993 THEN
            exp_f := 179;
        ELSIF x =- 4992 THEN
            exp_f := 179;
        ELSIF x =- 4991 THEN
            exp_f := 179;
        ELSIF x =- 4990 THEN
            exp_f := 179;
        ELSIF x =- 4989 THEN
            exp_f := 179;
        ELSIF x =- 4988 THEN
            exp_f := 179;
        ELSIF x =- 4987 THEN
            exp_f := 179;
        ELSIF x =- 4986 THEN
            exp_f := 180;
        ELSIF x =- 4985 THEN
            exp_f := 180;
        ELSIF x =- 4984 THEN
            exp_f := 180;
        ELSIF x =- 4983 THEN
            exp_f := 180;
        ELSIF x =- 4982 THEN
            exp_f := 180;
        ELSIF x =- 4981 THEN
            exp_f := 180;
        ELSIF x =- 4980 THEN
            exp_f := 180;
        ELSIF x =- 4979 THEN
            exp_f := 180;
        ELSIF x =- 4978 THEN
            exp_f := 180;
        ELSIF x =- 4977 THEN
            exp_f := 180;
        ELSIF x =- 4976 THEN
            exp_f := 180;
        ELSIF x =- 4975 THEN
            exp_f := 180;
        ELSIF x =- 4974 THEN
            exp_f := 180;
        ELSIF x =- 4973 THEN
            exp_f := 181;
        ELSIF x =- 4972 THEN
            exp_f := 181;
        ELSIF x =- 4971 THEN
            exp_f := 181;
        ELSIF x =- 4970 THEN
            exp_f := 181;
        ELSIF x =- 4969 THEN
            exp_f := 181;
        ELSIF x =- 4968 THEN
            exp_f := 181;
        ELSIF x =- 4967 THEN
            exp_f := 181;
        ELSIF x =- 4966 THEN
            exp_f := 181;
        ELSIF x =- 4965 THEN
            exp_f := 181;
        ELSIF x =- 4964 THEN
            exp_f := 181;
        ELSIF x =- 4963 THEN
            exp_f := 181;
        ELSIF x =- 4962 THEN
            exp_f := 181;
        ELSIF x =- 4961 THEN
            exp_f := 181;
        ELSIF x =- 4960 THEN
            exp_f := 183;
        ELSIF x =- 4959 THEN
            exp_f := 183;
        ELSIF x =- 4958 THEN
            exp_f := 183;
        ELSIF x =- 4957 THEN
            exp_f := 183;
        ELSIF x =- 4956 THEN
            exp_f := 183;
        ELSIF x =- 4955 THEN
            exp_f := 183;
        ELSIF x =- 4954 THEN
            exp_f := 183;
        ELSIF x =- 4953 THEN
            exp_f := 183;
        ELSIF x =- 4952 THEN
            exp_f := 183;
        ELSIF x =- 4951 THEN
            exp_f := 183;
        ELSIF x =- 4950 THEN
            exp_f := 183;
        ELSIF x =- 4949 THEN
            exp_f := 183;
        ELSIF x =- 4948 THEN
            exp_f := 184;
        ELSIF x =- 4947 THEN
            exp_f := 184;
        ELSIF x =- 4946 THEN
            exp_f := 184;
        ELSIF x =- 4945 THEN
            exp_f := 184;
        ELSIF x =- 4944 THEN
            exp_f := 184;
        ELSIF x =- 4943 THEN
            exp_f := 184;
        ELSIF x =- 4942 THEN
            exp_f := 184;
        ELSIF x =- 4941 THEN
            exp_f := 184;
        ELSIF x =- 4940 THEN
            exp_f := 184;
        ELSIF x =- 4939 THEN
            exp_f := 184;
        ELSIF x =- 4938 THEN
            exp_f := 184;
        ELSIF x =- 4937 THEN
            exp_f := 184;
        ELSIF x =- 4936 THEN
            exp_f := 184;
        ELSIF x =- 4935 THEN
            exp_f := 185;
        ELSIF x =- 4934 THEN
            exp_f := 185;
        ELSIF x =- 4933 THEN
            exp_f := 185;
        ELSIF x =- 4932 THEN
            exp_f := 185;
        ELSIF x =- 4931 THEN
            exp_f := 185;
        ELSIF x =- 4930 THEN
            exp_f := 185;
        ELSIF x =- 4929 THEN
            exp_f := 185;
        ELSIF x =- 4928 THEN
            exp_f := 185;
        ELSIF x =- 4927 THEN
            exp_f := 185;
        ELSIF x =- 4926 THEN
            exp_f := 185;
        ELSIF x =- 4925 THEN
            exp_f := 185;
        ELSIF x =- 4924 THEN
            exp_f := 185;
        ELSIF x =- 4923 THEN
            exp_f := 185;
        ELSIF x =- 4922 THEN
            exp_f := 186;
        ELSIF x =- 4921 THEN
            exp_f := 186;
        ELSIF x =- 4920 THEN
            exp_f := 186;
        ELSIF x =- 4919 THEN
            exp_f := 186;
        ELSIF x =- 4918 THEN
            exp_f := 186;
        ELSIF x =- 4917 THEN
            exp_f := 186;
        ELSIF x =- 4916 THEN
            exp_f := 186;
        ELSIF x =- 4915 THEN
            exp_f := 186;
        ELSIF x =- 4914 THEN
            exp_f := 186;
        ELSIF x =- 4913 THEN
            exp_f := 186;
        ELSIF x =- 4912 THEN
            exp_f := 186;
        ELSIF x =- 4911 THEN
            exp_f := 186;
        ELSIF x =- 4910 THEN
            exp_f := 187;
        ELSIF x =- 4909 THEN
            exp_f := 187;
        ELSIF x =- 4908 THEN
            exp_f := 187;
        ELSIF x =- 4907 THEN
            exp_f := 187;
        ELSIF x =- 4906 THEN
            exp_f := 187;
        ELSIF x =- 4905 THEN
            exp_f := 187;
        ELSIF x =- 4904 THEN
            exp_f := 187;
        ELSIF x =- 4903 THEN
            exp_f := 187;
        ELSIF x =- 4902 THEN
            exp_f := 187;
        ELSIF x =- 4901 THEN
            exp_f := 187;
        ELSIF x =- 4900 THEN
            exp_f := 187;
        ELSIF x =- 4899 THEN
            exp_f := 187;
        ELSIF x =- 4898 THEN
            exp_f := 187;
        ELSIF x =- 4897 THEN
            exp_f := 188;
        ELSIF x =- 4896 THEN
            exp_f := 188;
        ELSIF x =- 4895 THEN
            exp_f := 188;
        ELSIF x =- 4894 THEN
            exp_f := 188;
        ELSIF x =- 4893 THEN
            exp_f := 188;
        ELSIF x =- 4892 THEN
            exp_f := 188;
        ELSIF x =- 4891 THEN
            exp_f := 188;
        ELSIF x =- 4890 THEN
            exp_f := 188;
        ELSIF x =- 4889 THEN
            exp_f := 188;
        ELSIF x =- 4888 THEN
            exp_f := 188;
        ELSIF x =- 4887 THEN
            exp_f := 188;
        ELSIF x =- 4886 THEN
            exp_f := 188;
        ELSIF x =- 4885 THEN
            exp_f := 188;
        ELSIF x =- 4884 THEN
            exp_f := 190;
        ELSIF x =- 4883 THEN
            exp_f := 190;
        ELSIF x =- 4882 THEN
            exp_f := 190;
        ELSIF x =- 4881 THEN
            exp_f := 190;
        ELSIF x =- 4880 THEN
            exp_f := 190;
        ELSIF x =- 4879 THEN
            exp_f := 190;
        ELSIF x =- 4878 THEN
            exp_f := 190;
        ELSIF x =- 4877 THEN
            exp_f := 190;
        ELSIF x =- 4876 THEN
            exp_f := 190;
        ELSIF x =- 4875 THEN
            exp_f := 190;
        ELSIF x =- 4874 THEN
            exp_f := 190;
        ELSIF x =- 4873 THEN
            exp_f := 190;
        ELSIF x =- 4872 THEN
            exp_f := 190;
        ELSIF x =- 4871 THEN
            exp_f := 191;
        ELSIF x =- 4870 THEN
            exp_f := 191;
        ELSIF x =- 4869 THEN
            exp_f := 191;
        ELSIF x =- 4868 THEN
            exp_f := 191;
        ELSIF x =- 4867 THEN
            exp_f := 191;
        ELSIF x =- 4866 THEN
            exp_f := 191;
        ELSIF x =- 4865 THEN
            exp_f := 191;
        ELSIF x =- 4864 THEN
            exp_f := 191;
        ELSIF x =- 4863 THEN
            exp_f := 191;
        ELSIF x =- 4862 THEN
            exp_f := 191;
        ELSIF x =- 4861 THEN
            exp_f := 191;
        ELSIF x =- 4860 THEN
            exp_f := 191;
        ELSIF x =- 4859 THEN
            exp_f := 192;
        ELSIF x =- 4858 THEN
            exp_f := 192;
        ELSIF x =- 4857 THEN
            exp_f := 192;
        ELSIF x =- 4856 THEN
            exp_f := 192;
        ELSIF x =- 4855 THEN
            exp_f := 192;
        ELSIF x =- 4854 THEN
            exp_f := 192;
        ELSIF x =- 4853 THEN
            exp_f := 192;
        ELSIF x =- 4852 THEN
            exp_f := 192;
        ELSIF x =- 4851 THEN
            exp_f := 192;
        ELSIF x =- 4850 THEN
            exp_f := 192;
        ELSIF x =- 4849 THEN
            exp_f := 192;
        ELSIF x =- 4848 THEN
            exp_f := 192;
        ELSIF x =- 4847 THEN
            exp_f := 192;
        ELSIF x =- 4846 THEN
            exp_f := 193;
        ELSIF x =- 4845 THEN
            exp_f := 193;
        ELSIF x =- 4844 THEN
            exp_f := 193;
        ELSIF x =- 4843 THEN
            exp_f := 193;
        ELSIF x =- 4842 THEN
            exp_f := 193;
        ELSIF x =- 4841 THEN
            exp_f := 193;
        ELSIF x =- 4840 THEN
            exp_f := 193;
        ELSIF x =- 4839 THEN
            exp_f := 193;
        ELSIF x =- 4838 THEN
            exp_f := 193;
        ELSIF x =- 4837 THEN
            exp_f := 193;
        ELSIF x =- 4836 THEN
            exp_f := 193;
        ELSIF x =- 4835 THEN
            exp_f := 193;
        ELSIF x =- 4834 THEN
            exp_f := 193;
        ELSIF x =- 4833 THEN
            exp_f := 194;
        ELSIF x =- 4832 THEN
            exp_f := 194;
        ELSIF x =- 4831 THEN
            exp_f := 194;
        ELSIF x =- 4830 THEN
            exp_f := 194;
        ELSIF x =- 4829 THEN
            exp_f := 194;
        ELSIF x =- 4828 THEN
            exp_f := 194;
        ELSIF x =- 4827 THEN
            exp_f := 194;
        ELSIF x =- 4826 THEN
            exp_f := 194;
        ELSIF x =- 4825 THEN
            exp_f := 194;
        ELSIF x =- 4824 THEN
            exp_f := 194;
        ELSIF x =- 4823 THEN
            exp_f := 194;
        ELSIF x =- 4822 THEN
            exp_f := 194;
        ELSIF x =- 4821 THEN
            exp_f := 196;
        ELSIF x =- 4820 THEN
            exp_f := 196;
        ELSIF x =- 4819 THEN
            exp_f := 196;
        ELSIF x =- 4818 THEN
            exp_f := 196;
        ELSIF x =- 4817 THEN
            exp_f := 196;
        ELSIF x =- 4816 THEN
            exp_f := 196;
        ELSIF x =- 4815 THEN
            exp_f := 196;
        ELSIF x =- 4814 THEN
            exp_f := 196;
        ELSIF x =- 4813 THEN
            exp_f := 196;
        ELSIF x =- 4812 THEN
            exp_f := 196;
        ELSIF x =- 4811 THEN
            exp_f := 196;
        ELSIF x =- 4810 THEN
            exp_f := 196;
        ELSIF x =- 4809 THEN
            exp_f := 196;
        ELSIF x =- 4808 THEN
            exp_f := 197;
        ELSIF x =- 4807 THEN
            exp_f := 197;
        ELSIF x =- 4806 THEN
            exp_f := 197;
        ELSIF x =- 4805 THEN
            exp_f := 197;
        ELSIF x =- 4804 THEN
            exp_f := 197;
        ELSIF x =- 4803 THEN
            exp_f := 197;
        ELSIF x =- 4802 THEN
            exp_f := 197;
        ELSIF x =- 4801 THEN
            exp_f := 197;
        ELSIF x =- 4800 THEN
            exp_f := 197;
        ELSIF x =- 4799 THEN
            exp_f := 197;
        ELSIF x =- 4798 THEN
            exp_f := 197;
        ELSIF x =- 4797 THEN
            exp_f := 197;
        ELSIF x =- 4796 THEN
            exp_f := 197;
        ELSIF x =- 4795 THEN
            exp_f := 198;
        ELSIF x =- 4794 THEN
            exp_f := 198;
        ELSIF x =- 4793 THEN
            exp_f := 198;
        ELSIF x =- 4792 THEN
            exp_f := 198;
        ELSIF x =- 4791 THEN
            exp_f := 198;
        ELSIF x =- 4790 THEN
            exp_f := 198;
        ELSIF x =- 4789 THEN
            exp_f := 198;
        ELSIF x =- 4788 THEN
            exp_f := 198;
        ELSIF x =- 4787 THEN
            exp_f := 198;
        ELSIF x =- 4786 THEN
            exp_f := 198;
        ELSIF x =- 4785 THEN
            exp_f := 198;
        ELSIF x =- 4784 THEN
            exp_f := 198;
        ELSIF x =- 4783 THEN
            exp_f := 198;
        ELSIF x =- 4782 THEN
            exp_f := 199;
        ELSIF x =- 4781 THEN
            exp_f := 199;
        ELSIF x =- 4780 THEN
            exp_f := 199;
        ELSIF x =- 4779 THEN
            exp_f := 199;
        ELSIF x =- 4778 THEN
            exp_f := 199;
        ELSIF x =- 4777 THEN
            exp_f := 199;
        ELSIF x =- 4776 THEN
            exp_f := 199;
        ELSIF x =- 4775 THEN
            exp_f := 199;
        ELSIF x =- 4774 THEN
            exp_f := 199;
        ELSIF x =- 4773 THEN
            exp_f := 199;
        ELSIF x =- 4772 THEN
            exp_f := 199;
        ELSIF x =- 4771 THEN
            exp_f := 199;
        ELSIF x =- 4770 THEN
            exp_f := 200;
        ELSIF x =- 4769 THEN
            exp_f := 200;
        ELSIF x =- 4768 THEN
            exp_f := 200;
        ELSIF x =- 4767 THEN
            exp_f := 200;
        ELSIF x =- 4766 THEN
            exp_f := 200;
        ELSIF x =- 4765 THEN
            exp_f := 200;
        ELSIF x =- 4764 THEN
            exp_f := 200;
        ELSIF x =- 4763 THEN
            exp_f := 200;
        ELSIF x =- 4762 THEN
            exp_f := 200;
        ELSIF x =- 4761 THEN
            exp_f := 200;
        ELSIF x =- 4760 THEN
            exp_f := 200;
        ELSIF x =- 4759 THEN
            exp_f := 200;
        ELSIF x =- 4758 THEN
            exp_f := 200;
        ELSIF x =- 4757 THEN
            exp_f := 202;
        ELSIF x =- 4756 THEN
            exp_f := 202;
        ELSIF x =- 4755 THEN
            exp_f := 202;
        ELSIF x =- 4754 THEN
            exp_f := 202;
        ELSIF x =- 4753 THEN
            exp_f := 202;
        ELSIF x =- 4752 THEN
            exp_f := 202;
        ELSIF x =- 4751 THEN
            exp_f := 202;
        ELSIF x =- 4750 THEN
            exp_f := 202;
        ELSIF x =- 4749 THEN
            exp_f := 202;
        ELSIF x =- 4748 THEN
            exp_f := 202;
        ELSIF x =- 4747 THEN
            exp_f := 202;
        ELSIF x =- 4746 THEN
            exp_f := 202;
        ELSIF x =- 4745 THEN
            exp_f := 202;
        ELSIF x =- 4744 THEN
            exp_f := 203;
        ELSIF x =- 4743 THEN
            exp_f := 203;
        ELSIF x =- 4742 THEN
            exp_f := 203;
        ELSIF x =- 4741 THEN
            exp_f := 203;
        ELSIF x =- 4740 THEN
            exp_f := 203;
        ELSIF x =- 4739 THEN
            exp_f := 203;
        ELSIF x =- 4738 THEN
            exp_f := 203;
        ELSIF x =- 4737 THEN
            exp_f := 203;
        ELSIF x =- 4736 THEN
            exp_f := 203;
        ELSIF x =- 4735 THEN
            exp_f := 203;
        ELSIF x =- 4734 THEN
            exp_f := 203;
        ELSIF x =- 4733 THEN
            exp_f := 203;
        ELSIF x =- 4732 THEN
            exp_f := 204;
        ELSIF x =- 4731 THEN
            exp_f := 204;
        ELSIF x =- 4730 THEN
            exp_f := 204;
        ELSIF x =- 4729 THEN
            exp_f := 204;
        ELSIF x =- 4728 THEN
            exp_f := 204;
        ELSIF x =- 4727 THEN
            exp_f := 204;
        ELSIF x =- 4726 THEN
            exp_f := 204;
        ELSIF x =- 4725 THEN
            exp_f := 204;
        ELSIF x =- 4724 THEN
            exp_f := 204;
        ELSIF x =- 4723 THEN
            exp_f := 204;
        ELSIF x =- 4722 THEN
            exp_f := 204;
        ELSIF x =- 4721 THEN
            exp_f := 204;
        ELSIF x =- 4720 THEN
            exp_f := 204;
        ELSIF x =- 4719 THEN
            exp_f := 205;
        ELSIF x =- 4718 THEN
            exp_f := 205;
        ELSIF x =- 4717 THEN
            exp_f := 205;
        ELSIF x =- 4716 THEN
            exp_f := 205;
        ELSIF x =- 4715 THEN
            exp_f := 205;
        ELSIF x =- 4714 THEN
            exp_f := 205;
        ELSIF x =- 4713 THEN
            exp_f := 205;
        ELSIF x =- 4712 THEN
            exp_f := 205;
        ELSIF x =- 4711 THEN
            exp_f := 205;
        ELSIF x =- 4710 THEN
            exp_f := 205;
        ELSIF x =- 4709 THEN
            exp_f := 205;
        ELSIF x =- 4708 THEN
            exp_f := 205;
        ELSIF x =- 4707 THEN
            exp_f := 205;
        ELSIF x =- 4706 THEN
            exp_f := 207;
        ELSIF x =- 4705 THEN
            exp_f := 207;
        ELSIF x =- 4704 THEN
            exp_f := 207;
        ELSIF x =- 4703 THEN
            exp_f := 207;
        ELSIF x =- 4702 THEN
            exp_f := 207;
        ELSIF x =- 4701 THEN
            exp_f := 207;
        ELSIF x =- 4700 THEN
            exp_f := 207;
        ELSIF x =- 4699 THEN
            exp_f := 207;
        ELSIF x =- 4698 THEN
            exp_f := 207;
        ELSIF x =- 4697 THEN
            exp_f := 207;
        ELSIF x =- 4696 THEN
            exp_f := 207;
        ELSIF x =- 4695 THEN
            exp_f := 207;
        ELSIF x =- 4694 THEN
            exp_f := 207;
        ELSIF x =- 4693 THEN
            exp_f := 208;
        ELSIF x =- 4692 THEN
            exp_f := 208;
        ELSIF x =- 4691 THEN
            exp_f := 208;
        ELSIF x =- 4690 THEN
            exp_f := 208;
        ELSIF x =- 4689 THEN
            exp_f := 208;
        ELSIF x =- 4688 THEN
            exp_f := 208;
        ELSIF x =- 4687 THEN
            exp_f := 208;
        ELSIF x =- 4686 THEN
            exp_f := 208;
        ELSIF x =- 4685 THEN
            exp_f := 208;
        ELSIF x =- 4684 THEN
            exp_f := 208;
        ELSIF x =- 4683 THEN
            exp_f := 208;
        ELSIF x =- 4682 THEN
            exp_f := 208;
        ELSIF x =- 4681 THEN
            exp_f := 209;
        ELSIF x =- 4680 THEN
            exp_f := 209;
        ELSIF x =- 4679 THEN
            exp_f := 209;
        ELSIF x =- 4678 THEN
            exp_f := 209;
        ELSIF x =- 4677 THEN
            exp_f := 209;
        ELSIF x =- 4676 THEN
            exp_f := 209;
        ELSIF x =- 4675 THEN
            exp_f := 209;
        ELSIF x =- 4674 THEN
            exp_f := 209;
        ELSIF x =- 4673 THEN
            exp_f := 209;
        ELSIF x =- 4672 THEN
            exp_f := 209;
        ELSIF x =- 4671 THEN
            exp_f := 209;
        ELSIF x =- 4670 THEN
            exp_f := 209;
        ELSIF x =- 4669 THEN
            exp_f := 209;
        ELSIF x =- 4668 THEN
            exp_f := 210;
        ELSIF x =- 4667 THEN
            exp_f := 210;
        ELSIF x =- 4666 THEN
            exp_f := 210;
        ELSIF x =- 4665 THEN
            exp_f := 210;
        ELSIF x =- 4664 THEN
            exp_f := 210;
        ELSIF x =- 4663 THEN
            exp_f := 210;
        ELSIF x =- 4662 THEN
            exp_f := 210;
        ELSIF x =- 4661 THEN
            exp_f := 210;
        ELSIF x =- 4660 THEN
            exp_f := 210;
        ELSIF x =- 4659 THEN
            exp_f := 210;
        ELSIF x =- 4658 THEN
            exp_f := 210;
        ELSIF x =- 4657 THEN
            exp_f := 210;
        ELSIF x =- 4656 THEN
            exp_f := 210;
        ELSIF x =- 4655 THEN
            exp_f := 211;
        ELSIF x =- 4654 THEN
            exp_f := 211;
        ELSIF x =- 4653 THEN
            exp_f := 211;
        ELSIF x =- 4652 THEN
            exp_f := 211;
        ELSIF x =- 4651 THEN
            exp_f := 211;
        ELSIF x =- 4650 THEN
            exp_f := 211;
        ELSIF x =- 4649 THEN
            exp_f := 211;
        ELSIF x =- 4648 THEN
            exp_f := 211;
        ELSIF x =- 4647 THEN
            exp_f := 211;
        ELSIF x =- 4646 THEN
            exp_f := 211;
        ELSIF x =- 4645 THEN
            exp_f := 211;
        ELSIF x =- 4644 THEN
            exp_f := 211;
        ELSIF x =- 4643 THEN
            exp_f := 211;
        ELSIF x =- 4642 THEN
            exp_f := 213;
        ELSIF x =- 4641 THEN
            exp_f := 213;
        ELSIF x =- 4640 THEN
            exp_f := 213;
        ELSIF x =- 4639 THEN
            exp_f := 213;
        ELSIF x =- 4638 THEN
            exp_f := 213;
        ELSIF x =- 4637 THEN
            exp_f := 213;
        ELSIF x =- 4636 THEN
            exp_f := 213;
        ELSIF x =- 4635 THEN
            exp_f := 213;
        ELSIF x =- 4634 THEN
            exp_f := 213;
        ELSIF x =- 4633 THEN
            exp_f := 213;
        ELSIF x =- 4632 THEN
            exp_f := 213;
        ELSIF x =- 4631 THEN
            exp_f := 213;
        ELSIF x =- 4630 THEN
            exp_f := 214;
        ELSIF x =- 4629 THEN
            exp_f := 214;
        ELSIF x =- 4628 THEN
            exp_f := 214;
        ELSIF x =- 4627 THEN
            exp_f := 214;
        ELSIF x =- 4626 THEN
            exp_f := 214;
        ELSIF x =- 4625 THEN
            exp_f := 214;
        ELSIF x =- 4624 THEN
            exp_f := 214;
        ELSIF x =- 4623 THEN
            exp_f := 214;
        ELSIF x =- 4622 THEN
            exp_f := 214;
        ELSIF x =- 4621 THEN
            exp_f := 214;
        ELSIF x =- 4620 THEN
            exp_f := 214;
        ELSIF x =- 4619 THEN
            exp_f := 214;
        ELSIF x =- 4618 THEN
            exp_f := 214;
        ELSIF x =- 4617 THEN
            exp_f := 215;
        ELSIF x =- 4616 THEN
            exp_f := 215;
        ELSIF x =- 4615 THEN
            exp_f := 215;
        ELSIF x =- 4614 THEN
            exp_f := 215;
        ELSIF x =- 4613 THEN
            exp_f := 215;
        ELSIF x =- 4612 THEN
            exp_f := 215;
        ELSIF x =- 4611 THEN
            exp_f := 215;
        ELSIF x =- 4610 THEN
            exp_f := 215;
        ELSIF x =- 4609 THEN
            exp_f := 215;
        ELSIF x =- 4608 THEN
            exp_f := 215;
        ELSIF x =- 4607 THEN
            exp_f := 215;
        ELSIF x =- 4606 THEN
            exp_f := 215;
        ELSIF x =- 4605 THEN
            exp_f := 216;
        ELSIF x =- 4604 THEN
            exp_f := 216;
        ELSIF x =- 4603 THEN
            exp_f := 216;
        ELSIF x =- 4602 THEN
            exp_f := 216;
        ELSIF x =- 4601 THEN
            exp_f := 216;
        ELSIF x =- 4600 THEN
            exp_f := 216;
        ELSIF x =- 4599 THEN
            exp_f := 216;
        ELSIF x =- 4598 THEN
            exp_f := 216;
        ELSIF x =- 4597 THEN
            exp_f := 216;
        ELSIF x =- 4596 THEN
            exp_f := 216;
        ELSIF x =- 4595 THEN
            exp_f := 216;
        ELSIF x =- 4594 THEN
            exp_f := 217;
        ELSIF x =- 4593 THEN
            exp_f := 217;
        ELSIF x =- 4592 THEN
            exp_f := 217;
        ELSIF x =- 4591 THEN
            exp_f := 217;
        ELSIF x =- 4590 THEN
            exp_f := 217;
        ELSIF x =- 4589 THEN
            exp_f := 217;
        ELSIF x =- 4588 THEN
            exp_f := 217;
        ELSIF x =- 4587 THEN
            exp_f := 217;
        ELSIF x =- 4586 THEN
            exp_f := 217;
        ELSIF x =- 4585 THEN
            exp_f := 217;
        ELSIF x =- 4584 THEN
            exp_f := 219;
        ELSIF x =- 4583 THEN
            exp_f := 219;
        ELSIF x =- 4582 THEN
            exp_f := 219;
        ELSIF x =- 4581 THEN
            exp_f := 219;
        ELSIF x =- 4580 THEN
            exp_f := 219;
        ELSIF x =- 4579 THEN
            exp_f := 219;
        ELSIF x =- 4578 THEN
            exp_f := 219;
        ELSIF x =- 4577 THEN
            exp_f := 219;
        ELSIF x =- 4576 THEN
            exp_f := 219;
        ELSIF x =- 4575 THEN
            exp_f := 219;
        ELSIF x =- 4574 THEN
            exp_f := 219;
        ELSIF x =- 4573 THEN
            exp_f := 220;
        ELSIF x =- 4572 THEN
            exp_f := 220;
        ELSIF x =- 4571 THEN
            exp_f := 220;
        ELSIF x =- 4570 THEN
            exp_f := 220;
        ELSIF x =- 4569 THEN
            exp_f := 220;
        ELSIF x =- 4568 THEN
            exp_f := 220;
        ELSIF x =- 4567 THEN
            exp_f := 220;
        ELSIF x =- 4566 THEN
            exp_f := 220;
        ELSIF x =- 4565 THEN
            exp_f := 220;
        ELSIF x =- 4564 THEN
            exp_f := 220;
        ELSIF x =- 4563 THEN
            exp_f := 220;
        ELSIF x =- 4562 THEN
            exp_f := 221;
        ELSIF x =- 4561 THEN
            exp_f := 221;
        ELSIF x =- 4560 THEN
            exp_f := 221;
        ELSIF x =- 4559 THEN
            exp_f := 221;
        ELSIF x =- 4558 THEN
            exp_f := 221;
        ELSIF x =- 4557 THEN
            exp_f := 221;
        ELSIF x =- 4556 THEN
            exp_f := 221;
        ELSIF x =- 4555 THEN
            exp_f := 221;
        ELSIF x =- 4554 THEN
            exp_f := 221;
        ELSIF x =- 4553 THEN
            exp_f := 221;
        ELSIF x =- 4552 THEN
            exp_f := 222;
        ELSIF x =- 4551 THEN
            exp_f := 222;
        ELSIF x =- 4550 THEN
            exp_f := 222;
        ELSIF x =- 4549 THEN
            exp_f := 222;
        ELSIF x =- 4548 THEN
            exp_f := 222;
        ELSIF x =- 4547 THEN
            exp_f := 222;
        ELSIF x =- 4546 THEN
            exp_f := 222;
        ELSIF x =- 4545 THEN
            exp_f := 222;
        ELSIF x =- 4544 THEN
            exp_f := 222;
        ELSIF x =- 4543 THEN
            exp_f := 222;
        ELSIF x =- 4542 THEN
            exp_f := 222;
        ELSIF x =- 4541 THEN
            exp_f := 224;
        ELSIF x =- 4540 THEN
            exp_f := 224;
        ELSIF x =- 4539 THEN
            exp_f := 224;
        ELSIF x =- 4538 THEN
            exp_f := 224;
        ELSIF x =- 4537 THEN
            exp_f := 224;
        ELSIF x =- 4536 THEN
            exp_f := 224;
        ELSIF x =- 4535 THEN
            exp_f := 224;
        ELSIF x =- 4534 THEN
            exp_f := 224;
        ELSIF x =- 4533 THEN
            exp_f := 224;
        ELSIF x =- 4532 THEN
            exp_f := 224;
        ELSIF x =- 4531 THEN
            exp_f := 225;
        ELSIF x =- 4530 THEN
            exp_f := 225;
        ELSIF x =- 4529 THEN
            exp_f := 225;
        ELSIF x =- 4528 THEN
            exp_f := 225;
        ELSIF x =- 4527 THEN
            exp_f := 225;
        ELSIF x =- 4526 THEN
            exp_f := 225;
        ELSIF x =- 4525 THEN
            exp_f := 225;
        ELSIF x =- 4524 THEN
            exp_f := 225;
        ELSIF x =- 4523 THEN
            exp_f := 225;
        ELSIF x =- 4522 THEN
            exp_f := 225;
        ELSIF x =- 4521 THEN
            exp_f := 225;
        ELSIF x =- 4520 THEN
            exp_f := 226;
        ELSIF x =- 4519 THEN
            exp_f := 226;
        ELSIF x =- 4518 THEN
            exp_f := 226;
        ELSIF x =- 4517 THEN
            exp_f := 226;
        ELSIF x =- 4516 THEN
            exp_f := 226;
        ELSIF x =- 4515 THEN
            exp_f := 226;
        ELSIF x =- 4514 THEN
            exp_f := 226;
        ELSIF x =- 4513 THEN
            exp_f := 226;
        ELSIF x =- 4512 THEN
            exp_f := 226;
        ELSIF x =- 4511 THEN
            exp_f := 226;
        ELSIF x =- 4510 THEN
            exp_f := 226;
        ELSIF x =- 4509 THEN
            exp_f := 227;
        ELSIF x =- 4508 THEN
            exp_f := 227;
        ELSIF x =- 4507 THEN
            exp_f := 227;
        ELSIF x =- 4506 THEN
            exp_f := 227;
        ELSIF x =- 4505 THEN
            exp_f := 227;
        ELSIF x =- 4504 THEN
            exp_f := 227;
        ELSIF x =- 4503 THEN
            exp_f := 227;
        ELSIF x =- 4502 THEN
            exp_f := 227;
        ELSIF x =- 4501 THEN
            exp_f := 227;
        ELSIF x =- 4500 THEN
            exp_f := 227;
        ELSIF x =- 4499 THEN
            exp_f := 229;
        ELSIF x =- 4498 THEN
            exp_f := 229;
        ELSIF x =- 4497 THEN
            exp_f := 229;
        ELSIF x =- 4496 THEN
            exp_f := 229;
        ELSIF x =- 4495 THEN
            exp_f := 229;
        ELSIF x =- 4494 THEN
            exp_f := 229;
        ELSIF x =- 4493 THEN
            exp_f := 229;
        ELSIF x =- 4492 THEN
            exp_f := 229;
        ELSIF x =- 4491 THEN
            exp_f := 229;
        ELSIF x =- 4490 THEN
            exp_f := 229;
        ELSIF x =- 4489 THEN
            exp_f := 229;
        ELSIF x =- 4488 THEN
            exp_f := 230;
        ELSIF x =- 4487 THEN
            exp_f := 230;
        ELSIF x =- 4486 THEN
            exp_f := 230;
        ELSIF x =- 4485 THEN
            exp_f := 230;
        ELSIF x =- 4484 THEN
            exp_f := 230;
        ELSIF x =- 4483 THEN
            exp_f := 230;
        ELSIF x =- 4482 THEN
            exp_f := 230;
        ELSIF x =- 4481 THEN
            exp_f := 230;
        ELSIF x =- 4480 THEN
            exp_f := 230;
        ELSIF x =- 4479 THEN
            exp_f := 230;
        ELSIF x =- 4478 THEN
            exp_f := 231;
        ELSIF x =- 4477 THEN
            exp_f := 231;
        ELSIF x =- 4476 THEN
            exp_f := 231;
        ELSIF x =- 4475 THEN
            exp_f := 231;
        ELSIF x =- 4474 THEN
            exp_f := 231;
        ELSIF x =- 4473 THEN
            exp_f := 231;
        ELSIF x =- 4472 THEN
            exp_f := 231;
        ELSIF x =- 4471 THEN
            exp_f := 231;
        ELSIF x =- 4470 THEN
            exp_f := 231;
        ELSIF x =- 4469 THEN
            exp_f := 231;
        ELSIF x =- 4468 THEN
            exp_f := 231;
        ELSIF x =- 4467 THEN
            exp_f := 232;
        ELSIF x =- 4466 THEN
            exp_f := 232;
        ELSIF x =- 4465 THEN
            exp_f := 232;
        ELSIF x =- 4464 THEN
            exp_f := 232;
        ELSIF x =- 4463 THEN
            exp_f := 232;
        ELSIF x =- 4462 THEN
            exp_f := 232;
        ELSIF x =- 4461 THEN
            exp_f := 232;
        ELSIF x =- 4460 THEN
            exp_f := 232;
        ELSIF x =- 4459 THEN
            exp_f := 232;
        ELSIF x =- 4458 THEN
            exp_f := 232;
        ELSIF x =- 4457 THEN
            exp_f := 232;
        ELSIF x =- 4456 THEN
            exp_f := 233;
        ELSIF x =- 4455 THEN
            exp_f := 233;
        ELSIF x =- 4454 THEN
            exp_f := 233;
        ELSIF x =- 4453 THEN
            exp_f := 233;
        ELSIF x =- 4452 THEN
            exp_f := 233;
        ELSIF x =- 4451 THEN
            exp_f := 233;
        ELSIF x =- 4450 THEN
            exp_f := 233;
        ELSIF x =- 4449 THEN
            exp_f := 233;
        ELSIF x =- 4448 THEN
            exp_f := 233;
        ELSIF x =- 4447 THEN
            exp_f := 233;
        ELSIF x =- 4446 THEN
            exp_f := 235;
        ELSIF x =- 4445 THEN
            exp_f := 235;
        ELSIF x =- 4444 THEN
            exp_f := 235;
        ELSIF x =- 4443 THEN
            exp_f := 235;
        ELSIF x =- 4442 THEN
            exp_f := 235;
        ELSIF x =- 4441 THEN
            exp_f := 235;
        ELSIF x =- 4440 THEN
            exp_f := 235;
        ELSIF x =- 4439 THEN
            exp_f := 235;
        ELSIF x =- 4438 THEN
            exp_f := 235;
        ELSIF x =- 4437 THEN
            exp_f := 235;
        ELSIF x =- 4436 THEN
            exp_f := 235;
        ELSIF x =- 4435 THEN
            exp_f := 236;
        ELSIF x =- 4434 THEN
            exp_f := 236;
        ELSIF x =- 4433 THEN
            exp_f := 236;
        ELSIF x =- 4432 THEN
            exp_f := 236;
        ELSIF x =- 4431 THEN
            exp_f := 236;
        ELSIF x =- 4430 THEN
            exp_f := 236;
        ELSIF x =- 4429 THEN
            exp_f := 236;
        ELSIF x =- 4428 THEN
            exp_f := 236;
        ELSIF x =- 4427 THEN
            exp_f := 236;
        ELSIF x =- 4426 THEN
            exp_f := 236;
        ELSIF x =- 4425 THEN
            exp_f := 236;
        ELSIF x =- 4424 THEN
            exp_f := 237;
        ELSIF x =- 4423 THEN
            exp_f := 237;
        ELSIF x =- 4422 THEN
            exp_f := 237;
        ELSIF x =- 4421 THEN
            exp_f := 237;
        ELSIF x =- 4420 THEN
            exp_f := 237;
        ELSIF x =- 4419 THEN
            exp_f := 237;
        ELSIF x =- 4418 THEN
            exp_f := 237;
        ELSIF x =- 4417 THEN
            exp_f := 237;
        ELSIF x =- 4416 THEN
            exp_f := 237;
        ELSIF x =- 4415 THEN
            exp_f := 237;
        ELSIF x =- 4414 THEN
            exp_f := 238;
        ELSIF x =- 4413 THEN
            exp_f := 238;
        ELSIF x =- 4412 THEN
            exp_f := 238;
        ELSIF x =- 4411 THEN
            exp_f := 238;
        ELSIF x =- 4410 THEN
            exp_f := 238;
        ELSIF x =- 4409 THEN
            exp_f := 238;
        ELSIF x =- 4408 THEN
            exp_f := 238;
        ELSIF x =- 4407 THEN
            exp_f := 238;
        ELSIF x =- 4406 THEN
            exp_f := 238;
        ELSIF x =- 4405 THEN
            exp_f := 238;
        ELSIF x =- 4404 THEN
            exp_f := 238;
        ELSIF x =- 4403 THEN
            exp_f := 240;
        ELSIF x =- 4402 THEN
            exp_f := 240;
        ELSIF x =- 4401 THEN
            exp_f := 240;
        ELSIF x =- 4400 THEN
            exp_f := 240;
        ELSIF x =- 4399 THEN
            exp_f := 240;
        ELSIF x =- 4398 THEN
            exp_f := 240;
        ELSIF x =- 4397 THEN
            exp_f := 240;
        ELSIF x =- 4396 THEN
            exp_f := 240;
        ELSIF x =- 4395 THEN
            exp_f := 240;
        ELSIF x =- 4394 THEN
            exp_f := 240;
        ELSIF x =- 4393 THEN
            exp_f := 241;
        ELSIF x =- 4392 THEN
            exp_f := 241;
        ELSIF x =- 4391 THEN
            exp_f := 241;
        ELSIF x =- 4390 THEN
            exp_f := 241;
        ELSIF x =- 4389 THEN
            exp_f := 241;
        ELSIF x =- 4388 THEN
            exp_f := 241;
        ELSIF x =- 4387 THEN
            exp_f := 241;
        ELSIF x =- 4386 THEN
            exp_f := 241;
        ELSIF x =- 4385 THEN
            exp_f := 241;
        ELSIF x =- 4384 THEN
            exp_f := 241;
        ELSIF x =- 4383 THEN
            exp_f := 241;
        ELSIF x =- 4382 THEN
            exp_f := 242;
        ELSIF x =- 4381 THEN
            exp_f := 242;
        ELSIF x =- 4380 THEN
            exp_f := 242;
        ELSIF x =- 4379 THEN
            exp_f := 242;
        ELSIF x =- 4378 THEN
            exp_f := 242;
        ELSIF x =- 4377 THEN
            exp_f := 242;
        ELSIF x =- 4376 THEN
            exp_f := 242;
        ELSIF x =- 4375 THEN
            exp_f := 242;
        ELSIF x =- 4374 THEN
            exp_f := 242;
        ELSIF x =- 4373 THEN
            exp_f := 242;
        ELSIF x =- 4372 THEN
            exp_f := 242;
        ELSIF x =- 4371 THEN
            exp_f := 243;
        ELSIF x =- 4370 THEN
            exp_f := 243;
        ELSIF x =- 4369 THEN
            exp_f := 243;
        ELSIF x =- 4368 THEN
            exp_f := 243;
        ELSIF x =- 4367 THEN
            exp_f := 243;
        ELSIF x =- 4366 THEN
            exp_f := 243;
        ELSIF x =- 4365 THEN
            exp_f := 243;
        ELSIF x =- 4364 THEN
            exp_f := 243;
        ELSIF x =- 4363 THEN
            exp_f := 243;
        ELSIF x =- 4362 THEN
            exp_f := 243;
        ELSIF x =- 4361 THEN
            exp_f := 245;
        ELSIF x =- 4360 THEN
            exp_f := 245;
        ELSIF x =- 4359 THEN
            exp_f := 245;
        ELSIF x =- 4358 THEN
            exp_f := 245;
        ELSIF x =- 4357 THEN
            exp_f := 245;
        ELSIF x =- 4356 THEN
            exp_f := 245;
        ELSIF x =- 4355 THEN
            exp_f := 245;
        ELSIF x =- 4354 THEN
            exp_f := 245;
        ELSIF x =- 4353 THEN
            exp_f := 245;
        ELSIF x =- 4352 THEN
            exp_f := 245;
        ELSIF x =- 4351 THEN
            exp_f := 245;
        ELSIF x =- 4350 THEN
            exp_f := 246;
        ELSIF x =- 4349 THEN
            exp_f := 246;
        ELSIF x =- 4348 THEN
            exp_f := 246;
        ELSIF x =- 4347 THEN
            exp_f := 246;
        ELSIF x =- 4346 THEN
            exp_f := 246;
        ELSIF x =- 4345 THEN
            exp_f := 246;
        ELSIF x =- 4344 THEN
            exp_f := 246;
        ELSIF x =- 4343 THEN
            exp_f := 246;
        ELSIF x =- 4342 THEN
            exp_f := 246;
        ELSIF x =- 4341 THEN
            exp_f := 246;
        ELSIF x =- 4340 THEN
            exp_f := 247;
        ELSIF x =- 4339 THEN
            exp_f := 247;
        ELSIF x =- 4338 THEN
            exp_f := 247;
        ELSIF x =- 4337 THEN
            exp_f := 247;
        ELSIF x =- 4336 THEN
            exp_f := 247;
        ELSIF x =- 4335 THEN
            exp_f := 247;
        ELSIF x =- 4334 THEN
            exp_f := 247;
        ELSIF x =- 4333 THEN
            exp_f := 247;
        ELSIF x =- 4332 THEN
            exp_f := 247;
        ELSIF x =- 4331 THEN
            exp_f := 247;
        ELSIF x =- 4330 THEN
            exp_f := 247;
        ELSIF x =- 4329 THEN
            exp_f := 248;
        ELSIF x =- 4328 THEN
            exp_f := 248;
        ELSIF x =- 4327 THEN
            exp_f := 248;
        ELSIF x =- 4326 THEN
            exp_f := 248;
        ELSIF x =- 4325 THEN
            exp_f := 248;
        ELSIF x =- 4324 THEN
            exp_f := 248;
        ELSIF x =- 4323 THEN
            exp_f := 248;
        ELSIF x =- 4322 THEN
            exp_f := 248;
        ELSIF x =- 4321 THEN
            exp_f := 248;
        ELSIF x =- 4320 THEN
            exp_f := 248;
        ELSIF x =- 4319 THEN
            exp_f := 248;
        ELSIF x =- 4318 THEN
            exp_f := 250;
        ELSIF x =- 4317 THEN
            exp_f := 250;
        ELSIF x =- 4316 THEN
            exp_f := 250;
        ELSIF x =- 4315 THEN
            exp_f := 250;
        ELSIF x =- 4314 THEN
            exp_f := 250;
        ELSIF x =- 4313 THEN
            exp_f := 250;
        ELSIF x =- 4312 THEN
            exp_f := 250;
        ELSIF x =- 4311 THEN
            exp_f := 250;
        ELSIF x =- 4310 THEN
            exp_f := 250;
        ELSIF x =- 4309 THEN
            exp_f := 250;
        ELSIF x =- 4308 THEN
            exp_f := 251;
        ELSIF x =- 4307 THEN
            exp_f := 251;
        ELSIF x =- 4306 THEN
            exp_f := 251;
        ELSIF x =- 4305 THEN
            exp_f := 251;
        ELSIF x =- 4304 THEN
            exp_f := 251;
        ELSIF x =- 4303 THEN
            exp_f := 251;
        ELSIF x =- 4302 THEN
            exp_f := 251;
        ELSIF x =- 4301 THEN
            exp_f := 251;
        ELSIF x =- 4300 THEN
            exp_f := 251;
        ELSIF x =- 4299 THEN
            exp_f := 251;
        ELSIF x =- 4298 THEN
            exp_f := 251;
        ELSIF x =- 4297 THEN
            exp_f := 252;
        ELSIF x =- 4296 THEN
            exp_f := 252;
        ELSIF x =- 4295 THEN
            exp_f := 252;
        ELSIF x =- 4294 THEN
            exp_f := 252;
        ELSIF x =- 4293 THEN
            exp_f := 252;
        ELSIF x =- 4292 THEN
            exp_f := 252;
        ELSIF x =- 4291 THEN
            exp_f := 252;
        ELSIF x =- 4290 THEN
            exp_f := 252;
        ELSIF x =- 4289 THEN
            exp_f := 252;
        ELSIF x =- 4288 THEN
            exp_f := 252;
        ELSIF x =- 4287 THEN
            exp_f := 254;
        ELSIF x =- 4286 THEN
            exp_f := 254;
        ELSIF x =- 4285 THEN
            exp_f := 254;
        ELSIF x =- 4284 THEN
            exp_f := 254;
        ELSIF x =- 4283 THEN
            exp_f := 254;
        ELSIF x =- 4282 THEN
            exp_f := 254;
        ELSIF x =- 4281 THEN
            exp_f := 254;
        ELSIF x =- 4280 THEN
            exp_f := 254;
        ELSIF x =- 4279 THEN
            exp_f := 254;
        ELSIF x =- 4278 THEN
            exp_f := 254;
        ELSIF x =- 4277 THEN
            exp_f := 254;
        ELSIF x =- 4276 THEN
            exp_f := 255;
        ELSIF x =- 4275 THEN
            exp_f := 255;
        ELSIF x =- 4274 THEN
            exp_f := 255;
        ELSIF x =- 4273 THEN
            exp_f := 255;
        ELSIF x =- 4272 THEN
            exp_f := 255;
        ELSIF x =- 4271 THEN
            exp_f := 255;
        ELSIF x =- 4270 THEN
            exp_f := 255;
        ELSIF x =- 4269 THEN
            exp_f := 255;
        ELSIF x =- 4268 THEN
            exp_f := 255;
        ELSIF x =- 4267 THEN
            exp_f := 255;
        ELSIF x =- 4266 THEN
            exp_f := 255;
        ELSIF x =- 4265 THEN
            exp_f := 256;
        ELSIF x =- 4264 THEN
            exp_f := 256;
        ELSIF x =- 4263 THEN
            exp_f := 256;
        ELSIF x =- 4262 THEN
            exp_f := 256;
        ELSIF x =- 4261 THEN
            exp_f := 256;
        ELSIF x =- 4260 THEN
            exp_f := 256;
        ELSIF x =- 4259 THEN
            exp_f := 256;
        ELSIF x =- 4258 THEN
            exp_f := 256;
        ELSIF x =- 4257 THEN
            exp_f := 256;
        ELSIF x =- 4256 THEN
            exp_f := 256;
        ELSIF x =- 4255 THEN
            exp_f := 257;
        ELSIF x =- 4254 THEN
            exp_f := 257;
        ELSIF x =- 4253 THEN
            exp_f := 257;
        ELSIF x =- 4252 THEN
            exp_f := 257;
        ELSIF x =- 4251 THEN
            exp_f := 257;
        ELSIF x =- 4250 THEN
            exp_f := 257;
        ELSIF x =- 4249 THEN
            exp_f := 257;
        ELSIF x =- 4248 THEN
            exp_f := 257;
        ELSIF x =- 4247 THEN
            exp_f := 257;
        ELSIF x =- 4246 THEN
            exp_f := 257;
        ELSIF x =- 4245 THEN
            exp_f := 257;
        ELSIF x =- 4244 THEN
            exp_f := 259;
        ELSIF x =- 4243 THEN
            exp_f := 259;
        ELSIF x =- 4242 THEN
            exp_f := 259;
        ELSIF x =- 4241 THEN
            exp_f := 259;
        ELSIF x =- 4240 THEN
            exp_f := 259;
        ELSIF x =- 4239 THEN
            exp_f := 259;
        ELSIF x =- 4238 THEN
            exp_f := 259;
        ELSIF x =- 4237 THEN
            exp_f := 259;
        ELSIF x =- 4236 THEN
            exp_f := 259;
        ELSIF x =- 4235 THEN
            exp_f := 259;
        ELSIF x =- 4234 THEN
            exp_f := 259;
        ELSIF x =- 4233 THEN
            exp_f := 260;
        ELSIF x =- 4232 THEN
            exp_f := 260;
        ELSIF x =- 4231 THEN
            exp_f := 260;
        ELSIF x =- 4230 THEN
            exp_f := 260;
        ELSIF x =- 4229 THEN
            exp_f := 260;
        ELSIF x =- 4228 THEN
            exp_f := 260;
        ELSIF x =- 4227 THEN
            exp_f := 260;
        ELSIF x =- 4226 THEN
            exp_f := 260;
        ELSIF x =- 4225 THEN
            exp_f := 260;
        ELSIF x =- 4224 THEN
            exp_f := 260;
        ELSIF x =- 4223 THEN
            exp_f := 261;
        ELSIF x =- 4222 THEN
            exp_f := 261;
        ELSIF x =- 4221 THEN
            exp_f := 261;
        ELSIF x =- 4220 THEN
            exp_f := 261;
        ELSIF x =- 4219 THEN
            exp_f := 261;
        ELSIF x =- 4218 THEN
            exp_f := 261;
        ELSIF x =- 4217 THEN
            exp_f := 261;
        ELSIF x =- 4216 THEN
            exp_f := 261;
        ELSIF x =- 4215 THEN
            exp_f := 261;
        ELSIF x =- 4214 THEN
            exp_f := 261;
        ELSIF x =- 4213 THEN
            exp_f := 261;
        ELSIF x =- 4212 THEN
            exp_f := 262;
        ELSIF x =- 4211 THEN
            exp_f := 262;
        ELSIF x =- 4210 THEN
            exp_f := 262;
        ELSIF x =- 4209 THEN
            exp_f := 262;
        ELSIF x =- 4208 THEN
            exp_f := 262;
        ELSIF x =- 4207 THEN
            exp_f := 262;
        ELSIF x =- 4206 THEN
            exp_f := 262;
        ELSIF x =- 4205 THEN
            exp_f := 262;
        ELSIF x =- 4204 THEN
            exp_f := 262;
        ELSIF x =- 4203 THEN
            exp_f := 262;
        ELSIF x =- 4202 THEN
            exp_f := 264;
        ELSIF x =- 4201 THEN
            exp_f := 264;
        ELSIF x =- 4200 THEN
            exp_f := 264;
        ELSIF x =- 4199 THEN
            exp_f := 264;
        ELSIF x =- 4198 THEN
            exp_f := 264;
        ELSIF x =- 4197 THEN
            exp_f := 264;
        ELSIF x =- 4196 THEN
            exp_f := 264;
        ELSIF x =- 4195 THEN
            exp_f := 264;
        ELSIF x =- 4194 THEN
            exp_f := 264;
        ELSIF x =- 4193 THEN
            exp_f := 264;
        ELSIF x =- 4192 THEN
            exp_f := 264;
        ELSIF x =- 4191 THEN
            exp_f := 265;
        ELSIF x =- 4190 THEN
            exp_f := 265;
        ELSIF x =- 4189 THEN
            exp_f := 265;
        ELSIF x =- 4188 THEN
            exp_f := 265;
        ELSIF x =- 4187 THEN
            exp_f := 265;
        ELSIF x =- 4186 THEN
            exp_f := 265;
        ELSIF x =- 4185 THEN
            exp_f := 265;
        ELSIF x =- 4184 THEN
            exp_f := 265;
        ELSIF x =- 4183 THEN
            exp_f := 265;
        ELSIF x =- 4182 THEN
            exp_f := 265;
        ELSIF x =- 4181 THEN
            exp_f := 265;
        ELSIF x =- 4180 THEN
            exp_f := 266;
        ELSIF x =- 4179 THEN
            exp_f := 266;
        ELSIF x =- 4178 THEN
            exp_f := 266;
        ELSIF x =- 4177 THEN
            exp_f := 266;
        ELSIF x =- 4176 THEN
            exp_f := 266;
        ELSIF x =- 4175 THEN
            exp_f := 266;
        ELSIF x =- 4174 THEN
            exp_f := 266;
        ELSIF x =- 4173 THEN
            exp_f := 266;
        ELSIF x =- 4172 THEN
            exp_f := 266;
        ELSIF x =- 4171 THEN
            exp_f := 266;
        ELSIF x =- 4170 THEN
            exp_f := 268;
        ELSIF x =- 4169 THEN
            exp_f := 268;
        ELSIF x =- 4168 THEN
            exp_f := 268;
        ELSIF x =- 4167 THEN
            exp_f := 268;
        ELSIF x =- 4166 THEN
            exp_f := 268;
        ELSIF x =- 4165 THEN
            exp_f := 268;
        ELSIF x =- 4164 THEN
            exp_f := 268;
        ELSIF x =- 4163 THEN
            exp_f := 268;
        ELSIF x =- 4162 THEN
            exp_f := 268;
        ELSIF x =- 4161 THEN
            exp_f := 268;
        ELSIF x =- 4160 THEN
            exp_f := 268;
        ELSIF x =- 4159 THEN
            exp_f := 269;
        ELSIF x =- 4158 THEN
            exp_f := 269;
        ELSIF x =- 4157 THEN
            exp_f := 269;
        ELSIF x =- 4156 THEN
            exp_f := 269;
        ELSIF x =- 4155 THEN
            exp_f := 269;
        ELSIF x =- 4154 THEN
            exp_f := 269;
        ELSIF x =- 4153 THEN
            exp_f := 269;
        ELSIF x =- 4152 THEN
            exp_f := 269;
        ELSIF x =- 4151 THEN
            exp_f := 269;
        ELSIF x =- 4150 THEN
            exp_f := 269;
        ELSIF x =- 4149 THEN
            exp_f := 270;
        ELSIF x =- 4148 THEN
            exp_f := 270;
        ELSIF x =- 4147 THEN
            exp_f := 270;
        ELSIF x =- 4146 THEN
            exp_f := 270;
        ELSIF x =- 4145 THEN
            exp_f := 270;
        ELSIF x =- 4144 THEN
            exp_f := 270;
        ELSIF x =- 4143 THEN
            exp_f := 270;
        ELSIF x =- 4142 THEN
            exp_f := 270;
        ELSIF x =- 4141 THEN
            exp_f := 270;
        ELSIF x =- 4140 THEN
            exp_f := 270;
        ELSIF x =- 4139 THEN
            exp_f := 270;
        ELSIF x =- 4138 THEN
            exp_f := 271;
        ELSIF x =- 4137 THEN
            exp_f := 271;
        ELSIF x =- 4136 THEN
            exp_f := 271;
        ELSIF x =- 4135 THEN
            exp_f := 271;
        ELSIF x =- 4134 THEN
            exp_f := 271;
        ELSIF x =- 4133 THEN
            exp_f := 271;
        ELSIF x =- 4132 THEN
            exp_f := 271;
        ELSIF x =- 4131 THEN
            exp_f := 271;
        ELSIF x =- 4130 THEN
            exp_f := 271;
        ELSIF x =- 4129 THEN
            exp_f := 271;
        ELSIF x =- 4128 THEN
            exp_f := 271;
        ELSIF x =- 4127 THEN
            exp_f := 273;
        ELSIF x =- 4126 THEN
            exp_f := 273;
        ELSIF x =- 4125 THEN
            exp_f := 273;
        ELSIF x =- 4124 THEN
            exp_f := 273;
        ELSIF x =- 4123 THEN
            exp_f := 273;
        ELSIF x =- 4122 THEN
            exp_f := 273;
        ELSIF x =- 4121 THEN
            exp_f := 273;
        ELSIF x =- 4120 THEN
            exp_f := 273;
        ELSIF x =- 4119 THEN
            exp_f := 273;
        ELSIF x =- 4118 THEN
            exp_f := 273;
        ELSIF x =- 4117 THEN
            exp_f := 274;
        ELSIF x =- 4116 THEN
            exp_f := 274;
        ELSIF x =- 4115 THEN
            exp_f := 274;
        ELSIF x =- 4114 THEN
            exp_f := 274;
        ELSIF x =- 4113 THEN
            exp_f := 274;
        ELSIF x =- 4112 THEN
            exp_f := 274;
        ELSIF x =- 4111 THEN
            exp_f := 274;
        ELSIF x =- 4110 THEN
            exp_f := 274;
        ELSIF x =- 4109 THEN
            exp_f := 274;
        ELSIF x =- 4108 THEN
            exp_f := 274;
        ELSIF x =- 4107 THEN
            exp_f := 274;
        ELSIF x =- 4106 THEN
            exp_f := 275;
        ELSIF x =- 4105 THEN
            exp_f := 275;
        ELSIF x =- 4104 THEN
            exp_f := 275;
        ELSIF x =- 4103 THEN
            exp_f := 275;
        ELSIF x =- 4102 THEN
            exp_f := 275;
        ELSIF x =- 4101 THEN
            exp_f := 275;
        ELSIF x =- 4100 THEN
            exp_f := 275;
        ELSIF x =- 4099 THEN
            exp_f := 275;
        ELSIF x =- 4098 THEN
            exp_f := 275;
        ELSIF x =- 4097 THEN
            exp_f := 275;
        ELSIF x =- 4096 THEN
            exp_f := 275;
        ELSIF x =- 4095 THEN
            exp_f := 277;
        ELSIF x =- 4094 THEN
            exp_f := 277;
        ELSIF x =- 4093 THEN
            exp_f := 277;
        ELSIF x =- 4092 THEN
            exp_f := 277;
        ELSIF x =- 4091 THEN
            exp_f := 277;
        ELSIF x =- 4090 THEN
            exp_f := 277;
        ELSIF x =- 4089 THEN
            exp_f := 277;
        ELSIF x =- 4088 THEN
            exp_f := 277;
        ELSIF x =- 4087 THEN
            exp_f := 278;
        ELSIF x =- 4086 THEN
            exp_f := 278;
        ELSIF x =- 4085 THEN
            exp_f := 278;
        ELSIF x =- 4084 THEN
            exp_f := 278;
        ELSIF x =- 4083 THEN
            exp_f := 278;
        ELSIF x =- 4082 THEN
            exp_f := 278;
        ELSIF x =- 4081 THEN
            exp_f := 278;
        ELSIF x =- 4080 THEN
            exp_f := 278;
        ELSIF x =- 4079 THEN
            exp_f := 278;
        ELSIF x =- 4078 THEN
            exp_f := 279;
        ELSIF x =- 4077 THEN
            exp_f := 279;
        ELSIF x =- 4076 THEN
            exp_f := 279;
        ELSIF x =- 4075 THEN
            exp_f := 279;
        ELSIF x =- 4074 THEN
            exp_f := 279;
        ELSIF x =- 4073 THEN
            exp_f := 279;
        ELSIF x =- 4072 THEN
            exp_f := 279;
        ELSIF x =- 4071 THEN
            exp_f := 279;
        ELSIF x =- 4070 THEN
            exp_f := 280;
        ELSIF x =- 4069 THEN
            exp_f := 280;
        ELSIF x =- 4068 THEN
            exp_f := 280;
        ELSIF x =- 4067 THEN
            exp_f := 280;
        ELSIF x =- 4066 THEN
            exp_f := 280;
        ELSIF x =- 4065 THEN
            exp_f := 280;
        ELSIF x =- 4064 THEN
            exp_f := 280;
        ELSIF x =- 4063 THEN
            exp_f := 280;
        ELSIF x =- 4062 THEN
            exp_f := 280;
        ELSIF x =- 4061 THEN
            exp_f := 282;
        ELSIF x =- 4060 THEN
            exp_f := 282;
        ELSIF x =- 4059 THEN
            exp_f := 282;
        ELSIF x =- 4058 THEN
            exp_f := 282;
        ELSIF x =- 4057 THEN
            exp_f := 282;
        ELSIF x =- 4056 THEN
            exp_f := 282;
        ELSIF x =- 4055 THEN
            exp_f := 282;
        ELSIF x =- 4054 THEN
            exp_f := 282;
        ELSIF x =- 4053 THEN
            exp_f := 282;
        ELSIF x =- 4052 THEN
            exp_f := 283;
        ELSIF x =- 4051 THEN
            exp_f := 283;
        ELSIF x =- 4050 THEN
            exp_f := 283;
        ELSIF x =- 4049 THEN
            exp_f := 283;
        ELSIF x =- 4048 THEN
            exp_f := 283;
        ELSIF x =- 4047 THEN
            exp_f := 283;
        ELSIF x =- 4046 THEN
            exp_f := 283;
        ELSIF x =- 4045 THEN
            exp_f := 283;
        ELSIF x =- 4044 THEN
            exp_f := 284;
        ELSIF x =- 4043 THEN
            exp_f := 284;
        ELSIF x =- 4042 THEN
            exp_f := 284;
        ELSIF x =- 4041 THEN
            exp_f := 284;
        ELSIF x =- 4040 THEN
            exp_f := 284;
        ELSIF x =- 4039 THEN
            exp_f := 284;
        ELSIF x =- 4038 THEN
            exp_f := 284;
        ELSIF x =- 4037 THEN
            exp_f := 284;
        ELSIF x =- 4036 THEN
            exp_f := 284;
        ELSIF x =- 4035 THEN
            exp_f := 286;
        ELSIF x =- 4034 THEN
            exp_f := 286;
        ELSIF x =- 4033 THEN
            exp_f := 286;
        ELSIF x =- 4032 THEN
            exp_f := 286;
        ELSIF x =- 4031 THEN
            exp_f := 286;
        ELSIF x =- 4030 THEN
            exp_f := 286;
        ELSIF x =- 4029 THEN
            exp_f := 286;
        ELSIF x =- 4028 THEN
            exp_f := 286;
        ELSIF x =- 4027 THEN
            exp_f := 287;
        ELSIF x =- 4026 THEN
            exp_f := 287;
        ELSIF x =- 4025 THEN
            exp_f := 287;
        ELSIF x =- 4024 THEN
            exp_f := 287;
        ELSIF x =- 4023 THEN
            exp_f := 287;
        ELSIF x =- 4022 THEN
            exp_f := 287;
        ELSIF x =- 4021 THEN
            exp_f := 287;
        ELSIF x =- 4020 THEN
            exp_f := 287;
        ELSIF x =- 4019 THEN
            exp_f := 287;
        ELSIF x =- 4018 THEN
            exp_f := 288;
        ELSIF x =- 4017 THEN
            exp_f := 288;
        ELSIF x =- 4016 THEN
            exp_f := 288;
        ELSIF x =- 4015 THEN
            exp_f := 288;
        ELSIF x =- 4014 THEN
            exp_f := 288;
        ELSIF x =- 4013 THEN
            exp_f := 288;
        ELSIF x =- 4012 THEN
            exp_f := 288;
        ELSIF x =- 4011 THEN
            exp_f := 288;
        ELSIF x =- 4010 THEN
            exp_f := 288;
        ELSIF x =- 4009 THEN
            exp_f := 289;
        ELSIF x =- 4008 THEN
            exp_f := 289;
        ELSIF x =- 4007 THEN
            exp_f := 289;
        ELSIF x =- 4006 THEN
            exp_f := 289;
        ELSIF x =- 4005 THEN
            exp_f := 289;
        ELSIF x =- 4004 THEN
            exp_f := 289;
        ELSIF x =- 4003 THEN
            exp_f := 289;
        ELSIF x =- 4002 THEN
            exp_f := 289;
        ELSIF x =- 4001 THEN
            exp_f := 291;
        ELSIF x =- 4000 THEN
            exp_f := 291;
        ELSIF x =- 3999 THEN
            exp_f := 291;
        ELSIF x =- 3998 THEN
            exp_f := 291;
        ELSIF x =- 3997 THEN
            exp_f := 291;
        ELSIF x =- 3996 THEN
            exp_f := 291;
        ELSIF x =- 3995 THEN
            exp_f := 291;
        ELSIF x =- 3994 THEN
            exp_f := 291;
        ELSIF x =- 3993 THEN
            exp_f := 291;
        ELSIF x =- 3992 THEN
            exp_f := 292;
        ELSIF x =- 3991 THEN
            exp_f := 292;
        ELSIF x =- 3990 THEN
            exp_f := 292;
        ELSIF x =- 3989 THEN
            exp_f := 292;
        ELSIF x =- 3988 THEN
            exp_f := 292;
        ELSIF x =- 3987 THEN
            exp_f := 292;
        ELSIF x =- 3986 THEN
            exp_f := 292;
        ELSIF x =- 3985 THEN
            exp_f := 292;
        ELSIF x =- 3984 THEN
            exp_f := 293;
        ELSIF x =- 3983 THEN
            exp_f := 293;
        ELSIF x =- 3982 THEN
            exp_f := 293;
        ELSIF x =- 3981 THEN
            exp_f := 293;
        ELSIF x =- 3980 THEN
            exp_f := 293;
        ELSIF x =- 3979 THEN
            exp_f := 293;
        ELSIF x =- 3978 THEN
            exp_f := 293;
        ELSIF x =- 3977 THEN
            exp_f := 293;
        ELSIF x =- 3976 THEN
            exp_f := 293;
        ELSIF x =- 3975 THEN
            exp_f := 295;
        ELSIF x =- 3974 THEN
            exp_f := 295;
        ELSIF x =- 3973 THEN
            exp_f := 295;
        ELSIF x =- 3972 THEN
            exp_f := 295;
        ELSIF x =- 3971 THEN
            exp_f := 295;
        ELSIF x =- 3970 THEN
            exp_f := 295;
        ELSIF x =- 3969 THEN
            exp_f := 295;
        ELSIF x =- 3968 THEN
            exp_f := 295;
        ELSIF x =- 3967 THEN
            exp_f := 295;
        ELSIF x =- 3966 THEN
            exp_f := 296;
        ELSIF x =- 3965 THEN
            exp_f := 296;
        ELSIF x =- 3964 THEN
            exp_f := 296;
        ELSIF x =- 3963 THEN
            exp_f := 296;
        ELSIF x =- 3962 THEN
            exp_f := 296;
        ELSIF x =- 3961 THEN
            exp_f := 296;
        ELSIF x =- 3960 THEN
            exp_f := 296;
        ELSIF x =- 3959 THEN
            exp_f := 296;
        ELSIF x =- 3958 THEN
            exp_f := 297;
        ELSIF x =- 3957 THEN
            exp_f := 297;
        ELSIF x =- 3956 THEN
            exp_f := 297;
        ELSIF x =- 3955 THEN
            exp_f := 297;
        ELSIF x =- 3954 THEN
            exp_f := 297;
        ELSIF x =- 3953 THEN
            exp_f := 297;
        ELSIF x =- 3952 THEN
            exp_f := 297;
        ELSIF x =- 3951 THEN
            exp_f := 297;
        ELSIF x =- 3950 THEN
            exp_f := 297;
        ELSIF x =- 3949 THEN
            exp_f := 299;
        ELSIF x =- 3948 THEN
            exp_f := 299;
        ELSIF x =- 3947 THEN
            exp_f := 299;
        ELSIF x =- 3946 THEN
            exp_f := 299;
        ELSIF x =- 3945 THEN
            exp_f := 299;
        ELSIF x =- 3944 THEN
            exp_f := 299;
        ELSIF x =- 3943 THEN
            exp_f := 299;
        ELSIF x =- 3942 THEN
            exp_f := 299;
        ELSIF x =- 3941 THEN
            exp_f := 300;
        ELSIF x =- 3940 THEN
            exp_f := 300;
        ELSIF x =- 3939 THEN
            exp_f := 300;
        ELSIF x =- 3938 THEN
            exp_f := 300;
        ELSIF x =- 3937 THEN
            exp_f := 300;
        ELSIF x =- 3936 THEN
            exp_f := 300;
        ELSIF x =- 3935 THEN
            exp_f := 300;
        ELSIF x =- 3934 THEN
            exp_f := 300;
        ELSIF x =- 3933 THEN
            exp_f := 300;
        ELSIF x =- 3932 THEN
            exp_f := 301;
        ELSIF x =- 3931 THEN
            exp_f := 301;
        ELSIF x =- 3930 THEN
            exp_f := 301;
        ELSIF x =- 3929 THEN
            exp_f := 301;
        ELSIF x =- 3928 THEN
            exp_f := 301;
        ELSIF x =- 3927 THEN
            exp_f := 301;
        ELSIF x =- 3926 THEN
            exp_f := 301;
        ELSIF x =- 3925 THEN
            exp_f := 301;
        ELSIF x =- 3924 THEN
            exp_f := 301;
        ELSIF x =- 3923 THEN
            exp_f := 303;
        ELSIF x =- 3922 THEN
            exp_f := 303;
        ELSIF x =- 3921 THEN
            exp_f := 303;
        ELSIF x =- 3920 THEN
            exp_f := 303;
        ELSIF x =- 3919 THEN
            exp_f := 303;
        ELSIF x =- 3918 THEN
            exp_f := 303;
        ELSIF x =- 3917 THEN
            exp_f := 303;
        ELSIF x =- 3916 THEN
            exp_f := 303;
        ELSIF x =- 3915 THEN
            exp_f := 304;
        ELSIF x =- 3914 THEN
            exp_f := 304;
        ELSIF x =- 3913 THEN
            exp_f := 304;
        ELSIF x =- 3912 THEN
            exp_f := 304;
        ELSIF x =- 3911 THEN
            exp_f := 304;
        ELSIF x =- 3910 THEN
            exp_f := 304;
        ELSIF x =- 3909 THEN
            exp_f := 304;
        ELSIF x =- 3908 THEN
            exp_f := 304;
        ELSIF x =- 3907 THEN
            exp_f := 304;
        ELSIF x =- 3906 THEN
            exp_f := 305;
        ELSIF x =- 3905 THEN
            exp_f := 305;
        ELSIF x =- 3904 THEN
            exp_f := 305;
        ELSIF x =- 3903 THEN
            exp_f := 305;
        ELSIF x =- 3902 THEN
            exp_f := 305;
        ELSIF x =- 3901 THEN
            exp_f := 305;
        ELSIF x =- 3900 THEN
            exp_f := 305;
        ELSIF x =- 3899 THEN
            exp_f := 305;
        ELSIF x =- 3898 THEN
            exp_f := 307;
        ELSIF x =- 3897 THEN
            exp_f := 307;
        ELSIF x =- 3896 THEN
            exp_f := 307;
        ELSIF x =- 3895 THEN
            exp_f := 307;
        ELSIF x =- 3894 THEN
            exp_f := 307;
        ELSIF x =- 3893 THEN
            exp_f := 307;
        ELSIF x =- 3892 THEN
            exp_f := 307;
        ELSIF x =- 3891 THEN
            exp_f := 307;
        ELSIF x =- 3890 THEN
            exp_f := 307;
        ELSIF x =- 3889 THEN
            exp_f := 308;
        ELSIF x =- 3888 THEN
            exp_f := 308;
        ELSIF x =- 3887 THEN
            exp_f := 308;
        ELSIF x =- 3886 THEN
            exp_f := 308;
        ELSIF x =- 3885 THEN
            exp_f := 308;
        ELSIF x =- 3884 THEN
            exp_f := 308;
        ELSIF x =- 3883 THEN
            exp_f := 308;
        ELSIF x =- 3882 THEN
            exp_f := 308;
        ELSIF x =- 3881 THEN
            exp_f := 308;
        ELSIF x =- 3880 THEN
            exp_f := 309;
        ELSIF x =- 3879 THEN
            exp_f := 309;
        ELSIF x =- 3878 THEN
            exp_f := 309;
        ELSIF x =- 3877 THEN
            exp_f := 309;
        ELSIF x =- 3876 THEN
            exp_f := 309;
        ELSIF x =- 3875 THEN
            exp_f := 309;
        ELSIF x =- 3874 THEN
            exp_f := 309;
        ELSIF x =- 3873 THEN
            exp_f := 309;
        ELSIF x =- 3872 THEN
            exp_f := 311;
        ELSIF x =- 3871 THEN
            exp_f := 311;
        ELSIF x =- 3870 THEN
            exp_f := 311;
        ELSIF x =- 3869 THEN
            exp_f := 311;
        ELSIF x =- 3868 THEN
            exp_f := 311;
        ELSIF x =- 3867 THEN
            exp_f := 311;
        ELSIF x =- 3866 THEN
            exp_f := 311;
        ELSIF x =- 3865 THEN
            exp_f := 311;
        ELSIF x =- 3864 THEN
            exp_f := 311;
        ELSIF x =- 3863 THEN
            exp_f := 312;
        ELSIF x =- 3862 THEN
            exp_f := 312;
        ELSIF x =- 3861 THEN
            exp_f := 312;
        ELSIF x =- 3860 THEN
            exp_f := 312;
        ELSIF x =- 3859 THEN
            exp_f := 312;
        ELSIF x =- 3858 THEN
            exp_f := 312;
        ELSIF x =- 3857 THEN
            exp_f := 312;
        ELSIF x =- 3856 THEN
            exp_f := 312;
        ELSIF x =- 3855 THEN
            exp_f := 313;
        ELSIF x =- 3854 THEN
            exp_f := 313;
        ELSIF x =- 3853 THEN
            exp_f := 313;
        ELSIF x =- 3852 THEN
            exp_f := 313;
        ELSIF x =- 3851 THEN
            exp_f := 313;
        ELSIF x =- 3850 THEN
            exp_f := 313;
        ELSIF x =- 3849 THEN
            exp_f := 313;
        ELSIF x =- 3848 THEN
            exp_f := 313;
        ELSIF x =- 3847 THEN
            exp_f := 313;
        ELSIF x =- 3846 THEN
            exp_f := 314;
        ELSIF x =- 3845 THEN
            exp_f := 314;
        ELSIF x =- 3844 THEN
            exp_f := 314;
        ELSIF x =- 3843 THEN
            exp_f := 314;
        ELSIF x =- 3842 THEN
            exp_f := 314;
        ELSIF x =- 3841 THEN
            exp_f := 314;
        ELSIF x =- 3840 THEN
            exp_f := 314;
        ELSIF x =- 3839 THEN
            exp_f := 314;
        ELSIF x =- 3838 THEN
            exp_f := 314;
        ELSIF x =- 3837 THEN
            exp_f := 316;
        ELSIF x =- 3836 THEN
            exp_f := 316;
        ELSIF x =- 3835 THEN
            exp_f := 316;
        ELSIF x =- 3834 THEN
            exp_f := 316;
        ELSIF x =- 3833 THEN
            exp_f := 316;
        ELSIF x =- 3832 THEN
            exp_f := 316;
        ELSIF x =- 3831 THEN
            exp_f := 316;
        ELSIF x =- 3830 THEN
            exp_f := 316;
        ELSIF x =- 3829 THEN
            exp_f := 317;
        ELSIF x =- 3828 THEN
            exp_f := 317;
        ELSIF x =- 3827 THEN
            exp_f := 317;
        ELSIF x =- 3826 THEN
            exp_f := 317;
        ELSIF x =- 3825 THEN
            exp_f := 317;
        ELSIF x =- 3824 THEN
            exp_f := 317;
        ELSIF x =- 3823 THEN
            exp_f := 317;
        ELSIF x =- 3822 THEN
            exp_f := 317;
        ELSIF x =- 3821 THEN
            exp_f := 317;
        ELSIF x =- 3820 THEN
            exp_f := 318;
        ELSIF x =- 3819 THEN
            exp_f := 318;
        ELSIF x =- 3818 THEN
            exp_f := 318;
        ELSIF x =- 3817 THEN
            exp_f := 318;
        ELSIF x =- 3816 THEN
            exp_f := 318;
        ELSIF x =- 3815 THEN
            exp_f := 318;
        ELSIF x =- 3814 THEN
            exp_f := 318;
        ELSIF x =- 3813 THEN
            exp_f := 318;
        ELSIF x =- 3812 THEN
            exp_f := 320;
        ELSIF x =- 3811 THEN
            exp_f := 320;
        ELSIF x =- 3810 THEN
            exp_f := 320;
        ELSIF x =- 3809 THEN
            exp_f := 320;
        ELSIF x =- 3808 THEN
            exp_f := 320;
        ELSIF x =- 3807 THEN
            exp_f := 320;
        ELSIF x =- 3806 THEN
            exp_f := 320;
        ELSIF x =- 3805 THEN
            exp_f := 320;
        ELSIF x =- 3804 THEN
            exp_f := 320;
        ELSIF x =- 3803 THEN
            exp_f := 321;
        ELSIF x =- 3802 THEN
            exp_f := 321;
        ELSIF x =- 3801 THEN
            exp_f := 321;
        ELSIF x =- 3800 THEN
            exp_f := 321;
        ELSIF x =- 3799 THEN
            exp_f := 321;
        ELSIF x =- 3798 THEN
            exp_f := 321;
        ELSIF x =- 3797 THEN
            exp_f := 321;
        ELSIF x =- 3796 THEN
            exp_f := 321;
        ELSIF x =- 3795 THEN
            exp_f := 321;
        ELSIF x =- 3794 THEN
            exp_f := 323;
        ELSIF x =- 3793 THEN
            exp_f := 323;
        ELSIF x =- 3792 THEN
            exp_f := 323;
        ELSIF x =- 3791 THEN
            exp_f := 323;
        ELSIF x =- 3790 THEN
            exp_f := 323;
        ELSIF x =- 3789 THEN
            exp_f := 323;
        ELSIF x =- 3788 THEN
            exp_f := 323;
        ELSIF x =- 3787 THEN
            exp_f := 323;
        ELSIF x =- 3786 THEN
            exp_f := 324;
        ELSIF x =- 3785 THEN
            exp_f := 324;
        ELSIF x =- 3784 THEN
            exp_f := 324;
        ELSIF x =- 3783 THEN
            exp_f := 324;
        ELSIF x =- 3782 THEN
            exp_f := 324;
        ELSIF x =- 3781 THEN
            exp_f := 324;
        ELSIF x =- 3780 THEN
            exp_f := 324;
        ELSIF x =- 3779 THEN
            exp_f := 324;
        ELSIF x =- 3778 THEN
            exp_f := 324;
        ELSIF x =- 3777 THEN
            exp_f := 325;
        ELSIF x =- 3776 THEN
            exp_f := 325;
        ELSIF x =- 3775 THEN
            exp_f := 325;
        ELSIF x =- 3774 THEN
            exp_f := 325;
        ELSIF x =- 3773 THEN
            exp_f := 325;
        ELSIF x =- 3772 THEN
            exp_f := 325;
        ELSIF x =- 3771 THEN
            exp_f := 325;
        ELSIF x =- 3770 THEN
            exp_f := 325;
        ELSIF x =- 3769 THEN
            exp_f := 327;
        ELSIF x =- 3768 THEN
            exp_f := 327;
        ELSIF x =- 3767 THEN
            exp_f := 327;
        ELSIF x =- 3766 THEN
            exp_f := 327;
        ELSIF x =- 3765 THEN
            exp_f := 327;
        ELSIF x =- 3764 THEN
            exp_f := 327;
        ELSIF x =- 3763 THEN
            exp_f := 327;
        ELSIF x =- 3762 THEN
            exp_f := 327;
        ELSIF x =- 3761 THEN
            exp_f := 327;
        ELSIF x =- 3760 THEN
            exp_f := 328;
        ELSIF x =- 3759 THEN
            exp_f := 328;
        ELSIF x =- 3758 THEN
            exp_f := 328;
        ELSIF x =- 3757 THEN
            exp_f := 328;
        ELSIF x =- 3756 THEN
            exp_f := 328;
        ELSIF x =- 3755 THEN
            exp_f := 328;
        ELSIF x =- 3754 THEN
            exp_f := 328;
        ELSIF x =- 3753 THEN
            exp_f := 328;
        ELSIF x =- 3752 THEN
            exp_f := 328;
        ELSIF x =- 3751 THEN
            exp_f := 329;
        ELSIF x =- 3750 THEN
            exp_f := 329;
        ELSIF x =- 3749 THEN
            exp_f := 329;
        ELSIF x =- 3748 THEN
            exp_f := 329;
        ELSIF x =- 3747 THEN
            exp_f := 329;
        ELSIF x =- 3746 THEN
            exp_f := 329;
        ELSIF x =- 3745 THEN
            exp_f := 329;
        ELSIF x =- 3744 THEN
            exp_f := 329;
        ELSIF x =- 3743 THEN
            exp_f := 331;
        ELSIF x =- 3742 THEN
            exp_f := 331;
        ELSIF x =- 3741 THEN
            exp_f := 331;
        ELSIF x =- 3740 THEN
            exp_f := 331;
        ELSIF x =- 3739 THEN
            exp_f := 331;
        ELSIF x =- 3738 THEN
            exp_f := 331;
        ELSIF x =- 3737 THEN
            exp_f := 331;
        ELSIF x =- 3736 THEN
            exp_f := 331;
        ELSIF x =- 3735 THEN
            exp_f := 331;
        ELSIF x =- 3734 THEN
            exp_f := 332;
        ELSIF x =- 3733 THEN
            exp_f := 332;
        ELSIF x =- 3732 THEN
            exp_f := 332;
        ELSIF x =- 3731 THEN
            exp_f := 332;
        ELSIF x =- 3730 THEN
            exp_f := 332;
        ELSIF x =- 3729 THEN
            exp_f := 332;
        ELSIF x =- 3728 THEN
            exp_f := 332;
        ELSIF x =- 3727 THEN
            exp_f := 332;
        ELSIF x =- 3726 THEN
            exp_f := 332;
        ELSIF x =- 3725 THEN
            exp_f := 333;
        ELSIF x =- 3724 THEN
            exp_f := 333;
        ELSIF x =- 3723 THEN
            exp_f := 333;
        ELSIF x =- 3722 THEN
            exp_f := 333;
        ELSIF x =- 3721 THEN
            exp_f := 333;
        ELSIF x =- 3720 THEN
            exp_f := 333;
        ELSIF x =- 3719 THEN
            exp_f := 333;
        ELSIF x =- 3718 THEN
            exp_f := 333;
        ELSIF x =- 3717 THEN
            exp_f := 335;
        ELSIF x =- 3716 THEN
            exp_f := 335;
        ELSIF x =- 3715 THEN
            exp_f := 335;
        ELSIF x =- 3714 THEN
            exp_f := 335;
        ELSIF x =- 3713 THEN
            exp_f := 335;
        ELSIF x =- 3712 THEN
            exp_f := 335;
        ELSIF x =- 3711 THEN
            exp_f := 335;
        ELSIF x =- 3710 THEN
            exp_f := 335;
        ELSIF x =- 3709 THEN
            exp_f := 335;
        ELSIF x =- 3708 THEN
            exp_f := 336;
        ELSIF x =- 3707 THEN
            exp_f := 336;
        ELSIF x =- 3706 THEN
            exp_f := 336;
        ELSIF x =- 3705 THEN
            exp_f := 336;
        ELSIF x =- 3704 THEN
            exp_f := 336;
        ELSIF x =- 3703 THEN
            exp_f := 336;
        ELSIF x =- 3702 THEN
            exp_f := 336;
        ELSIF x =- 3701 THEN
            exp_f := 336;
        ELSIF x =- 3700 THEN
            exp_f := 337;
        ELSIF x =- 3699 THEN
            exp_f := 337;
        ELSIF x =- 3698 THEN
            exp_f := 337;
        ELSIF x =- 3697 THEN
            exp_f := 337;
        ELSIF x =- 3696 THEN
            exp_f := 337;
        ELSIF x =- 3695 THEN
            exp_f := 337;
        ELSIF x =- 3694 THEN
            exp_f := 337;
        ELSIF x =- 3693 THEN
            exp_f := 337;
        ELSIF x =- 3692 THEN
            exp_f := 337;
        ELSIF x =- 3691 THEN
            exp_f := 339;
        ELSIF x =- 3690 THEN
            exp_f := 339;
        ELSIF x =- 3689 THEN
            exp_f := 339;
        ELSIF x =- 3688 THEN
            exp_f := 339;
        ELSIF x =- 3687 THEN
            exp_f := 339;
        ELSIF x =- 3686 THEN
            exp_f := 339;
        ELSIF x =- 3685 THEN
            exp_f := 339;
        ELSIF x =- 3684 THEN
            exp_f := 339;
        ELSIF x =- 3683 THEN
            exp_f := 339;
        ELSIF x =- 3682 THEN
            exp_f := 340;
        ELSIF x =- 3681 THEN
            exp_f := 340;
        ELSIF x =- 3680 THEN
            exp_f := 340;
        ELSIF x =- 3679 THEN
            exp_f := 340;
        ELSIF x =- 3678 THEN
            exp_f := 340;
        ELSIF x =- 3677 THEN
            exp_f := 340;
        ELSIF x =- 3676 THEN
            exp_f := 340;
        ELSIF x =- 3675 THEN
            exp_f := 340;
        ELSIF x =- 3674 THEN
            exp_f := 341;
        ELSIF x =- 3673 THEN
            exp_f := 341;
        ELSIF x =- 3672 THEN
            exp_f := 341;
        ELSIF x =- 3671 THEN
            exp_f := 341;
        ELSIF x =- 3670 THEN
            exp_f := 341;
        ELSIF x =- 3669 THEN
            exp_f := 341;
        ELSIF x =- 3668 THEN
            exp_f := 341;
        ELSIF x =- 3667 THEN
            exp_f := 341;
        ELSIF x =- 3666 THEN
            exp_f := 341;
        ELSIF x =- 3665 THEN
            exp_f := 343;
        ELSIF x =- 3664 THEN
            exp_f := 343;
        ELSIF x =- 3663 THEN
            exp_f := 343;
        ELSIF x =- 3662 THEN
            exp_f := 343;
        ELSIF x =- 3661 THEN
            exp_f := 343;
        ELSIF x =- 3660 THEN
            exp_f := 343;
        ELSIF x =- 3659 THEN
            exp_f := 343;
        ELSIF x =- 3658 THEN
            exp_f := 343;
        ELSIF x =- 3657 THEN
            exp_f := 344;
        ELSIF x =- 3656 THEN
            exp_f := 344;
        ELSIF x =- 3655 THEN
            exp_f := 344;
        ELSIF x =- 3654 THEN
            exp_f := 344;
        ELSIF x =- 3653 THEN
            exp_f := 344;
        ELSIF x =- 3652 THEN
            exp_f := 344;
        ELSIF x =- 3651 THEN
            exp_f := 344;
        ELSIF x =- 3650 THEN
            exp_f := 344;
        ELSIF x =- 3649 THEN
            exp_f := 344;
        ELSIF x =- 3648 THEN
            exp_f := 346;
        ELSIF x =- 3647 THEN
            exp_f := 346;
        ELSIF x =- 3646 THEN
            exp_f := 346;
        ELSIF x =- 3645 THEN
            exp_f := 346;
        ELSIF x =- 3644 THEN
            exp_f := 346;
        ELSIF x =- 3643 THEN
            exp_f := 346;
        ELSIF x =- 3642 THEN
            exp_f := 346;
        ELSIF x =- 3641 THEN
            exp_f := 346;
        ELSIF x =- 3640 THEN
            exp_f := 346;
        ELSIF x =- 3639 THEN
            exp_f := 347;
        ELSIF x =- 3638 THEN
            exp_f := 347;
        ELSIF x =- 3637 THEN
            exp_f := 347;
        ELSIF x =- 3636 THEN
            exp_f := 347;
        ELSIF x =- 3635 THEN
            exp_f := 347;
        ELSIF x =- 3634 THEN
            exp_f := 347;
        ELSIF x =- 3633 THEN
            exp_f := 347;
        ELSIF x =- 3632 THEN
            exp_f := 347;
        ELSIF x =- 3631 THEN
            exp_f := 348;
        ELSIF x =- 3630 THEN
            exp_f := 348;
        ELSIF x =- 3629 THEN
            exp_f := 348;
        ELSIF x =- 3628 THEN
            exp_f := 348;
        ELSIF x =- 3627 THEN
            exp_f := 348;
        ELSIF x =- 3626 THEN
            exp_f := 348;
        ELSIF x =- 3625 THEN
            exp_f := 348;
        ELSIF x =- 3624 THEN
            exp_f := 348;
        ELSIF x =- 3623 THEN
            exp_f := 348;
        ELSIF x =- 3622 THEN
            exp_f := 350;
        ELSIF x =- 3621 THEN
            exp_f := 350;
        ELSIF x =- 3620 THEN
            exp_f := 350;
        ELSIF x =- 3619 THEN
            exp_f := 350;
        ELSIF x =- 3618 THEN
            exp_f := 350;
        ELSIF x =- 3617 THEN
            exp_f := 350;
        ELSIF x =- 3616 THEN
            exp_f := 350;
        ELSIF x =- 3615 THEN
            exp_f := 350;
        ELSIF x =- 3614 THEN
            exp_f := 351;
        ELSIF x =- 3613 THEN
            exp_f := 351;
        ELSIF x =- 3612 THEN
            exp_f := 351;
        ELSIF x =- 3611 THEN
            exp_f := 351;
        ELSIF x =- 3610 THEN
            exp_f := 351;
        ELSIF x =- 3609 THEN
            exp_f := 351;
        ELSIF x =- 3608 THEN
            exp_f := 351;
        ELSIF x =- 3607 THEN
            exp_f := 351;
        ELSIF x =- 3606 THEN
            exp_f := 351;
        ELSIF x =- 3605 THEN
            exp_f := 352;
        ELSIF x =- 3604 THEN
            exp_f := 352;
        ELSIF x =- 3603 THEN
            exp_f := 352;
        ELSIF x =- 3602 THEN
            exp_f := 352;
        ELSIF x =- 3601 THEN
            exp_f := 352;
        ELSIF x =- 3600 THEN
            exp_f := 352;
        ELSIF x =- 3599 THEN
            exp_f := 352;
        ELSIF x =- 3598 THEN
            exp_f := 352;
        ELSIF x =- 3597 THEN
            exp_f := 352;
        ELSIF x =- 3596 THEN
            exp_f := 354;
        ELSIF x =- 3595 THEN
            exp_f := 354;
        ELSIF x =- 3594 THEN
            exp_f := 354;
        ELSIF x =- 3593 THEN
            exp_f := 354;
        ELSIF x =- 3592 THEN
            exp_f := 354;
        ELSIF x =- 3591 THEN
            exp_f := 354;
        ELSIF x =- 3590 THEN
            exp_f := 354;
        ELSIF x =- 3589 THEN
            exp_f := 354;
        ELSIF x =- 3588 THEN
            exp_f := 355;
        ELSIF x =- 3587 THEN
            exp_f := 355;
        ELSIF x =- 3586 THEN
            exp_f := 355;
        ELSIF x =- 3585 THEN
            exp_f := 355;
        ELSIF x =- 3584 THEN
            exp_f := 355;
        ELSIF x =- 3583 THEN
            exp_f := 355;
        ELSIF x =- 3582 THEN
            exp_f := 355;
        ELSIF x =- 3581 THEN
            exp_f := 355;
        ELSIF x =- 3580 THEN
            exp_f := 355;
        ELSIF x =- 3579 THEN
            exp_f := 355;
        ELSIF x =- 3578 THEN
            exp_f := 356;
        ELSIF x =- 3577 THEN
            exp_f := 356;
        ELSIF x =- 3576 THEN
            exp_f := 356;
        ELSIF x =- 3575 THEN
            exp_f := 356;
        ELSIF x =- 3574 THEN
            exp_f := 356;
        ELSIF x =- 3573 THEN
            exp_f := 356;
        ELSIF x =- 3572 THEN
            exp_f := 356;
        ELSIF x =- 3571 THEN
            exp_f := 358;
        ELSIF x =- 3570 THEN
            exp_f := 358;
        ELSIF x =- 3569 THEN
            exp_f := 358;
        ELSIF x =- 3568 THEN
            exp_f := 358;
        ELSIF x =- 3567 THEN
            exp_f := 358;
        ELSIF x =- 3566 THEN
            exp_f := 358;
        ELSIF x =- 3565 THEN
            exp_f := 358;
        ELSIF x =- 3564 THEN
            exp_f := 358;
        ELSIF x =- 3563 THEN
            exp_f := 359;
        ELSIF x =- 3562 THEN
            exp_f := 359;
        ELSIF x =- 3561 THEN
            exp_f := 359;
        ELSIF x =- 3560 THEN
            exp_f := 359;
        ELSIF x =- 3559 THEN
            exp_f := 359;
        ELSIF x =- 3558 THEN
            exp_f := 359;
        ELSIF x =- 3557 THEN
            exp_f := 359;
        ELSIF x =- 3556 THEN
            exp_f := 361;
        ELSIF x =- 3555 THEN
            exp_f := 361;
        ELSIF x =- 3554 THEN
            exp_f := 361;
        ELSIF x =- 3553 THEN
            exp_f := 361;
        ELSIF x =- 3552 THEN
            exp_f := 361;
        ELSIF x =- 3551 THEN
            exp_f := 361;
        ELSIF x =- 3550 THEN
            exp_f := 361;
        ELSIF x =- 3549 THEN
            exp_f := 362;
        ELSIF x =- 3548 THEN
            exp_f := 362;
        ELSIF x =- 3547 THEN
            exp_f := 362;
        ELSIF x =- 3546 THEN
            exp_f := 362;
        ELSIF x =- 3545 THEN
            exp_f := 362;
        ELSIF x =- 3544 THEN
            exp_f := 362;
        ELSIF x =- 3543 THEN
            exp_f := 362;
        ELSIF x =- 3542 THEN
            exp_f := 363;
        ELSIF x =- 3541 THEN
            exp_f := 363;
        ELSIF x =- 3540 THEN
            exp_f := 363;
        ELSIF x =- 3539 THEN
            exp_f := 363;
        ELSIF x =- 3538 THEN
            exp_f := 363;
        ELSIF x =- 3537 THEN
            exp_f := 363;
        ELSIF x =- 3536 THEN
            exp_f := 363;
        ELSIF x =- 3535 THEN
            exp_f := 363;
        ELSIF x =- 3534 THEN
            exp_f := 365;
        ELSIF x =- 3533 THEN
            exp_f := 365;
        ELSIF x =- 3532 THEN
            exp_f := 365;
        ELSIF x =- 3531 THEN
            exp_f := 365;
        ELSIF x =- 3530 THEN
            exp_f := 365;
        ELSIF x =- 3529 THEN
            exp_f := 365;
        ELSIF x =- 3528 THEN
            exp_f := 365;
        ELSIF x =- 3527 THEN
            exp_f := 366;
        ELSIF x =- 3526 THEN
            exp_f := 366;
        ELSIF x =- 3525 THEN
            exp_f := 366;
        ELSIF x =- 3524 THEN
            exp_f := 366;
        ELSIF x =- 3523 THEN
            exp_f := 366;
        ELSIF x =- 3522 THEN
            exp_f := 366;
        ELSIF x =- 3521 THEN
            exp_f := 366;
        ELSIF x =- 3520 THEN
            exp_f := 368;
        ELSIF x =- 3519 THEN
            exp_f := 368;
        ELSIF x =- 3518 THEN
            exp_f := 368;
        ELSIF x =- 3517 THEN
            exp_f := 368;
        ELSIF x =- 3516 THEN
            exp_f := 368;
        ELSIF x =- 3515 THEN
            exp_f := 368;
        ELSIF x =- 3514 THEN
            exp_f := 368;
        ELSIF x =- 3513 THEN
            exp_f := 368;
        ELSIF x =- 3512 THEN
            exp_f := 369;
        ELSIF x =- 3511 THEN
            exp_f := 369;
        ELSIF x =- 3510 THEN
            exp_f := 369;
        ELSIF x =- 3509 THEN
            exp_f := 369;
        ELSIF x =- 3508 THEN
            exp_f := 369;
        ELSIF x =- 3507 THEN
            exp_f := 369;
        ELSIF x =- 3506 THEN
            exp_f := 369;
        ELSIF x =- 3505 THEN
            exp_f := 370;
        ELSIF x =- 3504 THEN
            exp_f := 370;
        ELSIF x =- 3503 THEN
            exp_f := 370;
        ELSIF x =- 3502 THEN
            exp_f := 370;
        ELSIF x =- 3501 THEN
            exp_f := 370;
        ELSIF x =- 3500 THEN
            exp_f := 370;
        ELSIF x =- 3499 THEN
            exp_f := 370;
        ELSIF x =- 3498 THEN
            exp_f := 372;
        ELSIF x =- 3497 THEN
            exp_f := 372;
        ELSIF x =- 3496 THEN
            exp_f := 372;
        ELSIF x =- 3495 THEN
            exp_f := 372;
        ELSIF x =- 3494 THEN
            exp_f := 372;
        ELSIF x =- 3493 THEN
            exp_f := 372;
        ELSIF x =- 3492 THEN
            exp_f := 372;
        ELSIF x =- 3491 THEN
            exp_f := 373;
        ELSIF x =- 3490 THEN
            exp_f := 373;
        ELSIF x =- 3489 THEN
            exp_f := 373;
        ELSIF x =- 3488 THEN
            exp_f := 373;
        ELSIF x =- 3487 THEN
            exp_f := 373;
        ELSIF x =- 3486 THEN
            exp_f := 373;
        ELSIF x =- 3485 THEN
            exp_f := 373;
        ELSIF x =- 3484 THEN
            exp_f := 373;
        ELSIF x =- 3483 THEN
            exp_f := 375;
        ELSIF x =- 3482 THEN
            exp_f := 375;
        ELSIF x =- 3481 THEN
            exp_f := 375;
        ELSIF x =- 3480 THEN
            exp_f := 375;
        ELSIF x =- 3479 THEN
            exp_f := 375;
        ELSIF x =- 3478 THEN
            exp_f := 375;
        ELSIF x =- 3477 THEN
            exp_f := 375;
        ELSIF x =- 3476 THEN
            exp_f := 376;
        ELSIF x =- 3475 THEN
            exp_f := 376;
        ELSIF x =- 3474 THEN
            exp_f := 376;
        ELSIF x =- 3473 THEN
            exp_f := 376;
        ELSIF x =- 3472 THEN
            exp_f := 376;
        ELSIF x =- 3471 THEN
            exp_f := 376;
        ELSIF x =- 3470 THEN
            exp_f := 376;
        ELSIF x =- 3469 THEN
            exp_f := 377;
        ELSIF x =- 3468 THEN
            exp_f := 377;
        ELSIF x =- 3467 THEN
            exp_f := 377;
        ELSIF x =- 3466 THEN
            exp_f := 377;
        ELSIF x =- 3465 THEN
            exp_f := 377;
        ELSIF x =- 3464 THEN
            exp_f := 377;
        ELSIF x =- 3463 THEN
            exp_f := 377;
        ELSIF x =- 3462 THEN
            exp_f := 377;
        ELSIF x =- 3461 THEN
            exp_f := 379;
        ELSIF x =- 3460 THEN
            exp_f := 379;
        ELSIF x =- 3459 THEN
            exp_f := 379;
        ELSIF x =- 3458 THEN
            exp_f := 379;
        ELSIF x =- 3457 THEN
            exp_f := 379;
        ELSIF x =- 3456 THEN
            exp_f := 379;
        ELSIF x =- 3455 THEN
            exp_f := 379;
        ELSIF x =- 3454 THEN
            exp_f := 380;
        ELSIF x =- 3453 THEN
            exp_f := 380;
        ELSIF x =- 3452 THEN
            exp_f := 380;
        ELSIF x =- 3451 THEN
            exp_f := 380;
        ELSIF x =- 3450 THEN
            exp_f := 380;
        ELSIF x =- 3449 THEN
            exp_f := 380;
        ELSIF x =- 3448 THEN
            exp_f := 380;
        ELSIF x =- 3447 THEN
            exp_f := 382;
        ELSIF x =- 3446 THEN
            exp_f := 382;
        ELSIF x =- 3445 THEN
            exp_f := 382;
        ELSIF x =- 3444 THEN
            exp_f := 382;
        ELSIF x =- 3443 THEN
            exp_f := 382;
        ELSIF x =- 3442 THEN
            exp_f := 382;
        ELSIF x =- 3441 THEN
            exp_f := 382;
        ELSIF x =- 3440 THEN
            exp_f := 383;
        ELSIF x =- 3439 THEN
            exp_f := 383;
        ELSIF x =- 3438 THEN
            exp_f := 383;
        ELSIF x =- 3437 THEN
            exp_f := 383;
        ELSIF x =- 3436 THEN
            exp_f := 383;
        ELSIF x =- 3435 THEN
            exp_f := 383;
        ELSIF x =- 3434 THEN
            exp_f := 383;
        ELSIF x =- 3433 THEN
            exp_f := 383;
        ELSIF x =- 3432 THEN
            exp_f := 384;
        ELSIF x =- 3431 THEN
            exp_f := 384;
        ELSIF x =- 3430 THEN
            exp_f := 384;
        ELSIF x =- 3429 THEN
            exp_f := 384;
        ELSIF x =- 3428 THEN
            exp_f := 384;
        ELSIF x =- 3427 THEN
            exp_f := 384;
        ELSIF x =- 3426 THEN
            exp_f := 384;
        ELSIF x =- 3425 THEN
            exp_f := 386;
        ELSIF x =- 3424 THEN
            exp_f := 386;
        ELSIF x =- 3423 THEN
            exp_f := 386;
        ELSIF x =- 3422 THEN
            exp_f := 386;
        ELSIF x =- 3421 THEN
            exp_f := 386;
        ELSIF x =- 3420 THEN
            exp_f := 386;
        ELSIF x =- 3419 THEN
            exp_f := 386;
        ELSIF x =- 3418 THEN
            exp_f := 387;
        ELSIF x =- 3417 THEN
            exp_f := 387;
        ELSIF x =- 3416 THEN
            exp_f := 387;
        ELSIF x =- 3415 THEN
            exp_f := 387;
        ELSIF x =- 3414 THEN
            exp_f := 387;
        ELSIF x =- 3413 THEN
            exp_f := 387;
        ELSIF x =- 3412 THEN
            exp_f := 387;
        ELSIF x =- 3411 THEN
            exp_f := 387;
        ELSIF x =- 3410 THEN
            exp_f := 389;
        ELSIF x =- 3409 THEN
            exp_f := 389;
        ELSIF x =- 3408 THEN
            exp_f := 389;
        ELSIF x =- 3407 THEN
            exp_f := 389;
        ELSIF x =- 3406 THEN
            exp_f := 389;
        ELSIF x =- 3405 THEN
            exp_f := 389;
        ELSIF x =- 3404 THEN
            exp_f := 389;
        ELSIF x =- 3403 THEN
            exp_f := 390;
        ELSIF x =- 3402 THEN
            exp_f := 390;
        ELSIF x =- 3401 THEN
            exp_f := 390;
        ELSIF x =- 3400 THEN
            exp_f := 390;
        ELSIF x =- 3399 THEN
            exp_f := 390;
        ELSIF x =- 3398 THEN
            exp_f := 390;
        ELSIF x =- 3397 THEN
            exp_f := 390;
        ELSIF x =- 3396 THEN
            exp_f := 391;
        ELSIF x =- 3395 THEN
            exp_f := 391;
        ELSIF x =- 3394 THEN
            exp_f := 391;
        ELSIF x =- 3393 THEN
            exp_f := 391;
        ELSIF x =- 3392 THEN
            exp_f := 391;
        ELSIF x =- 3391 THEN
            exp_f := 391;
        ELSIF x =- 3390 THEN
            exp_f := 391;
        ELSIF x =- 3389 THEN
            exp_f := 393;
        ELSIF x =- 3388 THEN
            exp_f := 393;
        ELSIF x =- 3387 THEN
            exp_f := 393;
        ELSIF x =- 3386 THEN
            exp_f := 393;
        ELSIF x =- 3385 THEN
            exp_f := 393;
        ELSIF x =- 3384 THEN
            exp_f := 393;
        ELSIF x =- 3383 THEN
            exp_f := 393;
        ELSIF x =- 3382 THEN
            exp_f := 393;
        ELSIF x =- 3381 THEN
            exp_f := 394;
        ELSIF x =- 3380 THEN
            exp_f := 394;
        ELSIF x =- 3379 THEN
            exp_f := 394;
        ELSIF x =- 3378 THEN
            exp_f := 394;
        ELSIF x =- 3377 THEN
            exp_f := 394;
        ELSIF x =- 3376 THEN
            exp_f := 394;
        ELSIF x =- 3375 THEN
            exp_f := 394;
        ELSIF x =- 3374 THEN
            exp_f := 396;
        ELSIF x =- 3373 THEN
            exp_f := 396;
        ELSIF x =- 3372 THEN
            exp_f := 396;
        ELSIF x =- 3371 THEN
            exp_f := 396;
        ELSIF x =- 3370 THEN
            exp_f := 396;
        ELSIF x =- 3369 THEN
            exp_f := 396;
        ELSIF x =- 3368 THEN
            exp_f := 396;
        ELSIF x =- 3367 THEN
            exp_f := 397;
        ELSIF x =- 3366 THEN
            exp_f := 397;
        ELSIF x =- 3365 THEN
            exp_f := 397;
        ELSIF x =- 3364 THEN
            exp_f := 397;
        ELSIF x =- 3363 THEN
            exp_f := 397;
        ELSIF x =- 3362 THEN
            exp_f := 397;
        ELSIF x =- 3361 THEN
            exp_f := 397;
        ELSIF x =- 3360 THEN
            exp_f := 397;
        ELSIF x =- 3359 THEN
            exp_f := 399;
        ELSIF x =- 3358 THEN
            exp_f := 399;
        ELSIF x =- 3357 THEN
            exp_f := 399;
        ELSIF x =- 3356 THEN
            exp_f := 399;
        ELSIF x =- 3355 THEN
            exp_f := 399;
        ELSIF x =- 3354 THEN
            exp_f := 399;
        ELSIF x =- 3353 THEN
            exp_f := 399;
        ELSIF x =- 3352 THEN
            exp_f := 400;
        ELSIF x =- 3351 THEN
            exp_f := 400;
        ELSIF x =- 3350 THEN
            exp_f := 400;
        ELSIF x =- 3349 THEN
            exp_f := 400;
        ELSIF x =- 3348 THEN
            exp_f := 400;
        ELSIF x =- 3347 THEN
            exp_f := 400;
        ELSIF x =- 3346 THEN
            exp_f := 400;
        ELSIF x =- 3345 THEN
            exp_f := 401;
        ELSIF x =- 3344 THEN
            exp_f := 401;
        ELSIF x =- 3343 THEN
            exp_f := 401;
        ELSIF x =- 3342 THEN
            exp_f := 401;
        ELSIF x =- 3341 THEN
            exp_f := 401;
        ELSIF x =- 3340 THEN
            exp_f := 401;
        ELSIF x =- 3339 THEN
            exp_f := 401;
        ELSIF x =- 3338 THEN
            exp_f := 403;
        ELSIF x =- 3337 THEN
            exp_f := 403;
        ELSIF x =- 3336 THEN
            exp_f := 403;
        ELSIF x =- 3335 THEN
            exp_f := 403;
        ELSIF x =- 3334 THEN
            exp_f := 403;
        ELSIF x =- 3333 THEN
            exp_f := 403;
        ELSIF x =- 3332 THEN
            exp_f := 403;
        ELSIF x =- 3331 THEN
            exp_f := 403;
        ELSIF x =- 3330 THEN
            exp_f := 404;
        ELSIF x =- 3329 THEN
            exp_f := 404;
        ELSIF x =- 3328 THEN
            exp_f := 404;
        ELSIF x =- 3327 THEN
            exp_f := 404;
        ELSIF x =- 3326 THEN
            exp_f := 404;
        ELSIF x =- 3325 THEN
            exp_f := 404;
        ELSIF x =- 3324 THEN
            exp_f := 404;
        ELSIF x =- 3323 THEN
            exp_f := 406;
        ELSIF x =- 3322 THEN
            exp_f := 406;
        ELSIF x =- 3321 THEN
            exp_f := 406;
        ELSIF x =- 3320 THEN
            exp_f := 406;
        ELSIF x =- 3319 THEN
            exp_f := 406;
        ELSIF x =- 3318 THEN
            exp_f := 406;
        ELSIF x =- 3317 THEN
            exp_f := 406;
        ELSIF x =- 3316 THEN
            exp_f := 407;
        ELSIF x =- 3315 THEN
            exp_f := 407;
        ELSIF x =- 3314 THEN
            exp_f := 407;
        ELSIF x =- 3313 THEN
            exp_f := 407;
        ELSIF x =- 3312 THEN
            exp_f := 407;
        ELSIF x =- 3311 THEN
            exp_f := 407;
        ELSIF x =- 3310 THEN
            exp_f := 407;
        ELSIF x =- 3309 THEN
            exp_f := 407;
        ELSIF x =- 3308 THEN
            exp_f := 409;
        ELSIF x =- 3307 THEN
            exp_f := 409;
        ELSIF x =- 3306 THEN
            exp_f := 409;
        ELSIF x =- 3305 THEN
            exp_f := 409;
        ELSIF x =- 3304 THEN
            exp_f := 409;
        ELSIF x =- 3303 THEN
            exp_f := 409;
        ELSIF x =- 3302 THEN
            exp_f := 409;
        ELSIF x =- 3301 THEN
            exp_f := 410;
        ELSIF x =- 3300 THEN
            exp_f := 410;
        ELSIF x =- 3299 THEN
            exp_f := 410;
        ELSIF x =- 3298 THEN
            exp_f := 410;
        ELSIF x =- 3297 THEN
            exp_f := 410;
        ELSIF x =- 3296 THEN
            exp_f := 410;
        ELSIF x =- 3295 THEN
            exp_f := 410;
        ELSIF x =- 3294 THEN
            exp_f := 412;
        ELSIF x =- 3293 THEN
            exp_f := 412;
        ELSIF x =- 3292 THEN
            exp_f := 412;
        ELSIF x =- 3291 THEN
            exp_f := 412;
        ELSIF x =- 3290 THEN
            exp_f := 412;
        ELSIF x =- 3289 THEN
            exp_f := 412;
        ELSIF x =- 3288 THEN
            exp_f := 412;
        ELSIF x =- 3287 THEN
            exp_f := 413;
        ELSIF x =- 3286 THEN
            exp_f := 413;
        ELSIF x =- 3285 THEN
            exp_f := 413;
        ELSIF x =- 3284 THEN
            exp_f := 413;
        ELSIF x =- 3283 THEN
            exp_f := 413;
        ELSIF x =- 3282 THEN
            exp_f := 413;
        ELSIF x =- 3281 THEN
            exp_f := 413;
        ELSIF x =- 3280 THEN
            exp_f := 413;
        ELSIF x =- 3279 THEN
            exp_f := 414;
        ELSIF x =- 3278 THEN
            exp_f := 414;
        ELSIF x =- 3277 THEN
            exp_f := 414;
        ELSIF x =- 3276 THEN
            exp_f := 414;
        ELSIF x =- 3275 THEN
            exp_f := 414;
        ELSIF x =- 3274 THEN
            exp_f := 414;
        ELSIF x =- 3273 THEN
            exp_f := 414;
        ELSIF x =- 3272 THEN
            exp_f := 416;
        ELSIF x =- 3271 THEN
            exp_f := 416;
        ELSIF x =- 3270 THEN
            exp_f := 416;
        ELSIF x =- 3269 THEN
            exp_f := 416;
        ELSIF x =- 3268 THEN
            exp_f := 416;
        ELSIF x =- 3267 THEN
            exp_f := 416;
        ELSIF x =- 3266 THEN
            exp_f := 416;
        ELSIF x =- 3265 THEN
            exp_f := 417;
        ELSIF x =- 3264 THEN
            exp_f := 417;
        ELSIF x =- 3263 THEN
            exp_f := 417;
        ELSIF x =- 3262 THEN
            exp_f := 417;
        ELSIF x =- 3261 THEN
            exp_f := 417;
        ELSIF x =- 3260 THEN
            exp_f := 417;
        ELSIF x =- 3259 THEN
            exp_f := 417;
        ELSIF x =- 3258 THEN
            exp_f := 417;
        ELSIF x =- 3257 THEN
            exp_f := 419;
        ELSIF x =- 3256 THEN
            exp_f := 419;
        ELSIF x =- 3255 THEN
            exp_f := 419;
        ELSIF x =- 3254 THEN
            exp_f := 419;
        ELSIF x =- 3253 THEN
            exp_f := 419;
        ELSIF x =- 3252 THEN
            exp_f := 419;
        ELSIF x =- 3251 THEN
            exp_f := 419;
        ELSIF x =- 3250 THEN
            exp_f := 420;
        ELSIF x =- 3249 THEN
            exp_f := 420;
        ELSIF x =- 3248 THEN
            exp_f := 420;
        ELSIF x =- 3247 THEN
            exp_f := 420;
        ELSIF x =- 3246 THEN
            exp_f := 420;
        ELSIF x =- 3245 THEN
            exp_f := 420;
        ELSIF x =- 3244 THEN
            exp_f := 420;
        ELSIF x =- 3243 THEN
            exp_f := 422;
        ELSIF x =- 3242 THEN
            exp_f := 422;
        ELSIF x =- 3241 THEN
            exp_f := 422;
        ELSIF x =- 3240 THEN
            exp_f := 422;
        ELSIF x =- 3239 THEN
            exp_f := 422;
        ELSIF x =- 3238 THEN
            exp_f := 422;
        ELSIF x =- 3237 THEN
            exp_f := 422;
        ELSIF x =- 3236 THEN
            exp_f := 422;
        ELSIF x =- 3235 THEN
            exp_f := 423;
        ELSIF x =- 3234 THEN
            exp_f := 423;
        ELSIF x =- 3233 THEN
            exp_f := 423;
        ELSIF x =- 3232 THEN
            exp_f := 423;
        ELSIF x =- 3231 THEN
            exp_f := 423;
        ELSIF x =- 3230 THEN
            exp_f := 423;
        ELSIF x =- 3229 THEN
            exp_f := 423;
        ELSIF x =- 3228 THEN
            exp_f := 425;
        ELSIF x =- 3227 THEN
            exp_f := 425;
        ELSIF x =- 3226 THEN
            exp_f := 425;
        ELSIF x =- 3225 THEN
            exp_f := 425;
        ELSIF x =- 3224 THEN
            exp_f := 425;
        ELSIF x =- 3223 THEN
            exp_f := 425;
        ELSIF x =- 3222 THEN
            exp_f := 425;
        ELSIF x =- 3221 THEN
            exp_f := 426;
        ELSIF x =- 3220 THEN
            exp_f := 426;
        ELSIF x =- 3219 THEN
            exp_f := 426;
        ELSIF x =- 3218 THEN
            exp_f := 426;
        ELSIF x =- 3217 THEN
            exp_f := 426;
        ELSIF x =- 3216 THEN
            exp_f := 426;
        ELSIF x =- 3215 THEN
            exp_f := 426;
        ELSIF x =- 3214 THEN
            exp_f := 427;
        ELSIF x =- 3213 THEN
            exp_f := 427;
        ELSIF x =- 3212 THEN
            exp_f := 427;
        ELSIF x =- 3211 THEN
            exp_f := 427;
        ELSIF x =- 3210 THEN
            exp_f := 427;
        ELSIF x =- 3209 THEN
            exp_f := 427;
        ELSIF x =- 3208 THEN
            exp_f := 427;
        ELSIF x =- 3207 THEN
            exp_f := 427;
        ELSIF x =- 3206 THEN
            exp_f := 429;
        ELSIF x =- 3205 THEN
            exp_f := 429;
        ELSIF x =- 3204 THEN
            exp_f := 429;
        ELSIF x =- 3203 THEN
            exp_f := 429;
        ELSIF x =- 3202 THEN
            exp_f := 429;
        ELSIF x =- 3201 THEN
            exp_f := 429;
        ELSIF x =- 3200 THEN
            exp_f := 429;
        ELSIF x =- 3199 THEN
            exp_f := 430;
        ELSIF x =- 3198 THEN
            exp_f := 430;
        ELSIF x =- 3197 THEN
            exp_f := 430;
        ELSIF x =- 3196 THEN
            exp_f := 430;
        ELSIF x =- 3195 THEN
            exp_f := 430;
        ELSIF x =- 3194 THEN
            exp_f := 430;
        ELSIF x =- 3193 THEN
            exp_f := 430;
        ELSIF x =- 3192 THEN
            exp_f := 432;
        ELSIF x =- 3191 THEN
            exp_f := 432;
        ELSIF x =- 3190 THEN
            exp_f := 432;
        ELSIF x =- 3189 THEN
            exp_f := 432;
        ELSIF x =- 3188 THEN
            exp_f := 432;
        ELSIF x =- 3187 THEN
            exp_f := 432;
        ELSIF x =- 3186 THEN
            exp_f := 432;
        ELSIF x =- 3185 THEN
            exp_f := 432;
        ELSIF x =- 3184 THEN
            exp_f := 433;
        ELSIF x =- 3183 THEN
            exp_f := 433;
        ELSIF x =- 3182 THEN
            exp_f := 433;
        ELSIF x =- 3181 THEN
            exp_f := 433;
        ELSIF x =- 3180 THEN
            exp_f := 433;
        ELSIF x =- 3179 THEN
            exp_f := 433;
        ELSIF x =- 3178 THEN
            exp_f := 433;
        ELSIF x =- 3177 THEN
            exp_f := 435;
        ELSIF x =- 3176 THEN
            exp_f := 435;
        ELSIF x =- 3175 THEN
            exp_f := 435;
        ELSIF x =- 3174 THEN
            exp_f := 435;
        ELSIF x =- 3173 THEN
            exp_f := 435;
        ELSIF x =- 3172 THEN
            exp_f := 435;
        ELSIF x =- 3171 THEN
            exp_f := 435;
        ELSIF x =- 3170 THEN
            exp_f := 436;
        ELSIF x =- 3169 THEN
            exp_f := 436;
        ELSIF x =- 3168 THEN
            exp_f := 436;
        ELSIF x =- 3167 THEN
            exp_f := 436;
        ELSIF x =- 3166 THEN
            exp_f := 436;
        ELSIF x =- 3165 THEN
            exp_f := 436;
        ELSIF x =- 3164 THEN
            exp_f := 436;
        ELSIF x =- 3163 THEN
            exp_f := 438;
        ELSIF x =- 3162 THEN
            exp_f := 438;
        ELSIF x =- 3161 THEN
            exp_f := 438;
        ELSIF x =- 3160 THEN
            exp_f := 438;
        ELSIF x =- 3159 THEN
            exp_f := 438;
        ELSIF x =- 3158 THEN
            exp_f := 438;
        ELSIF x =- 3157 THEN
            exp_f := 438;
        ELSIF x =- 3156 THEN
            exp_f := 438;
        ELSIF x =- 3155 THEN
            exp_f := 439;
        ELSIF x =- 3154 THEN
            exp_f := 439;
        ELSIF x =- 3153 THEN
            exp_f := 439;
        ELSIF x =- 3152 THEN
            exp_f := 439;
        ELSIF x =- 3151 THEN
            exp_f := 439;
        ELSIF x =- 3150 THEN
            exp_f := 439;
        ELSIF x =- 3149 THEN
            exp_f := 439;
        ELSIF x =- 3148 THEN
            exp_f := 441;
        ELSIF x =- 3147 THEN
            exp_f := 441;
        ELSIF x =- 3146 THEN
            exp_f := 441;
        ELSIF x =- 3145 THEN
            exp_f := 441;
        ELSIF x =- 3144 THEN
            exp_f := 441;
        ELSIF x =- 3143 THEN
            exp_f := 441;
        ELSIF x =- 3142 THEN
            exp_f := 441;
        ELSIF x =- 3141 THEN
            exp_f := 442;
        ELSIF x =- 3140 THEN
            exp_f := 442;
        ELSIF x =- 3139 THEN
            exp_f := 442;
        ELSIF x =- 3138 THEN
            exp_f := 442;
        ELSIF x =- 3137 THEN
            exp_f := 442;
        ELSIF x =- 3136 THEN
            exp_f := 442;
        ELSIF x =- 3135 THEN
            exp_f := 442;
        ELSIF x =- 3134 THEN
            exp_f := 442;
        ELSIF x =- 3133 THEN
            exp_f := 444;
        ELSIF x =- 3132 THEN
            exp_f := 444;
        ELSIF x =- 3131 THEN
            exp_f := 444;
        ELSIF x =- 3130 THEN
            exp_f := 444;
        ELSIF x =- 3129 THEN
            exp_f := 444;
        ELSIF x =- 3128 THEN
            exp_f := 444;
        ELSIF x =- 3127 THEN
            exp_f := 444;
        ELSIF x =- 3126 THEN
            exp_f := 445;
        ELSIF x =- 3125 THEN
            exp_f := 445;
        ELSIF x =- 3124 THEN
            exp_f := 445;
        ELSIF x =- 3123 THEN
            exp_f := 445;
        ELSIF x =- 3122 THEN
            exp_f := 445;
        ELSIF x =- 3121 THEN
            exp_f := 445;
        ELSIF x =- 3120 THEN
            exp_f := 445;
        ELSIF x =- 3119 THEN
            exp_f := 447;
        ELSIF x =- 3118 THEN
            exp_f := 447;
        ELSIF x =- 3117 THEN
            exp_f := 447;
        ELSIF x =- 3116 THEN
            exp_f := 447;
        ELSIF x =- 3115 THEN
            exp_f := 447;
        ELSIF x =- 3114 THEN
            exp_f := 447;
        ELSIF x =- 3113 THEN
            exp_f := 447;
        ELSIF x =- 3112 THEN
            exp_f := 448;
        ELSIF x =- 3111 THEN
            exp_f := 448;
        ELSIF x =- 3110 THEN
            exp_f := 448;
        ELSIF x =- 3109 THEN
            exp_f := 448;
        ELSIF x =- 3108 THEN
            exp_f := 448;
        ELSIF x =- 3107 THEN
            exp_f := 448;
        ELSIF x =- 3106 THEN
            exp_f := 448;
        ELSIF x =- 3105 THEN
            exp_f := 448;
        ELSIF x =- 3104 THEN
            exp_f := 450;
        ELSIF x =- 3103 THEN
            exp_f := 450;
        ELSIF x =- 3102 THEN
            exp_f := 450;
        ELSIF x =- 3101 THEN
            exp_f := 450;
        ELSIF x =- 3100 THEN
            exp_f := 450;
        ELSIF x =- 3099 THEN
            exp_f := 450;
        ELSIF x =- 3098 THEN
            exp_f := 450;
        ELSIF x =- 3097 THEN
            exp_f := 451;
        ELSIF x =- 3096 THEN
            exp_f := 451;
        ELSIF x =- 3095 THEN
            exp_f := 451;
        ELSIF x =- 3094 THEN
            exp_f := 451;
        ELSIF x =- 3093 THEN
            exp_f := 451;
        ELSIF x =- 3092 THEN
            exp_f := 451;
        ELSIF x =- 3091 THEN
            exp_f := 451;
        ELSIF x =- 3090 THEN
            exp_f := 453;
        ELSIF x =- 3089 THEN
            exp_f := 453;
        ELSIF x =- 3088 THEN
            exp_f := 453;
        ELSIF x =- 3087 THEN
            exp_f := 453;
        ELSIF x =- 3086 THEN
            exp_f := 453;
        ELSIF x =- 3085 THEN
            exp_f := 453;
        ELSIF x =- 3084 THEN
            exp_f := 453;
        ELSIF x =- 3083 THEN
            exp_f := 453;
        ELSIF x =- 3082 THEN
            exp_f := 454;
        ELSIF x =- 3081 THEN
            exp_f := 454;
        ELSIF x =- 3080 THEN
            exp_f := 454;
        ELSIF x =- 3079 THEN
            exp_f := 454;
        ELSIF x =- 3078 THEN
            exp_f := 454;
        ELSIF x =- 3077 THEN
            exp_f := 454;
        ELSIF x =- 3076 THEN
            exp_f := 454;
        ELSIF x =- 3075 THEN
            exp_f := 456;
        ELSIF x =- 3074 THEN
            exp_f := 456;
        ELSIF x =- 3073 THEN
            exp_f := 456;
        ELSIF x =- 3072 THEN
            exp_f := 456;
        ELSIF x =- 3071 THEN
            exp_f := 456;
        ELSIF x =- 3070 THEN
            exp_f := 456;
        ELSIF x =- 3069 THEN
            exp_f := 456;
        ELSIF x =- 3068 THEN
            exp_f := 457;
        ELSIF x =- 3067 THEN
            exp_f := 457;
        ELSIF x =- 3066 THEN
            exp_f := 457;
        ELSIF x =- 3065 THEN
            exp_f := 457;
        ELSIF x =- 3064 THEN
            exp_f := 457;
        ELSIF x =- 3063 THEN
            exp_f := 457;
        ELSIF x =- 3062 THEN
            exp_f := 459;
        ELSIF x =- 3061 THEN
            exp_f := 459;
        ELSIF x =- 3060 THEN
            exp_f := 459;
        ELSIF x =- 3059 THEN
            exp_f := 459;
        ELSIF x =- 3058 THEN
            exp_f := 459;
        ELSIF x =- 3057 THEN
            exp_f := 459;
        ELSIF x =- 3056 THEN
            exp_f := 460;
        ELSIF x =- 3055 THEN
            exp_f := 460;
        ELSIF x =- 3054 THEN
            exp_f := 460;
        ELSIF x =- 3053 THEN
            exp_f := 460;
        ELSIF x =- 3052 THEN
            exp_f := 460;
        ELSIF x =- 3051 THEN
            exp_f := 460;
        ELSIF x =- 3050 THEN
            exp_f := 462;
        ELSIF x =- 3049 THEN
            exp_f := 462;
        ELSIF x =- 3048 THEN
            exp_f := 462;
        ELSIF x =- 3047 THEN
            exp_f := 462;
        ELSIF x =- 3046 THEN
            exp_f := 462;
        ELSIF x =- 3045 THEN
            exp_f := 462;
        ELSIF x =- 3044 THEN
            exp_f := 462;
        ELSIF x =- 3043 THEN
            exp_f := 463;
        ELSIF x =- 3042 THEN
            exp_f := 463;
        ELSIF x =- 3041 THEN
            exp_f := 463;
        ELSIF x =- 3040 THEN
            exp_f := 463;
        ELSIF x =- 3039 THEN
            exp_f := 463;
        ELSIF x =- 3038 THEN
            exp_f := 463;
        ELSIF x =- 3037 THEN
            exp_f := 465;
        ELSIF x =- 3036 THEN
            exp_f := 465;
        ELSIF x =- 3035 THEN
            exp_f := 465;
        ELSIF x =- 3034 THEN
            exp_f := 465;
        ELSIF x =- 3033 THEN
            exp_f := 465;
        ELSIF x =- 3032 THEN
            exp_f := 465;
        ELSIF x =- 3031 THEN
            exp_f := 466;
        ELSIF x =- 3030 THEN
            exp_f := 466;
        ELSIF x =- 3029 THEN
            exp_f := 466;
        ELSIF x =- 3028 THEN
            exp_f := 466;
        ELSIF x =- 3027 THEN
            exp_f := 466;
        ELSIF x =- 3026 THEN
            exp_f := 466;
        ELSIF x =- 3025 THEN
            exp_f := 468;
        ELSIF x =- 3024 THEN
            exp_f := 468;
        ELSIF x =- 3023 THEN
            exp_f := 468;
        ELSIF x =- 3022 THEN
            exp_f := 468;
        ELSIF x =- 3021 THEN
            exp_f := 468;
        ELSIF x =- 3020 THEN
            exp_f := 468;
        ELSIF x =- 3019 THEN
            exp_f := 469;
        ELSIF x =- 3018 THEN
            exp_f := 469;
        ELSIF x =- 3017 THEN
            exp_f := 469;
        ELSIF x =- 3016 THEN
            exp_f := 469;
        ELSIF x =- 3015 THEN
            exp_f := 469;
        ELSIF x =- 3014 THEN
            exp_f := 469;
        ELSIF x =- 3013 THEN
            exp_f := 469;
        ELSIF x =- 3012 THEN
            exp_f := 471;
        ELSIF x =- 3011 THEN
            exp_f := 471;
        ELSIF x =- 3010 THEN
            exp_f := 471;
        ELSIF x =- 3009 THEN
            exp_f := 471;
        ELSIF x =- 3008 THEN
            exp_f := 471;
        ELSIF x =- 3007 THEN
            exp_f := 471;
        ELSIF x =- 3006 THEN
            exp_f := 472;
        ELSIF x =- 3005 THEN
            exp_f := 472;
        ELSIF x =- 3004 THEN
            exp_f := 472;
        ELSIF x =- 3003 THEN
            exp_f := 472;
        ELSIF x =- 3002 THEN
            exp_f := 472;
        ELSIF x =- 3001 THEN
            exp_f := 472;
        ELSIF x =- 3000 THEN
            exp_f := 474;
        ELSIF x =- 2999 THEN
            exp_f := 474;
        ELSIF x =- 2998 THEN
            exp_f := 474;
        ELSIF x =- 2997 THEN
            exp_f := 474;
        ELSIF x =- 2996 THEN
            exp_f := 474;
        ELSIF x =- 2995 THEN
            exp_f := 474;
        ELSIF x =- 2994 THEN
            exp_f := 475;
        ELSIF x =- 2993 THEN
            exp_f := 475;
        ELSIF x =- 2992 THEN
            exp_f := 475;
        ELSIF x =- 2991 THEN
            exp_f := 475;
        ELSIF x =- 2990 THEN
            exp_f := 475;
        ELSIF x =- 2989 THEN
            exp_f := 475;
        ELSIF x =- 2988 THEN
            exp_f := 475;
        ELSIF x =- 2987 THEN
            exp_f := 477;
        ELSIF x =- 2986 THEN
            exp_f := 477;
        ELSIF x =- 2985 THEN
            exp_f := 477;
        ELSIF x =- 2984 THEN
            exp_f := 477;
        ELSIF x =- 2983 THEN
            exp_f := 477;
        ELSIF x =- 2982 THEN
            exp_f := 477;
        ELSIF x =- 2981 THEN
            exp_f := 478;
        ELSIF x =- 2980 THEN
            exp_f := 478;
        ELSIF x =- 2979 THEN
            exp_f := 478;
        ELSIF x =- 2978 THEN
            exp_f := 478;
        ELSIF x =- 2977 THEN
            exp_f := 478;
        ELSIF x =- 2976 THEN
            exp_f := 478;
        ELSIF x =- 2975 THEN
            exp_f := 480;
        ELSIF x =- 2974 THEN
            exp_f := 480;
        ELSIF x =- 2973 THEN
            exp_f := 480;
        ELSIF x =- 2972 THEN
            exp_f := 480;
        ELSIF x =- 2971 THEN
            exp_f := 480;
        ELSIF x =- 2970 THEN
            exp_f := 480;
        ELSIF x =- 2969 THEN
            exp_f := 481;
        ELSIF x =- 2968 THEN
            exp_f := 481;
        ELSIF x =- 2967 THEN
            exp_f := 481;
        ELSIF x =- 2966 THEN
            exp_f := 481;
        ELSIF x =- 2965 THEN
            exp_f := 481;
        ELSIF x =- 2964 THEN
            exp_f := 481;
        ELSIF x =- 2963 THEN
            exp_f := 483;
        ELSIF x =- 2962 THEN
            exp_f := 483;
        ELSIF x =- 2961 THEN
            exp_f := 483;
        ELSIF x =- 2960 THEN
            exp_f := 483;
        ELSIF x =- 2959 THEN
            exp_f := 483;
        ELSIF x =- 2958 THEN
            exp_f := 483;
        ELSIF x =- 2957 THEN
            exp_f := 483;
        ELSIF x =- 2956 THEN
            exp_f := 484;
        ELSIF x =- 2955 THEN
            exp_f := 484;
        ELSIF x =- 2954 THEN
            exp_f := 484;
        ELSIF x =- 2953 THEN
            exp_f := 484;
        ELSIF x =- 2952 THEN
            exp_f := 484;
        ELSIF x =- 2951 THEN
            exp_f := 484;
        ELSIF x =- 2950 THEN
            exp_f := 486;
        ELSIF x =- 2949 THEN
            exp_f := 486;
        ELSIF x =- 2948 THEN
            exp_f := 486;
        ELSIF x =- 2947 THEN
            exp_f := 486;
        ELSIF x =- 2946 THEN
            exp_f := 486;
        ELSIF x =- 2945 THEN
            exp_f := 486;
        ELSIF x =- 2944 THEN
            exp_f := 487;
        ELSIF x =- 2943 THEN
            exp_f := 487;
        ELSIF x =- 2942 THEN
            exp_f := 487;
        ELSIF x =- 2941 THEN
            exp_f := 487;
        ELSIF x =- 2940 THEN
            exp_f := 487;
        ELSIF x =- 2939 THEN
            exp_f := 487;
        ELSIF x =- 2938 THEN
            exp_f := 489;
        ELSIF x =- 2937 THEN
            exp_f := 489;
        ELSIF x =- 2936 THEN
            exp_f := 489;
        ELSIF x =- 2935 THEN
            exp_f := 489;
        ELSIF x =- 2934 THEN
            exp_f := 489;
        ELSIF x =- 2933 THEN
            exp_f := 489;
        ELSIF x =- 2932 THEN
            exp_f := 489;
        ELSIF x =- 2931 THEN
            exp_f := 490;
        ELSIF x =- 2930 THEN
            exp_f := 490;
        ELSIF x =- 2929 THEN
            exp_f := 490;
        ELSIF x =- 2928 THEN
            exp_f := 490;
        ELSIF x =- 2927 THEN
            exp_f := 490;
        ELSIF x =- 2926 THEN
            exp_f := 490;
        ELSIF x =- 2925 THEN
            exp_f := 492;
        ELSIF x =- 2924 THEN
            exp_f := 492;
        ELSIF x =- 2923 THEN
            exp_f := 492;
        ELSIF x =- 2922 THEN
            exp_f := 492;
        ELSIF x =- 2921 THEN
            exp_f := 492;
        ELSIF x =- 2920 THEN
            exp_f := 492;
        ELSIF x =- 2919 THEN
            exp_f := 494;
        ELSIF x =- 2918 THEN
            exp_f := 494;
        ELSIF x =- 2917 THEN
            exp_f := 494;
        ELSIF x =- 2916 THEN
            exp_f := 494;
        ELSIF x =- 2915 THEN
            exp_f := 494;
        ELSIF x =- 2914 THEN
            exp_f := 494;
        ELSIF x =- 2913 THEN
            exp_f := 495;
        ELSIF x =- 2912 THEN
            exp_f := 495;
        ELSIF x =- 2911 THEN
            exp_f := 495;
        ELSIF x =- 2910 THEN
            exp_f := 495;
        ELSIF x =- 2909 THEN
            exp_f := 495;
        ELSIF x =- 2908 THEN
            exp_f := 495;
        ELSIF x =- 2907 THEN
            exp_f := 497;
        ELSIF x =- 2906 THEN
            exp_f := 497;
        ELSIF x =- 2905 THEN
            exp_f := 497;
        ELSIF x =- 2904 THEN
            exp_f := 497;
        ELSIF x =- 2903 THEN
            exp_f := 497;
        ELSIF x =- 2902 THEN
            exp_f := 497;
        ELSIF x =- 2901 THEN
            exp_f := 497;
        ELSIF x =- 2900 THEN
            exp_f := 498;
        ELSIF x =- 2899 THEN
            exp_f := 498;
        ELSIF x =- 2898 THEN
            exp_f := 498;
        ELSIF x =- 2897 THEN
            exp_f := 498;
        ELSIF x =- 2896 THEN
            exp_f := 498;
        ELSIF x =- 2895 THEN
            exp_f := 498;
        ELSIF x =- 2894 THEN
            exp_f := 500;
        ELSIF x =- 2893 THEN
            exp_f := 500;
        ELSIF x =- 2892 THEN
            exp_f := 500;
        ELSIF x =- 2891 THEN
            exp_f := 500;
        ELSIF x =- 2890 THEN
            exp_f := 500;
        ELSIF x =- 2889 THEN
            exp_f := 500;
        ELSIF x =- 2888 THEN
            exp_f := 501;
        ELSIF x =- 2887 THEN
            exp_f := 501;
        ELSIF x =- 2886 THEN
            exp_f := 501;
        ELSIF x =- 2885 THEN
            exp_f := 501;
        ELSIF x =- 2884 THEN
            exp_f := 501;
        ELSIF x =- 2883 THEN
            exp_f := 501;
        ELSIF x =- 2882 THEN
            exp_f := 503;
        ELSIF x =- 2881 THEN
            exp_f := 503;
        ELSIF x =- 2880 THEN
            exp_f := 503;
        ELSIF x =- 2879 THEN
            exp_f := 503;
        ELSIF x =- 2878 THEN
            exp_f := 503;
        ELSIF x =- 2877 THEN
            exp_f := 503;
        ELSIF x =- 2876 THEN
            exp_f := 503;
        ELSIF x =- 2875 THEN
            exp_f := 504;
        ELSIF x =- 2874 THEN
            exp_f := 504;
        ELSIF x =- 2873 THEN
            exp_f := 504;
        ELSIF x =- 2872 THEN
            exp_f := 504;
        ELSIF x =- 2871 THEN
            exp_f := 504;
        ELSIF x =- 2870 THEN
            exp_f := 504;
        ELSIF x =- 2869 THEN
            exp_f := 506;
        ELSIF x =- 2868 THEN
            exp_f := 506;
        ELSIF x =- 2867 THEN
            exp_f := 506;
        ELSIF x =- 2866 THEN
            exp_f := 506;
        ELSIF x =- 2865 THEN
            exp_f := 506;
        ELSIF x =- 2864 THEN
            exp_f := 506;
        ELSIF x =- 2863 THEN
            exp_f := 507;
        ELSIF x =- 2862 THEN
            exp_f := 507;
        ELSIF x =- 2861 THEN
            exp_f := 507;
        ELSIF x =- 2860 THEN
            exp_f := 507;
        ELSIF x =- 2859 THEN
            exp_f := 507;
        ELSIF x =- 2858 THEN
            exp_f := 507;
        ELSIF x =- 2857 THEN
            exp_f := 509;
        ELSIF x =- 2856 THEN
            exp_f := 509;
        ELSIF x =- 2855 THEN
            exp_f := 509;
        ELSIF x =- 2854 THEN
            exp_f := 509;
        ELSIF x =- 2853 THEN
            exp_f := 509;
        ELSIF x =- 2852 THEN
            exp_f := 509;
        ELSIF x =- 2851 THEN
            exp_f := 511;
        ELSIF x =- 2850 THEN
            exp_f := 511;
        ELSIF x =- 2849 THEN
            exp_f := 511;
        ELSIF x =- 2848 THEN
            exp_f := 511;
        ELSIF x =- 2847 THEN
            exp_f := 511;
        ELSIF x =- 2846 THEN
            exp_f := 511;
        ELSIF x =- 2845 THEN
            exp_f := 511;
        ELSIF x =- 2844 THEN
            exp_f := 512;
        ELSIF x =- 2843 THEN
            exp_f := 512;
        ELSIF x =- 2842 THEN
            exp_f := 512;
        ELSIF x =- 2841 THEN
            exp_f := 512;
        ELSIF x =- 2840 THEN
            exp_f := 512;
        ELSIF x =- 2839 THEN
            exp_f := 512;
        ELSIF x =- 2838 THEN
            exp_f := 514;
        ELSIF x =- 2837 THEN
            exp_f := 514;
        ELSIF x =- 2836 THEN
            exp_f := 514;
        ELSIF x =- 2835 THEN
            exp_f := 514;
        ELSIF x =- 2834 THEN
            exp_f := 514;
        ELSIF x =- 2833 THEN
            exp_f := 514;
        ELSIF x =- 2832 THEN
            exp_f := 515;
        ELSIF x =- 2831 THEN
            exp_f := 515;
        ELSIF x =- 2830 THEN
            exp_f := 515;
        ELSIF x =- 2829 THEN
            exp_f := 515;
        ELSIF x =- 2828 THEN
            exp_f := 515;
        ELSIF x =- 2827 THEN
            exp_f := 515;
        ELSIF x =- 2826 THEN
            exp_f := 517;
        ELSIF x =- 2825 THEN
            exp_f := 517;
        ELSIF x =- 2824 THEN
            exp_f := 517;
        ELSIF x =- 2823 THEN
            exp_f := 517;
        ELSIF x =- 2822 THEN
            exp_f := 517;
        ELSIF x =- 2821 THEN
            exp_f := 517;
        ELSIF x =- 2820 THEN
            exp_f := 517;
        ELSIF x =- 2819 THEN
            exp_f := 518;
        ELSIF x =- 2818 THEN
            exp_f := 518;
        ELSIF x =- 2817 THEN
            exp_f := 518;
        ELSIF x =- 2816 THEN
            exp_f := 518;
        ELSIF x =- 2815 THEN
            exp_f := 518;
        ELSIF x =- 2814 THEN
            exp_f := 518;
        ELSIF x =- 2813 THEN
            exp_f := 520;
        ELSIF x =- 2812 THEN
            exp_f := 520;
        ELSIF x =- 2811 THEN
            exp_f := 520;
        ELSIF x =- 2810 THEN
            exp_f := 520;
        ELSIF x =- 2809 THEN
            exp_f := 520;
        ELSIF x =- 2808 THEN
            exp_f := 520;
        ELSIF x =- 2807 THEN
            exp_f := 522;
        ELSIF x =- 2806 THEN
            exp_f := 522;
        ELSIF x =- 2805 THEN
            exp_f := 522;
        ELSIF x =- 2804 THEN
            exp_f := 522;
        ELSIF x =- 2803 THEN
            exp_f := 522;
        ELSIF x =- 2802 THEN
            exp_f := 522;
        ELSIF x =- 2801 THEN
            exp_f := 523;
        ELSIF x =- 2800 THEN
            exp_f := 523;
        ELSIF x =- 2799 THEN
            exp_f := 523;
        ELSIF x =- 2798 THEN
            exp_f := 523;
        ELSIF x =- 2797 THEN
            exp_f := 523;
        ELSIF x =- 2796 THEN
            exp_f := 523;
        ELSIF x =- 2795 THEN
            exp_f := 523;
        ELSIF x =- 2794 THEN
            exp_f := 525;
        ELSIF x =- 2793 THEN
            exp_f := 525;
        ELSIF x =- 2792 THEN
            exp_f := 525;
        ELSIF x =- 2791 THEN
            exp_f := 525;
        ELSIF x =- 2790 THEN
            exp_f := 525;
        ELSIF x =- 2789 THEN
            exp_f := 525;
        ELSIF x =- 2788 THEN
            exp_f := 526;
        ELSIF x =- 2787 THEN
            exp_f := 526;
        ELSIF x =- 2786 THEN
            exp_f := 526;
        ELSIF x =- 2785 THEN
            exp_f := 526;
        ELSIF x =- 2784 THEN
            exp_f := 526;
        ELSIF x =- 2783 THEN
            exp_f := 526;
        ELSIF x =- 2782 THEN
            exp_f := 528;
        ELSIF x =- 2781 THEN
            exp_f := 528;
        ELSIF x =- 2780 THEN
            exp_f := 528;
        ELSIF x =- 2779 THEN
            exp_f := 528;
        ELSIF x =- 2778 THEN
            exp_f := 528;
        ELSIF x =- 2777 THEN
            exp_f := 528;
        ELSIF x =- 2776 THEN
            exp_f := 529;
        ELSIF x =- 2775 THEN
            exp_f := 529;
        ELSIF x =- 2774 THEN
            exp_f := 529;
        ELSIF x =- 2773 THEN
            exp_f := 529;
        ELSIF x =- 2772 THEN
            exp_f := 529;
        ELSIF x =- 2771 THEN
            exp_f := 529;
        ELSIF x =- 2770 THEN
            exp_f := 531;
        ELSIF x =- 2769 THEN
            exp_f := 531;
        ELSIF x =- 2768 THEN
            exp_f := 531;
        ELSIF x =- 2767 THEN
            exp_f := 531;
        ELSIF x =- 2766 THEN
            exp_f := 531;
        ELSIF x =- 2765 THEN
            exp_f := 531;
        ELSIF x =- 2764 THEN
            exp_f := 531;
        ELSIF x =- 2763 THEN
            exp_f := 533;
        ELSIF x =- 2762 THEN
            exp_f := 533;
        ELSIF x =- 2761 THEN
            exp_f := 533;
        ELSIF x =- 2760 THEN
            exp_f := 533;
        ELSIF x =- 2759 THEN
            exp_f := 533;
        ELSIF x =- 2758 THEN
            exp_f := 533;
        ELSIF x =- 2757 THEN
            exp_f := 534;
        ELSIF x =- 2756 THEN
            exp_f := 534;
        ELSIF x =- 2755 THEN
            exp_f := 534;
        ELSIF x =- 2754 THEN
            exp_f := 534;
        ELSIF x =- 2753 THEN
            exp_f := 534;
        ELSIF x =- 2752 THEN
            exp_f := 534;
        ELSIF x =- 2751 THEN
            exp_f := 536;
        ELSIF x =- 2750 THEN
            exp_f := 536;
        ELSIF x =- 2749 THEN
            exp_f := 536;
        ELSIF x =- 2748 THEN
            exp_f := 536;
        ELSIF x =- 2747 THEN
            exp_f := 536;
        ELSIF x =- 2746 THEN
            exp_f := 536;
        ELSIF x =- 2745 THEN
            exp_f := 537;
        ELSIF x =- 2744 THEN
            exp_f := 537;
        ELSIF x =- 2743 THEN
            exp_f := 537;
        ELSIF x =- 2742 THEN
            exp_f := 537;
        ELSIF x =- 2741 THEN
            exp_f := 537;
        ELSIF x =- 2740 THEN
            exp_f := 537;
        ELSIF x =- 2739 THEN
            exp_f := 537;
        ELSIF x =- 2738 THEN
            exp_f := 539;
        ELSIF x =- 2737 THEN
            exp_f := 539;
        ELSIF x =- 2736 THEN
            exp_f := 539;
        ELSIF x =- 2735 THEN
            exp_f := 539;
        ELSIF x =- 2734 THEN
            exp_f := 539;
        ELSIF x =- 2733 THEN
            exp_f := 539;
        ELSIF x =- 2732 THEN
            exp_f := 541;
        ELSIF x =- 2731 THEN
            exp_f := 541;
        ELSIF x =- 2730 THEN
            exp_f := 541;
        ELSIF x =- 2729 THEN
            exp_f := 541;
        ELSIF x =- 2728 THEN
            exp_f := 541;
        ELSIF x =- 2727 THEN
            exp_f := 541;
        ELSIF x =- 2726 THEN
            exp_f := 542;
        ELSIF x =- 2725 THEN
            exp_f := 542;
        ELSIF x =- 2724 THEN
            exp_f := 542;
        ELSIF x =- 2723 THEN
            exp_f := 542;
        ELSIF x =- 2722 THEN
            exp_f := 542;
        ELSIF x =- 2721 THEN
            exp_f := 542;
        ELSIF x =- 2720 THEN
            exp_f := 544;
        ELSIF x =- 2719 THEN
            exp_f := 544;
        ELSIF x =- 2718 THEN
            exp_f := 544;
        ELSIF x =- 2717 THEN
            exp_f := 544;
        ELSIF x =- 2716 THEN
            exp_f := 544;
        ELSIF x =- 2715 THEN
            exp_f := 544;
        ELSIF x =- 2714 THEN
            exp_f := 545;
        ELSIF x =- 2713 THEN
            exp_f := 545;
        ELSIF x =- 2712 THEN
            exp_f := 545;
        ELSIF x =- 2711 THEN
            exp_f := 545;
        ELSIF x =- 2710 THEN
            exp_f := 545;
        ELSIF x =- 2709 THEN
            exp_f := 545;
        ELSIF x =- 2708 THEN
            exp_f := 545;
        ELSIF x =- 2707 THEN
            exp_f := 547;
        ELSIF x =- 2706 THEN
            exp_f := 547;
        ELSIF x =- 2705 THEN
            exp_f := 547;
        ELSIF x =- 2704 THEN
            exp_f := 547;
        ELSIF x =- 2703 THEN
            exp_f := 547;
        ELSIF x =- 2702 THEN
            exp_f := 547;
        ELSIF x =- 2701 THEN
            exp_f := 549;
        ELSIF x =- 2700 THEN
            exp_f := 549;
        ELSIF x =- 2699 THEN
            exp_f := 549;
        ELSIF x =- 2698 THEN
            exp_f := 549;
        ELSIF x =- 2697 THEN
            exp_f := 549;
        ELSIF x =- 2696 THEN
            exp_f := 549;
        ELSIF x =- 2695 THEN
            exp_f := 550;
        ELSIF x =- 2694 THEN
            exp_f := 550;
        ELSIF x =- 2693 THEN
            exp_f := 550;
        ELSIF x =- 2692 THEN
            exp_f := 550;
        ELSIF x =- 2691 THEN
            exp_f := 550;
        ELSIF x =- 2690 THEN
            exp_f := 550;
        ELSIF x =- 2689 THEN
            exp_f := 552;
        ELSIF x =- 2688 THEN
            exp_f := 552;
        ELSIF x =- 2687 THEN
            exp_f := 552;
        ELSIF x =- 2686 THEN
            exp_f := 552;
        ELSIF x =- 2685 THEN
            exp_f := 552;
        ELSIF x =- 2684 THEN
            exp_f := 552;
        ELSIF x =- 2683 THEN
            exp_f := 552;
        ELSIF x =- 2682 THEN
            exp_f := 553;
        ELSIF x =- 2681 THEN
            exp_f := 553;
        ELSIF x =- 2680 THEN
            exp_f := 553;
        ELSIF x =- 2679 THEN
            exp_f := 553;
        ELSIF x =- 2678 THEN
            exp_f := 553;
        ELSIF x =- 2677 THEN
            exp_f := 553;
        ELSIF x =- 2676 THEN
            exp_f := 555;
        ELSIF x =- 2675 THEN
            exp_f := 555;
        ELSIF x =- 2674 THEN
            exp_f := 555;
        ELSIF x =- 2673 THEN
            exp_f := 555;
        ELSIF x =- 2672 THEN
            exp_f := 555;
        ELSIF x =- 2671 THEN
            exp_f := 555;
        ELSIF x =- 2670 THEN
            exp_f := 557;
        ELSIF x =- 2669 THEN
            exp_f := 557;
        ELSIF x =- 2668 THEN
            exp_f := 557;
        ELSIF x =- 2667 THEN
            exp_f := 557;
        ELSIF x =- 2666 THEN
            exp_f := 557;
        ELSIF x =- 2665 THEN
            exp_f := 557;
        ELSIF x =- 2664 THEN
            exp_f := 558;
        ELSIF x =- 2663 THEN
            exp_f := 558;
        ELSIF x =- 2662 THEN
            exp_f := 558;
        ELSIF x =- 2661 THEN
            exp_f := 558;
        ELSIF x =- 2660 THEN
            exp_f := 558;
        ELSIF x =- 2659 THEN
            exp_f := 558;
        ELSIF x =- 2658 THEN
            exp_f := 560;
        ELSIF x =- 2657 THEN
            exp_f := 560;
        ELSIF x =- 2656 THEN
            exp_f := 560;
        ELSIF x =- 2655 THEN
            exp_f := 560;
        ELSIF x =- 2654 THEN
            exp_f := 560;
        ELSIF x =- 2653 THEN
            exp_f := 560;
        ELSIF x =- 2652 THEN
            exp_f := 560;
        ELSIF x =- 2651 THEN
            exp_f := 562;
        ELSIF x =- 2650 THEN
            exp_f := 562;
        ELSIF x =- 2649 THEN
            exp_f := 562;
        ELSIF x =- 2648 THEN
            exp_f := 562;
        ELSIF x =- 2647 THEN
            exp_f := 562;
        ELSIF x =- 2646 THEN
            exp_f := 562;
        ELSIF x =- 2645 THEN
            exp_f := 563;
        ELSIF x =- 2644 THEN
            exp_f := 563;
        ELSIF x =- 2643 THEN
            exp_f := 563;
        ELSIF x =- 2642 THEN
            exp_f := 563;
        ELSIF x =- 2641 THEN
            exp_f := 563;
        ELSIF x =- 2640 THEN
            exp_f := 563;
        ELSIF x =- 2639 THEN
            exp_f := 565;
        ELSIF x =- 2638 THEN
            exp_f := 565;
        ELSIF x =- 2637 THEN
            exp_f := 565;
        ELSIF x =- 2636 THEN
            exp_f := 565;
        ELSIF x =- 2635 THEN
            exp_f := 565;
        ELSIF x =- 2634 THEN
            exp_f := 565;
        ELSIF x =- 2633 THEN
            exp_f := 566;
        ELSIF x =- 2632 THEN
            exp_f := 566;
        ELSIF x =- 2631 THEN
            exp_f := 566;
        ELSIF x =- 2630 THEN
            exp_f := 566;
        ELSIF x =- 2629 THEN
            exp_f := 566;
        ELSIF x =- 2628 THEN
            exp_f := 566;
        ELSIF x =- 2627 THEN
            exp_f := 566;
        ELSIF x =- 2626 THEN
            exp_f := 568;
        ELSIF x =- 2625 THEN
            exp_f := 568;
        ELSIF x =- 2624 THEN
            exp_f := 568;
        ELSIF x =- 2623 THEN
            exp_f := 568;
        ELSIF x =- 2622 THEN
            exp_f := 568;
        ELSIF x =- 2621 THEN
            exp_f := 568;
        ELSIF x =- 2620 THEN
            exp_f := 570;
        ELSIF x =- 2619 THEN
            exp_f := 570;
        ELSIF x =- 2618 THEN
            exp_f := 570;
        ELSIF x =- 2617 THEN
            exp_f := 570;
        ELSIF x =- 2616 THEN
            exp_f := 570;
        ELSIF x =- 2615 THEN
            exp_f := 570;
        ELSIF x =- 2614 THEN
            exp_f := 571;
        ELSIF x =- 2613 THEN
            exp_f := 571;
        ELSIF x =- 2612 THEN
            exp_f := 571;
        ELSIF x =- 2611 THEN
            exp_f := 571;
        ELSIF x =- 2610 THEN
            exp_f := 571;
        ELSIF x =- 2609 THEN
            exp_f := 571;
        ELSIF x =- 2608 THEN
            exp_f := 573;
        ELSIF x =- 2607 THEN
            exp_f := 573;
        ELSIF x =- 2606 THEN
            exp_f := 573;
        ELSIF x =- 2605 THEN
            exp_f := 573;
        ELSIF x =- 2604 THEN
            exp_f := 573;
        ELSIF x =- 2603 THEN
            exp_f := 573;
        ELSIF x =- 2602 THEN
            exp_f := 575;
        ELSIF x =- 2601 THEN
            exp_f := 575;
        ELSIF x =- 2600 THEN
            exp_f := 575;
        ELSIF x =- 2599 THEN
            exp_f := 575;
        ELSIF x =- 2598 THEN
            exp_f := 575;
        ELSIF x =- 2597 THEN
            exp_f := 575;
        ELSIF x =- 2596 THEN
            exp_f := 575;
        ELSIF x =- 2595 THEN
            exp_f := 576;
        ELSIF x =- 2594 THEN
            exp_f := 576;
        ELSIF x =- 2593 THEN
            exp_f := 576;
        ELSIF x =- 2592 THEN
            exp_f := 576;
        ELSIF x =- 2591 THEN
            exp_f := 576;
        ELSIF x =- 2590 THEN
            exp_f := 576;
        ELSIF x =- 2589 THEN
            exp_f := 578;
        ELSIF x =- 2588 THEN
            exp_f := 578;
        ELSIF x =- 2587 THEN
            exp_f := 578;
        ELSIF x =- 2586 THEN
            exp_f := 578;
        ELSIF x =- 2585 THEN
            exp_f := 578;
        ELSIF x =- 2584 THEN
            exp_f := 578;
        ELSIF x =- 2583 THEN
            exp_f := 580;
        ELSIF x =- 2582 THEN
            exp_f := 580;
        ELSIF x =- 2581 THEN
            exp_f := 580;
        ELSIF x =- 2580 THEN
            exp_f := 580;
        ELSIF x =- 2579 THEN
            exp_f := 580;
        ELSIF x =- 2578 THEN
            exp_f := 580;
        ELSIF x =- 2577 THEN
            exp_f := 581;
        ELSIF x =- 2576 THEN
            exp_f := 581;
        ELSIF x =- 2575 THEN
            exp_f := 581;
        ELSIF x =- 2574 THEN
            exp_f := 581;
        ELSIF x =- 2573 THEN
            exp_f := 581;
        ELSIF x =- 2572 THEN
            exp_f := 581;
        ELSIF x =- 2571 THEN
            exp_f := 581;
        ELSIF x =- 2570 THEN
            exp_f := 583;
        ELSIF x =- 2569 THEN
            exp_f := 583;
        ELSIF x =- 2568 THEN
            exp_f := 583;
        ELSIF x =- 2567 THEN
            exp_f := 583;
        ELSIF x =- 2566 THEN
            exp_f := 583;
        ELSIF x =- 2565 THEN
            exp_f := 583;
        ELSIF x =- 2564 THEN
            exp_f := 584;
        ELSIF x =- 2563 THEN
            exp_f := 584;
        ELSIF x =- 2562 THEN
            exp_f := 584;
        ELSIF x =- 2561 THEN
            exp_f := 584;
        ELSIF x =- 2560 THEN
            exp_f := 584;
        ELSIF x =- 2559 THEN
            exp_f := 584;
        ELSIF x =- 2558 THEN
            exp_f := 586;
        ELSIF x =- 2557 THEN
            exp_f := 586;
        ELSIF x =- 2556 THEN
            exp_f := 586;
        ELSIF x =- 2555 THEN
            exp_f := 586;
        ELSIF x =- 2554 THEN
            exp_f := 586;
        ELSIF x =- 2553 THEN
            exp_f := 588;
        ELSIF x =- 2552 THEN
            exp_f := 588;
        ELSIF x =- 2551 THEN
            exp_f := 588;
        ELSIF x =- 2550 THEN
            exp_f := 588;
        ELSIF x =- 2549 THEN
            exp_f := 588;
        ELSIF x =- 2548 THEN
            exp_f := 588;
        ELSIF x =- 2547 THEN
            exp_f := 589;
        ELSIF x =- 2546 THEN
            exp_f := 589;
        ELSIF x =- 2545 THEN
            exp_f := 589;
        ELSIF x =- 2544 THEN
            exp_f := 589;
        ELSIF x =- 2543 THEN
            exp_f := 589;
        ELSIF x =- 2542 THEN
            exp_f := 591;
        ELSIF x =- 2541 THEN
            exp_f := 591;
        ELSIF x =- 2540 THEN
            exp_f := 591;
        ELSIF x =- 2539 THEN
            exp_f := 591;
        ELSIF x =- 2538 THEN
            exp_f := 591;
        ELSIF x =- 2537 THEN
            exp_f := 593;
        ELSIF x =- 2536 THEN
            exp_f := 593;
        ELSIF x =- 2535 THEN
            exp_f := 593;
        ELSIF x =- 2534 THEN
            exp_f := 593;
        ELSIF x =- 2533 THEN
            exp_f := 593;
        ELSIF x =- 2532 THEN
            exp_f := 593;
        ELSIF x =- 2531 THEN
            exp_f := 594;
        ELSIF x =- 2530 THEN
            exp_f := 594;
        ELSIF x =- 2529 THEN
            exp_f := 594;
        ELSIF x =- 2528 THEN
            exp_f := 594;
        ELSIF x =- 2527 THEN
            exp_f := 594;
        ELSIF x =- 2526 THEN
            exp_f := 596;
        ELSIF x =- 2525 THEN
            exp_f := 596;
        ELSIF x =- 2524 THEN
            exp_f := 596;
        ELSIF x =- 2523 THEN
            exp_f := 596;
        ELSIF x =- 2522 THEN
            exp_f := 596;
        ELSIF x =- 2521 THEN
            exp_f := 598;
        ELSIF x =- 2520 THEN
            exp_f := 598;
        ELSIF x =- 2519 THEN
            exp_f := 598;
        ELSIF x =- 2518 THEN
            exp_f := 598;
        ELSIF x =- 2517 THEN
            exp_f := 598;
        ELSIF x =- 2516 THEN
            exp_f := 598;
        ELSIF x =- 2515 THEN
            exp_f := 599;
        ELSIF x =- 2514 THEN
            exp_f := 599;
        ELSIF x =- 2513 THEN
            exp_f := 599;
        ELSIF x =- 2512 THEN
            exp_f := 599;
        ELSIF x =- 2511 THEN
            exp_f := 599;
        ELSIF x =- 2510 THEN
            exp_f := 601;
        ELSIF x =- 2509 THEN
            exp_f := 601;
        ELSIF x =- 2508 THEN
            exp_f := 601;
        ELSIF x =- 2507 THEN
            exp_f := 601;
        ELSIF x =- 2506 THEN
            exp_f := 601;
        ELSIF x =- 2505 THEN
            exp_f := 601;
        ELSIF x =- 2504 THEN
            exp_f := 603;
        ELSIF x =- 2503 THEN
            exp_f := 603;
        ELSIF x =- 2502 THEN
            exp_f := 603;
        ELSIF x =- 2501 THEN
            exp_f := 603;
        ELSIF x =- 2500 THEN
            exp_f := 603;
        ELSIF x =- 2499 THEN
            exp_f := 604;
        ELSIF x =- 2498 THEN
            exp_f := 604;
        ELSIF x =- 2497 THEN
            exp_f := 604;
        ELSIF x =- 2496 THEN
            exp_f := 604;
        ELSIF x =- 2495 THEN
            exp_f := 604;
        ELSIF x =- 2494 THEN
            exp_f := 606;
        ELSIF x =- 2493 THEN
            exp_f := 606;
        ELSIF x =- 2492 THEN
            exp_f := 606;
        ELSIF x =- 2491 THEN
            exp_f := 606;
        ELSIF x =- 2490 THEN
            exp_f := 606;
        ELSIF x =- 2489 THEN
            exp_f := 606;
        ELSIF x =- 2488 THEN
            exp_f := 608;
        ELSIF x =- 2487 THEN
            exp_f := 608;
        ELSIF x =- 2486 THEN
            exp_f := 608;
        ELSIF x =- 2485 THEN
            exp_f := 608;
        ELSIF x =- 2484 THEN
            exp_f := 608;
        ELSIF x =- 2483 THEN
            exp_f := 609;
        ELSIF x =- 2482 THEN
            exp_f := 609;
        ELSIF x =- 2481 THEN
            exp_f := 609;
        ELSIF x =- 2480 THEN
            exp_f := 609;
        ELSIF x =- 2479 THEN
            exp_f := 609;
        ELSIF x =- 2478 THEN
            exp_f := 611;
        ELSIF x =- 2477 THEN
            exp_f := 611;
        ELSIF x =- 2476 THEN
            exp_f := 611;
        ELSIF x =- 2475 THEN
            exp_f := 611;
        ELSIF x =- 2474 THEN
            exp_f := 611;
        ELSIF x =- 2473 THEN
            exp_f := 611;
        ELSIF x =- 2472 THEN
            exp_f := 613;
        ELSIF x =- 2471 THEN
            exp_f := 613;
        ELSIF x =- 2470 THEN
            exp_f := 613;
        ELSIF x =- 2469 THEN
            exp_f := 613;
        ELSIF x =- 2468 THEN
            exp_f := 613;
        ELSIF x =- 2467 THEN
            exp_f := 615;
        ELSIF x =- 2466 THEN
            exp_f := 615;
        ELSIF x =- 2465 THEN
            exp_f := 615;
        ELSIF x =- 2464 THEN
            exp_f := 615;
        ELSIF x =- 2463 THEN
            exp_f := 615;
        ELSIF x =- 2462 THEN
            exp_f := 615;
        ELSIF x =- 2461 THEN
            exp_f := 616;
        ELSIF x =- 2460 THEN
            exp_f := 616;
        ELSIF x =- 2459 THEN
            exp_f := 616;
        ELSIF x =- 2458 THEN
            exp_f := 616;
        ELSIF x =- 2457 THEN
            exp_f := 616;
        ELSIF x =- 2456 THEN
            exp_f := 618;
        ELSIF x =- 2455 THEN
            exp_f := 618;
        ELSIF x =- 2454 THEN
            exp_f := 618;
        ELSIF x =- 2453 THEN
            exp_f := 618;
        ELSIF x =- 2452 THEN
            exp_f := 618;
        ELSIF x =- 2451 THEN
            exp_f := 620;
        ELSIF x =- 2450 THEN
            exp_f := 620;
        ELSIF x =- 2449 THEN
            exp_f := 620;
        ELSIF x =- 2448 THEN
            exp_f := 620;
        ELSIF x =- 2447 THEN
            exp_f := 620;
        ELSIF x =- 2446 THEN
            exp_f := 620;
        ELSIF x =- 2445 THEN
            exp_f := 621;
        ELSIF x =- 2444 THEN
            exp_f := 621;
        ELSIF x =- 2443 THEN
            exp_f := 621;
        ELSIF x =- 2442 THEN
            exp_f := 621;
        ELSIF x =- 2441 THEN
            exp_f := 621;
        ELSIF x =- 2440 THEN
            exp_f := 623;
        ELSIF x =- 2439 THEN
            exp_f := 623;
        ELSIF x =- 2438 THEN
            exp_f := 623;
        ELSIF x =- 2437 THEN
            exp_f := 623;
        ELSIF x =- 2436 THEN
            exp_f := 623;
        ELSIF x =- 2435 THEN
            exp_f := 625;
        ELSIF x =- 2434 THEN
            exp_f := 625;
        ELSIF x =- 2433 THEN
            exp_f := 625;
        ELSIF x =- 2432 THEN
            exp_f := 625;
        ELSIF x =- 2431 THEN
            exp_f := 625;
        ELSIF x =- 2430 THEN
            exp_f := 625;
        ELSIF x =- 2429 THEN
            exp_f := 626;
        ELSIF x =- 2428 THEN
            exp_f := 626;
        ELSIF x =- 2427 THEN
            exp_f := 626;
        ELSIF x =- 2426 THEN
            exp_f := 626;
        ELSIF x =- 2425 THEN
            exp_f := 626;
        ELSIF x =- 2424 THEN
            exp_f := 628;
        ELSIF x =- 2423 THEN
            exp_f := 628;
        ELSIF x =- 2422 THEN
            exp_f := 628;
        ELSIF x =- 2421 THEN
            exp_f := 628;
        ELSIF x =- 2420 THEN
            exp_f := 628;
        ELSIF x =- 2419 THEN
            exp_f := 628;
        ELSIF x =- 2418 THEN
            exp_f := 630;
        ELSIF x =- 2417 THEN
            exp_f := 630;
        ELSIF x =- 2416 THEN
            exp_f := 630;
        ELSIF x =- 2415 THEN
            exp_f := 630;
        ELSIF x =- 2414 THEN
            exp_f := 630;
        ELSIF x =- 2413 THEN
            exp_f := 632;
        ELSIF x =- 2412 THEN
            exp_f := 632;
        ELSIF x =- 2411 THEN
            exp_f := 632;
        ELSIF x =- 2410 THEN
            exp_f := 632;
        ELSIF x =- 2409 THEN
            exp_f := 632;
        ELSIF x =- 2408 THEN
            exp_f := 633;
        ELSIF x =- 2407 THEN
            exp_f := 633;
        ELSIF x =- 2406 THEN
            exp_f := 633;
        ELSIF x =- 2405 THEN
            exp_f := 633;
        ELSIF x =- 2404 THEN
            exp_f := 633;
        ELSIF x =- 2403 THEN
            exp_f := 633;
        ELSIF x =- 2402 THEN
            exp_f := 635;
        ELSIF x =- 2401 THEN
            exp_f := 635;
        ELSIF x =- 2400 THEN
            exp_f := 635;
        ELSIF x =- 2399 THEN
            exp_f := 635;
        ELSIF x =- 2398 THEN
            exp_f := 635;
        ELSIF x =- 2397 THEN
            exp_f := 637;
        ELSIF x =- 2396 THEN
            exp_f := 637;
        ELSIF x =- 2395 THEN
            exp_f := 637;
        ELSIF x =- 2394 THEN
            exp_f := 637;
        ELSIF x =- 2393 THEN
            exp_f := 637;
        ELSIF x =- 2392 THEN
            exp_f := 638;
        ELSIF x =- 2391 THEN
            exp_f := 638;
        ELSIF x =- 2390 THEN
            exp_f := 638;
        ELSIF x =- 2389 THEN
            exp_f := 638;
        ELSIF x =- 2388 THEN
            exp_f := 638;
        ELSIF x =- 2387 THEN
            exp_f := 638;
        ELSIF x =- 2386 THEN
            exp_f := 640;
        ELSIF x =- 2385 THEN
            exp_f := 640;
        ELSIF x =- 2384 THEN
            exp_f := 640;
        ELSIF x =- 2383 THEN
            exp_f := 640;
        ELSIF x =- 2382 THEN
            exp_f := 640;
        ELSIF x =- 2381 THEN
            exp_f := 642;
        ELSIF x =- 2380 THEN
            exp_f := 642;
        ELSIF x =- 2379 THEN
            exp_f := 642;
        ELSIF x =- 2378 THEN
            exp_f := 642;
        ELSIF x =- 2377 THEN
            exp_f := 642;
        ELSIF x =- 2376 THEN
            exp_f := 642;
        ELSIF x =- 2375 THEN
            exp_f := 644;
        ELSIF x =- 2374 THEN
            exp_f := 644;
        ELSIF x =- 2373 THEN
            exp_f := 644;
        ELSIF x =- 2372 THEN
            exp_f := 644;
        ELSIF x =- 2371 THEN
            exp_f := 644;
        ELSIF x =- 2370 THEN
            exp_f := 645;
        ELSIF x =- 2369 THEN
            exp_f := 645;
        ELSIF x =- 2368 THEN
            exp_f := 645;
        ELSIF x =- 2367 THEN
            exp_f := 645;
        ELSIF x =- 2366 THEN
            exp_f := 645;
        ELSIF x =- 2365 THEN
            exp_f := 647;
        ELSIF x =- 2364 THEN
            exp_f := 647;
        ELSIF x =- 2363 THEN
            exp_f := 647;
        ELSIF x =- 2362 THEN
            exp_f := 647;
        ELSIF x =- 2361 THEN
            exp_f := 647;
        ELSIF x =- 2360 THEN
            exp_f := 647;
        ELSIF x =- 2359 THEN
            exp_f := 649;
        ELSIF x =- 2358 THEN
            exp_f := 649;
        ELSIF x =- 2357 THEN
            exp_f := 649;
        ELSIF x =- 2356 THEN
            exp_f := 649;
        ELSIF x =- 2355 THEN
            exp_f := 649;
        ELSIF x =- 2354 THEN
            exp_f := 651;
        ELSIF x =- 2353 THEN
            exp_f := 651;
        ELSIF x =- 2352 THEN
            exp_f := 651;
        ELSIF x =- 2351 THEN
            exp_f := 651;
        ELSIF x =- 2350 THEN
            exp_f := 651;
        ELSIF x =- 2349 THEN
            exp_f := 652;
        ELSIF x =- 2348 THEN
            exp_f := 652;
        ELSIF x =- 2347 THEN
            exp_f := 652;
        ELSIF x =- 2346 THEN
            exp_f := 652;
        ELSIF x =- 2345 THEN
            exp_f := 652;
        ELSIF x =- 2344 THEN
            exp_f := 652;
        ELSIF x =- 2343 THEN
            exp_f := 654;
        ELSIF x =- 2342 THEN
            exp_f := 654;
        ELSIF x =- 2341 THEN
            exp_f := 654;
        ELSIF x =- 2340 THEN
            exp_f := 654;
        ELSIF x =- 2339 THEN
            exp_f := 654;
        ELSIF x =- 2338 THEN
            exp_f := 656;
        ELSIF x =- 2337 THEN
            exp_f := 656;
        ELSIF x =- 2336 THEN
            exp_f := 656;
        ELSIF x =- 2335 THEN
            exp_f := 656;
        ELSIF x =- 2334 THEN
            exp_f := 656;
        ELSIF x =- 2333 THEN
            exp_f := 656;
        ELSIF x =- 2332 THEN
            exp_f := 658;
        ELSIF x =- 2331 THEN
            exp_f := 658;
        ELSIF x =- 2330 THEN
            exp_f := 658;
        ELSIF x =- 2329 THEN
            exp_f := 658;
        ELSIF x =- 2328 THEN
            exp_f := 658;
        ELSIF x =- 2327 THEN
            exp_f := 659;
        ELSIF x =- 2326 THEN
            exp_f := 659;
        ELSIF x =- 2325 THEN
            exp_f := 659;
        ELSIF x =- 2324 THEN
            exp_f := 659;
        ELSIF x =- 2323 THEN
            exp_f := 659;
        ELSIF x =- 2322 THEN
            exp_f := 661;
        ELSIF x =- 2321 THEN
            exp_f := 661;
        ELSIF x =- 2320 THEN
            exp_f := 661;
        ELSIF x =- 2319 THEN
            exp_f := 661;
        ELSIF x =- 2318 THEN
            exp_f := 661;
        ELSIF x =- 2317 THEN
            exp_f := 661;
        ELSIF x =- 2316 THEN
            exp_f := 663;
        ELSIF x =- 2315 THEN
            exp_f := 663;
        ELSIF x =- 2314 THEN
            exp_f := 663;
        ELSIF x =- 2313 THEN
            exp_f := 663;
        ELSIF x =- 2312 THEN
            exp_f := 663;
        ELSIF x =- 2311 THEN
            exp_f := 665;
        ELSIF x =- 2310 THEN
            exp_f := 665;
        ELSIF x =- 2309 THEN
            exp_f := 665;
        ELSIF x =- 2308 THEN
            exp_f := 665;
        ELSIF x =- 2307 THEN
            exp_f := 665;
        ELSIF x =- 2306 THEN
            exp_f := 666;
        ELSIF x =- 2305 THEN
            exp_f := 666;
        ELSIF x =- 2304 THEN
            exp_f := 666;
        ELSIF x =- 2303 THEN
            exp_f := 666;
        ELSIF x =- 2302 THEN
            exp_f := 666;
        ELSIF x =- 2301 THEN
            exp_f := 666;
        ELSIF x =- 2300 THEN
            exp_f := 668;
        ELSIF x =- 2299 THEN
            exp_f := 668;
        ELSIF x =- 2298 THEN
            exp_f := 668;
        ELSIF x =- 2297 THEN
            exp_f := 668;
        ELSIF x =- 2296 THEN
            exp_f := 668;
        ELSIF x =- 2295 THEN
            exp_f := 670;
        ELSIF x =- 2294 THEN
            exp_f := 670;
        ELSIF x =- 2293 THEN
            exp_f := 670;
        ELSIF x =- 2292 THEN
            exp_f := 670;
        ELSIF x =- 2291 THEN
            exp_f := 670;
        ELSIF x =- 2290 THEN
            exp_f := 670;
        ELSIF x =- 2289 THEN
            exp_f := 672;
        ELSIF x =- 2288 THEN
            exp_f := 672;
        ELSIF x =- 2287 THEN
            exp_f := 672;
        ELSIF x =- 2286 THEN
            exp_f := 672;
        ELSIF x =- 2285 THEN
            exp_f := 672;
        ELSIF x =- 2284 THEN
            exp_f := 673;
        ELSIF x =- 2283 THEN
            exp_f := 673;
        ELSIF x =- 2282 THEN
            exp_f := 673;
        ELSIF x =- 2281 THEN
            exp_f := 673;
        ELSIF x =- 2280 THEN
            exp_f := 673;
        ELSIF x =- 2279 THEN
            exp_f := 675;
        ELSIF x =- 2278 THEN
            exp_f := 675;
        ELSIF x =- 2277 THEN
            exp_f := 675;
        ELSIF x =- 2276 THEN
            exp_f := 675;
        ELSIF x =- 2275 THEN
            exp_f := 675;
        ELSIF x =- 2274 THEN
            exp_f := 675;
        ELSIF x =- 2273 THEN
            exp_f := 677;
        ELSIF x =- 2272 THEN
            exp_f := 677;
        ELSIF x =- 2271 THEN
            exp_f := 677;
        ELSIF x =- 2270 THEN
            exp_f := 677;
        ELSIF x =- 2269 THEN
            exp_f := 677;
        ELSIF x =- 2268 THEN
            exp_f := 679;
        ELSIF x =- 2267 THEN
            exp_f := 679;
        ELSIF x =- 2266 THEN
            exp_f := 679;
        ELSIF x =- 2265 THEN
            exp_f := 679;
        ELSIF x =- 2264 THEN
            exp_f := 679;
        ELSIF x =- 2263 THEN
            exp_f := 680;
        ELSIF x =- 2262 THEN
            exp_f := 680;
        ELSIF x =- 2261 THEN
            exp_f := 680;
        ELSIF x =- 2260 THEN
            exp_f := 680;
        ELSIF x =- 2259 THEN
            exp_f := 680;
        ELSIF x =- 2258 THEN
            exp_f := 680;
        ELSIF x =- 2257 THEN
            exp_f := 682;
        ELSIF x =- 2256 THEN
            exp_f := 682;
        ELSIF x =- 2255 THEN
            exp_f := 682;
        ELSIF x =- 2254 THEN
            exp_f := 682;
        ELSIF x =- 2253 THEN
            exp_f := 682;
        ELSIF x =- 2252 THEN
            exp_f := 684;
        ELSIF x =- 2251 THEN
            exp_f := 684;
        ELSIF x =- 2250 THEN
            exp_f := 684;
        ELSIF x =- 2249 THEN
            exp_f := 684;
        ELSIF x =- 2248 THEN
            exp_f := 684;
        ELSIF x =- 2247 THEN
            exp_f := 684;
        ELSIF x =- 2246 THEN
            exp_f := 686;
        ELSIF x =- 2245 THEN
            exp_f := 686;
        ELSIF x =- 2244 THEN
            exp_f := 686;
        ELSIF x =- 2243 THEN
            exp_f := 686;
        ELSIF x =- 2242 THEN
            exp_f := 686;
        ELSIF x =- 2241 THEN
            exp_f := 688;
        ELSIF x =- 2240 THEN
            exp_f := 688;
        ELSIF x =- 2239 THEN
            exp_f := 688;
        ELSIF x =- 2238 THEN
            exp_f := 688;
        ELSIF x =- 2237 THEN
            exp_f := 688;
        ELSIF x =- 2236 THEN
            exp_f := 689;
        ELSIF x =- 2235 THEN
            exp_f := 689;
        ELSIF x =- 2234 THEN
            exp_f := 689;
        ELSIF x =- 2233 THEN
            exp_f := 689;
        ELSIF x =- 2232 THEN
            exp_f := 689;
        ELSIF x =- 2231 THEN
            exp_f := 689;
        ELSIF x =- 2230 THEN
            exp_f := 691;
        ELSIF x =- 2229 THEN
            exp_f := 691;
        ELSIF x =- 2228 THEN
            exp_f := 691;
        ELSIF x =- 2227 THEN
            exp_f := 691;
        ELSIF x =- 2226 THEN
            exp_f := 691;
        ELSIF x =- 2225 THEN
            exp_f := 693;
        ELSIF x =- 2224 THEN
            exp_f := 693;
        ELSIF x =- 2223 THEN
            exp_f := 693;
        ELSIF x =- 2222 THEN
            exp_f := 693;
        ELSIF x =- 2221 THEN
            exp_f := 693;
        ELSIF x =- 2220 THEN
            exp_f := 695;
        ELSIF x =- 2219 THEN
            exp_f := 695;
        ELSIF x =- 2218 THEN
            exp_f := 695;
        ELSIF x =- 2217 THEN
            exp_f := 695;
        ELSIF x =- 2216 THEN
            exp_f := 695;
        ELSIF x =- 2215 THEN
            exp_f := 695;
        ELSIF x =- 2214 THEN
            exp_f := 696;
        ELSIF x =- 2213 THEN
            exp_f := 696;
        ELSIF x =- 2212 THEN
            exp_f := 696;
        ELSIF x =- 2211 THEN
            exp_f := 696;
        ELSIF x =- 2210 THEN
            exp_f := 696;
        ELSIF x =- 2209 THEN
            exp_f := 698;
        ELSIF x =- 2208 THEN
            exp_f := 698;
        ELSIF x =- 2207 THEN
            exp_f := 698;
        ELSIF x =- 2206 THEN
            exp_f := 698;
        ELSIF x =- 2205 THEN
            exp_f := 698;
        ELSIF x =- 2204 THEN
            exp_f := 698;
        ELSIF x =- 2203 THEN
            exp_f := 700;
        ELSIF x =- 2202 THEN
            exp_f := 700;
        ELSIF x =- 2201 THEN
            exp_f := 700;
        ELSIF x =- 2200 THEN
            exp_f := 700;
        ELSIF x =- 2199 THEN
            exp_f := 700;
        ELSIF x =- 2198 THEN
            exp_f := 702;
        ELSIF x =- 2197 THEN
            exp_f := 702;
        ELSIF x =- 2196 THEN
            exp_f := 702;
        ELSIF x =- 2195 THEN
            exp_f := 702;
        ELSIF x =- 2194 THEN
            exp_f := 702;
        ELSIF x =- 2193 THEN
            exp_f := 704;
        ELSIF x =- 2192 THEN
            exp_f := 704;
        ELSIF x =- 2191 THEN
            exp_f := 704;
        ELSIF x =- 2190 THEN
            exp_f := 704;
        ELSIF x =- 2189 THEN
            exp_f := 704;
        ELSIF x =- 2188 THEN
            exp_f := 704;
        ELSIF x =- 2187 THEN
            exp_f := 705;
        ELSIF x =- 2186 THEN
            exp_f := 705;
        ELSIF x =- 2185 THEN
            exp_f := 705;
        ELSIF x =- 2184 THEN
            exp_f := 705;
        ELSIF x =- 2183 THEN
            exp_f := 705;
        ELSIF x =- 2182 THEN
            exp_f := 707;
        ELSIF x =- 2181 THEN
            exp_f := 707;
        ELSIF x =- 2180 THEN
            exp_f := 707;
        ELSIF x =- 2179 THEN
            exp_f := 707;
        ELSIF x =- 2178 THEN
            exp_f := 707;
        ELSIF x =- 2177 THEN
            exp_f := 709;
        ELSIF x =- 2176 THEN
            exp_f := 709;
        ELSIF x =- 2175 THEN
            exp_f := 709;
        ELSIF x =- 2174 THEN
            exp_f := 709;
        ELSIF x =- 2173 THEN
            exp_f := 709;
        ELSIF x =- 2172 THEN
            exp_f := 709;
        ELSIF x =- 2171 THEN
            exp_f := 711;
        ELSIF x =- 2170 THEN
            exp_f := 711;
        ELSIF x =- 2169 THEN
            exp_f := 711;
        ELSIF x =- 2168 THEN
            exp_f := 711;
        ELSIF x =- 2167 THEN
            exp_f := 711;
        ELSIF x =- 2166 THEN
            exp_f := 713;
        ELSIF x =- 2165 THEN
            exp_f := 713;
        ELSIF x =- 2164 THEN
            exp_f := 713;
        ELSIF x =- 2163 THEN
            exp_f := 713;
        ELSIF x =- 2162 THEN
            exp_f := 713;
        ELSIF x =- 2161 THEN
            exp_f := 713;
        ELSIF x =- 2160 THEN
            exp_f := 715;
        ELSIF x =- 2159 THEN
            exp_f := 715;
        ELSIF x =- 2158 THEN
            exp_f := 715;
        ELSIF x =- 2157 THEN
            exp_f := 715;
        ELSIF x =- 2156 THEN
            exp_f := 715;
        ELSIF x =- 2155 THEN
            exp_f := 716;
        ELSIF x =- 2154 THEN
            exp_f := 716;
        ELSIF x =- 2153 THEN
            exp_f := 716;
        ELSIF x =- 2152 THEN
            exp_f := 716;
        ELSIF x =- 2151 THEN
            exp_f := 716;
        ELSIF x =- 2150 THEN
            exp_f := 718;
        ELSIF x =- 2149 THEN
            exp_f := 718;
        ELSIF x =- 2148 THEN
            exp_f := 718;
        ELSIF x =- 2147 THEN
            exp_f := 718;
        ELSIF x =- 2146 THEN
            exp_f := 718;
        ELSIF x =- 2145 THEN
            exp_f := 718;
        ELSIF x =- 2144 THEN
            exp_f := 720;
        ELSIF x =- 2143 THEN
            exp_f := 720;
        ELSIF x =- 2142 THEN
            exp_f := 720;
        ELSIF x =- 2141 THEN
            exp_f := 720;
        ELSIF x =- 2140 THEN
            exp_f := 720;
        ELSIF x =- 2139 THEN
            exp_f := 722;
        ELSIF x =- 2138 THEN
            exp_f := 722;
        ELSIF x =- 2137 THEN
            exp_f := 722;
        ELSIF x =- 2136 THEN
            exp_f := 722;
        ELSIF x =- 2135 THEN
            exp_f := 722;
        ELSIF x =- 2134 THEN
            exp_f := 724;
        ELSIF x =- 2133 THEN
            exp_f := 724;
        ELSIF x =- 2132 THEN
            exp_f := 724;
        ELSIF x =- 2131 THEN
            exp_f := 724;
        ELSIF x =- 2130 THEN
            exp_f := 724;
        ELSIF x =- 2129 THEN
            exp_f := 724;
        ELSIF x =- 2128 THEN
            exp_f := 726;
        ELSIF x =- 2127 THEN
            exp_f := 726;
        ELSIF x =- 2126 THEN
            exp_f := 726;
        ELSIF x =- 2125 THEN
            exp_f := 726;
        ELSIF x =- 2124 THEN
            exp_f := 726;
        ELSIF x =- 2123 THEN
            exp_f := 727;
        ELSIF x =- 2122 THEN
            exp_f := 727;
        ELSIF x =- 2121 THEN
            exp_f := 727;
        ELSIF x =- 2120 THEN
            exp_f := 727;
        ELSIF x =- 2119 THEN
            exp_f := 727;
        ELSIF x =- 2118 THEN
            exp_f := 727;
        ELSIF x =- 2117 THEN
            exp_f := 729;
        ELSIF x =- 2116 THEN
            exp_f := 729;
        ELSIF x =- 2115 THEN
            exp_f := 729;
        ELSIF x =- 2114 THEN
            exp_f := 729;
        ELSIF x =- 2113 THEN
            exp_f := 729;
        ELSIF x =- 2112 THEN
            exp_f := 731;
        ELSIF x =- 2111 THEN
            exp_f := 731;
        ELSIF x =- 2110 THEN
            exp_f := 731;
        ELSIF x =- 2109 THEN
            exp_f := 731;
        ELSIF x =- 2108 THEN
            exp_f := 731;
        ELSIF x =- 2107 THEN
            exp_f := 733;
        ELSIF x =- 2106 THEN
            exp_f := 733;
        ELSIF x =- 2105 THEN
            exp_f := 733;
        ELSIF x =- 2104 THEN
            exp_f := 733;
        ELSIF x =- 2103 THEN
            exp_f := 733;
        ELSIF x =- 2102 THEN
            exp_f := 733;
        ELSIF x =- 2101 THEN
            exp_f := 735;
        ELSIF x =- 2100 THEN
            exp_f := 735;
        ELSIF x =- 2099 THEN
            exp_f := 735;
        ELSIF x =- 2098 THEN
            exp_f := 735;
        ELSIF x =- 2097 THEN
            exp_f := 735;
        ELSIF x =- 2096 THEN
            exp_f := 737;
        ELSIF x =- 2095 THEN
            exp_f := 737;
        ELSIF x =- 2094 THEN
            exp_f := 737;
        ELSIF x =- 2093 THEN
            exp_f := 737;
        ELSIF x =- 2092 THEN
            exp_f := 737;
        ELSIF x =- 2091 THEN
            exp_f := 738;
        ELSIF x =- 2090 THEN
            exp_f := 738;
        ELSIF x =- 2089 THEN
            exp_f := 738;
        ELSIF x =- 2088 THEN
            exp_f := 738;
        ELSIF x =- 2087 THEN
            exp_f := 738;
        ELSIF x =- 2086 THEN
            exp_f := 738;
        ELSIF x =- 2085 THEN
            exp_f := 740;
        ELSIF x =- 2084 THEN
            exp_f := 740;
        ELSIF x =- 2083 THEN
            exp_f := 740;
        ELSIF x =- 2082 THEN
            exp_f := 740;
        ELSIF x =- 2081 THEN
            exp_f := 740;
        ELSIF x =- 2080 THEN
            exp_f := 742;
        ELSIF x =- 2079 THEN
            exp_f := 742;
        ELSIF x =- 2078 THEN
            exp_f := 742;
        ELSIF x =- 2077 THEN
            exp_f := 742;
        ELSIF x =- 2076 THEN
            exp_f := 742;
        ELSIF x =- 2075 THEN
            exp_f := 742;
        ELSIF x =- 2074 THEN
            exp_f := 744;
        ELSIF x =- 2073 THEN
            exp_f := 744;
        ELSIF x =- 2072 THEN
            exp_f := 744;
        ELSIF x =- 2071 THEN
            exp_f := 744;
        ELSIF x =- 2070 THEN
            exp_f := 744;
        ELSIF x =- 2069 THEN
            exp_f := 746;
        ELSIF x =- 2068 THEN
            exp_f := 746;
        ELSIF x =- 2067 THEN
            exp_f := 746;
        ELSIF x =- 2066 THEN
            exp_f := 746;
        ELSIF x =- 2065 THEN
            exp_f := 746;
        ELSIF x =- 2064 THEN
            exp_f := 748;
        ELSIF x =- 2063 THEN
            exp_f := 748;
        ELSIF x =- 2062 THEN
            exp_f := 748;
        ELSIF x =- 2061 THEN
            exp_f := 748;
        ELSIF x =- 2060 THEN
            exp_f := 748;
        ELSIF x =- 2059 THEN
            exp_f := 748;
        ELSIF x =- 2058 THEN
            exp_f := 750;
        ELSIF x =- 2057 THEN
            exp_f := 750;
        ELSIF x =- 2056 THEN
            exp_f := 750;
        ELSIF x =- 2055 THEN
            exp_f := 750;
        ELSIF x =- 2054 THEN
            exp_f := 750;
        ELSIF x =- 2053 THEN
            exp_f := 751;
        ELSIF x =- 2052 THEN
            exp_f := 751;
        ELSIF x =- 2051 THEN
            exp_f := 751;
        ELSIF x =- 2050 THEN
            exp_f := 751;
        ELSIF x =- 2049 THEN
            exp_f := 751;
        ELSIF x =- 2048 THEN
            exp_f := 751;
        ELSIF x =- 2047 THEN
            exp_f := 753;
        ELSIF x =- 2046 THEN
            exp_f := 753;
        ELSIF x =- 2045 THEN
            exp_f := 753;
        ELSIF x =- 2044 THEN
            exp_f := 753;
        ELSIF x =- 2043 THEN
            exp_f := 755;
        ELSIF x =- 2042 THEN
            exp_f := 755;
        ELSIF x =- 2041 THEN
            exp_f := 755;
        ELSIF x =- 2040 THEN
            exp_f := 755;
        ELSIF x =- 2039 THEN
            exp_f := 755;
        ELSIF x =- 2038 THEN
            exp_f := 757;
        ELSIF x =- 2037 THEN
            exp_f := 757;
        ELSIF x =- 2036 THEN
            exp_f := 757;
        ELSIF x =- 2035 THEN
            exp_f := 757;
        ELSIF x =- 2034 THEN
            exp_f := 757;
        ELSIF x =- 2033 THEN
            exp_f := 759;
        ELSIF x =- 2032 THEN
            exp_f := 759;
        ELSIF x =- 2031 THEN
            exp_f := 759;
        ELSIF x =- 2030 THEN
            exp_f := 759;
        ELSIF x =- 2029 THEN
            exp_f := 759;
        ELSIF x =- 2028 THEN
            exp_f := 761;
        ELSIF x =- 2027 THEN
            exp_f := 761;
        ELSIF x =- 2026 THEN
            exp_f := 761;
        ELSIF x =- 2025 THEN
            exp_f := 761;
        ELSIF x =- 2024 THEN
            exp_f := 761;
        ELSIF x =- 2023 THEN
            exp_f := 763;
        ELSIF x =- 2022 THEN
            exp_f := 763;
        ELSIF x =- 2021 THEN
            exp_f := 763;
        ELSIF x =- 2020 THEN
            exp_f := 763;
        ELSIF x =- 2019 THEN
            exp_f := 765;
        ELSIF x =- 2018 THEN
            exp_f := 765;
        ELSIF x =- 2017 THEN
            exp_f := 765;
        ELSIF x =- 2016 THEN
            exp_f := 765;
        ELSIF x =- 2015 THEN
            exp_f := 765;
        ELSIF x =- 2014 THEN
            exp_f := 766;
        ELSIF x =- 2013 THEN
            exp_f := 766;
        ELSIF x =- 2012 THEN
            exp_f := 766;
        ELSIF x =- 2011 THEN
            exp_f := 766;
        ELSIF x =- 2010 THEN
            exp_f := 766;
        ELSIF x =- 2009 THEN
            exp_f := 768;
        ELSIF x =- 2008 THEN
            exp_f := 768;
        ELSIF x =- 2007 THEN
            exp_f := 768;
        ELSIF x =- 2006 THEN
            exp_f := 768;
        ELSIF x =- 2005 THEN
            exp_f := 768;
        ELSIF x =- 2004 THEN
            exp_f := 770;
        ELSIF x =- 2003 THEN
            exp_f := 770;
        ELSIF x =- 2002 THEN
            exp_f := 770;
        ELSIF x =- 2001 THEN
            exp_f := 770;
        ELSIF x =- 2000 THEN
            exp_f := 770;
        ELSIF x =- 1999 THEN
            exp_f := 772;
        ELSIF x =- 1998 THEN
            exp_f := 772;
        ELSIF x =- 1997 THEN
            exp_f := 772;
        ELSIF x =- 1996 THEN
            exp_f := 772;
        ELSIF x =- 1995 THEN
            exp_f := 772;
        ELSIF x =- 1994 THEN
            exp_f := 774;
        ELSIF x =- 1993 THEN
            exp_f := 774;
        ELSIF x =- 1992 THEN
            exp_f := 774;
        ELSIF x =- 1991 THEN
            exp_f := 774;
        ELSIF x =- 1990 THEN
            exp_f := 776;
        ELSIF x =- 1989 THEN
            exp_f := 776;
        ELSIF x =- 1988 THEN
            exp_f := 776;
        ELSIF x =- 1987 THEN
            exp_f := 776;
        ELSIF x =- 1986 THEN
            exp_f := 776;
        ELSIF x =- 1985 THEN
            exp_f := 778;
        ELSIF x =- 1984 THEN
            exp_f := 778;
        ELSIF x =- 1983 THEN
            exp_f := 778;
        ELSIF x =- 1982 THEN
            exp_f := 778;
        ELSIF x =- 1981 THEN
            exp_f := 778;
        ELSIF x =- 1980 THEN
            exp_f := 780;
        ELSIF x =- 1979 THEN
            exp_f := 780;
        ELSIF x =- 1978 THEN
            exp_f := 780;
        ELSIF x =- 1977 THEN
            exp_f := 780;
        ELSIF x =- 1976 THEN
            exp_f := 780;
        ELSIF x =- 1975 THEN
            exp_f := 782;
        ELSIF x =- 1974 THEN
            exp_f := 782;
        ELSIF x =- 1973 THEN
            exp_f := 782;
        ELSIF x =- 1972 THEN
            exp_f := 782;
        ELSIF x =- 1971 THEN
            exp_f := 782;
        ELSIF x =- 1970 THEN
            exp_f := 784;
        ELSIF x =- 1969 THEN
            exp_f := 784;
        ELSIF x =- 1968 THEN
            exp_f := 784;
        ELSIF x =- 1967 THEN
            exp_f := 784;
        ELSIF x =- 1966 THEN
            exp_f := 784;
        ELSIF x =- 1965 THEN
            exp_f := 785;
        ELSIF x =- 1964 THEN
            exp_f := 785;
        ELSIF x =- 1963 THEN
            exp_f := 785;
        ELSIF x =- 1962 THEN
            exp_f := 785;
        ELSIF x =- 1961 THEN
            exp_f := 787;
        ELSIF x =- 1960 THEN
            exp_f := 787;
        ELSIF x =- 1959 THEN
            exp_f := 787;
        ELSIF x =- 1958 THEN
            exp_f := 787;
        ELSIF x =- 1957 THEN
            exp_f := 787;
        ELSIF x =- 1956 THEN
            exp_f := 789;
        ELSIF x =- 1955 THEN
            exp_f := 789;
        ELSIF x =- 1954 THEN
            exp_f := 789;
        ELSIF x =- 1953 THEN
            exp_f := 789;
        ELSIF x =- 1952 THEN
            exp_f := 789;
        ELSIF x =- 1951 THEN
            exp_f := 791;
        ELSIF x =- 1950 THEN
            exp_f := 791;
        ELSIF x =- 1949 THEN
            exp_f := 791;
        ELSIF x =- 1948 THEN
            exp_f := 791;
        ELSIF x =- 1947 THEN
            exp_f := 791;
        ELSIF x =- 1946 THEN
            exp_f := 793;
        ELSIF x =- 1945 THEN
            exp_f := 793;
        ELSIF x =- 1944 THEN
            exp_f := 793;
        ELSIF x =- 1943 THEN
            exp_f := 793;
        ELSIF x =- 1942 THEN
            exp_f := 793;
        ELSIF x =- 1941 THEN
            exp_f := 795;
        ELSIF x =- 1940 THEN
            exp_f := 795;
        ELSIF x =- 1939 THEN
            exp_f := 795;
        ELSIF x =- 1938 THEN
            exp_f := 795;
        ELSIF x =- 1937 THEN
            exp_f := 795;
        ELSIF x =- 1936 THEN
            exp_f := 797;
        ELSIF x =- 1935 THEN
            exp_f := 797;
        ELSIF x =- 1934 THEN
            exp_f := 797;
        ELSIF x =- 1933 THEN
            exp_f := 797;
        ELSIF x =- 1932 THEN
            exp_f := 799;
        ELSIF x =- 1931 THEN
            exp_f := 799;
        ELSIF x =- 1930 THEN
            exp_f := 799;
        ELSIF x =- 1929 THEN
            exp_f := 799;
        ELSIF x =- 1928 THEN
            exp_f := 799;
        ELSIF x =- 1927 THEN
            exp_f := 801;
        ELSIF x =- 1926 THEN
            exp_f := 801;
        ELSIF x =- 1925 THEN
            exp_f := 801;
        ELSIF x =- 1924 THEN
            exp_f := 801;
        ELSIF x =- 1923 THEN
            exp_f := 801;
        ELSIF x =- 1922 THEN
            exp_f := 803;
        ELSIF x =- 1921 THEN
            exp_f := 803;
        ELSIF x =- 1920 THEN
            exp_f := 803;
        ELSIF x =- 1919 THEN
            exp_f := 803;
        ELSIF x =- 1918 THEN
            exp_f := 803;
        ELSIF x =- 1917 THEN
            exp_f := 805;
        ELSIF x =- 1916 THEN
            exp_f := 805;
        ELSIF x =- 1915 THEN
            exp_f := 805;
        ELSIF x =- 1914 THEN
            exp_f := 805;
        ELSIF x =- 1913 THEN
            exp_f := 805;
        ELSIF x =- 1912 THEN
            exp_f := 807;
        ELSIF x =- 1911 THEN
            exp_f := 807;
        ELSIF x =- 1910 THEN
            exp_f := 807;
        ELSIF x =- 1909 THEN
            exp_f := 807;
        ELSIF x =- 1908 THEN
            exp_f := 807;
        ELSIF x =- 1907 THEN
            exp_f := 809;
        ELSIF x =- 1906 THEN
            exp_f := 809;
        ELSIF x =- 1905 THEN
            exp_f := 809;
        ELSIF x =- 1904 THEN
            exp_f := 809;
        ELSIF x =- 1903 THEN
            exp_f := 811;
        ELSIF x =- 1902 THEN
            exp_f := 811;
        ELSIF x =- 1901 THEN
            exp_f := 811;
        ELSIF x =- 1900 THEN
            exp_f := 811;
        ELSIF x =- 1899 THEN
            exp_f := 811;
        ELSIF x =- 1898 THEN
            exp_f := 813;
        ELSIF x =- 1897 THEN
            exp_f := 813;
        ELSIF x =- 1896 THEN
            exp_f := 813;
        ELSIF x =- 1895 THEN
            exp_f := 813;
        ELSIF x =- 1894 THEN
            exp_f := 813;
        ELSIF x =- 1893 THEN
            exp_f := 815;
        ELSIF x =- 1892 THEN
            exp_f := 815;
        ELSIF x =- 1891 THEN
            exp_f := 815;
        ELSIF x =- 1890 THEN
            exp_f := 815;
        ELSIF x =- 1889 THEN
            exp_f := 815;
        ELSIF x =- 1888 THEN
            exp_f := 816;
        ELSIF x =- 1887 THEN
            exp_f := 816;
        ELSIF x =- 1886 THEN
            exp_f := 816;
        ELSIF x =- 1885 THEN
            exp_f := 816;
        ELSIF x =- 1884 THEN
            exp_f := 816;
        ELSIF x =- 1883 THEN
            exp_f := 818;
        ELSIF x =- 1882 THEN
            exp_f := 818;
        ELSIF x =- 1881 THEN
            exp_f := 818;
        ELSIF x =- 1880 THEN
            exp_f := 818;
        ELSIF x =- 1879 THEN
            exp_f := 818;
        ELSIF x =- 1878 THEN
            exp_f := 820;
        ELSIF x =- 1877 THEN
            exp_f := 820;
        ELSIF x =- 1876 THEN
            exp_f := 820;
        ELSIF x =- 1875 THEN
            exp_f := 820;
        ELSIF x =- 1874 THEN
            exp_f := 822;
        ELSIF x =- 1873 THEN
            exp_f := 822;
        ELSIF x =- 1872 THEN
            exp_f := 822;
        ELSIF x =- 1871 THEN
            exp_f := 822;
        ELSIF x =- 1870 THEN
            exp_f := 822;
        ELSIF x =- 1869 THEN
            exp_f := 824;
        ELSIF x =- 1868 THEN
            exp_f := 824;
        ELSIF x =- 1867 THEN
            exp_f := 824;
        ELSIF x =- 1866 THEN
            exp_f := 824;
        ELSIF x =- 1865 THEN
            exp_f := 824;
        ELSIF x =- 1864 THEN
            exp_f := 826;
        ELSIF x =- 1863 THEN
            exp_f := 826;
        ELSIF x =- 1862 THEN
            exp_f := 826;
        ELSIF x =- 1861 THEN
            exp_f := 826;
        ELSIF x =- 1860 THEN
            exp_f := 826;
        ELSIF x =- 1859 THEN
            exp_f := 828;
        ELSIF x =- 1858 THEN
            exp_f := 828;
        ELSIF x =- 1857 THEN
            exp_f := 828;
        ELSIF x =- 1856 THEN
            exp_f := 828;
        ELSIF x =- 1855 THEN
            exp_f := 828;
        ELSIF x =- 1854 THEN
            exp_f := 830;
        ELSIF x =- 1853 THEN
            exp_f := 830;
        ELSIF x =- 1852 THEN
            exp_f := 830;
        ELSIF x =- 1851 THEN
            exp_f := 830;
        ELSIF x =- 1850 THEN
            exp_f := 830;
        ELSIF x =- 1849 THEN
            exp_f := 832;
        ELSIF x =- 1848 THEN
            exp_f := 832;
        ELSIF x =- 1847 THEN
            exp_f := 832;
        ELSIF x =- 1846 THEN
            exp_f := 832;
        ELSIF x =- 1845 THEN
            exp_f := 834;
        ELSIF x =- 1844 THEN
            exp_f := 834;
        ELSIF x =- 1843 THEN
            exp_f := 834;
        ELSIF x =- 1842 THEN
            exp_f := 834;
        ELSIF x =- 1841 THEN
            exp_f := 834;
        ELSIF x =- 1840 THEN
            exp_f := 836;
        ELSIF x =- 1839 THEN
            exp_f := 836;
        ELSIF x =- 1838 THEN
            exp_f := 836;
        ELSIF x =- 1837 THEN
            exp_f := 836;
        ELSIF x =- 1836 THEN
            exp_f := 836;
        ELSIF x =- 1835 THEN
            exp_f := 838;
        ELSIF x =- 1834 THEN
            exp_f := 838;
        ELSIF x =- 1833 THEN
            exp_f := 838;
        ELSIF x =- 1832 THEN
            exp_f := 838;
        ELSIF x =- 1831 THEN
            exp_f := 838;
        ELSIF x =- 1830 THEN
            exp_f := 840;
        ELSIF x =- 1829 THEN
            exp_f := 840;
        ELSIF x =- 1828 THEN
            exp_f := 840;
        ELSIF x =- 1827 THEN
            exp_f := 840;
        ELSIF x =- 1826 THEN
            exp_f := 840;
        ELSIF x =- 1825 THEN
            exp_f := 842;
        ELSIF x =- 1824 THEN
            exp_f := 842;
        ELSIF x =- 1823 THEN
            exp_f := 842;
        ELSIF x =- 1822 THEN
            exp_f := 842;
        ELSIF x =- 1821 THEN
            exp_f := 842;
        ELSIF x =- 1820 THEN
            exp_f := 844;
        ELSIF x =- 1819 THEN
            exp_f := 844;
        ELSIF x =- 1818 THEN
            exp_f := 844;
        ELSIF x =- 1817 THEN
            exp_f := 844;
        ELSIF x =- 1816 THEN
            exp_f := 846;
        ELSIF x =- 1815 THEN
            exp_f := 846;
        ELSIF x =- 1814 THEN
            exp_f := 846;
        ELSIF x =- 1813 THEN
            exp_f := 846;
        ELSIF x =- 1812 THEN
            exp_f := 846;
        ELSIF x =- 1811 THEN
            exp_f := 848;
        ELSIF x =- 1810 THEN
            exp_f := 848;
        ELSIF x =- 1809 THEN
            exp_f := 848;
        ELSIF x =- 1808 THEN
            exp_f := 848;
        ELSIF x =- 1807 THEN
            exp_f := 848;
        ELSIF x =- 1806 THEN
            exp_f := 850;
        ELSIF x =- 1805 THEN
            exp_f := 850;
        ELSIF x =- 1804 THEN
            exp_f := 850;
        ELSIF x =- 1803 THEN
            exp_f := 850;
        ELSIF x =- 1802 THEN
            exp_f := 850;
        ELSIF x =- 1801 THEN
            exp_f := 852;
        ELSIF x =- 1800 THEN
            exp_f := 852;
        ELSIF x =- 1799 THEN
            exp_f := 852;
        ELSIF x =- 1798 THEN
            exp_f := 852;
        ELSIF x =- 1797 THEN
            exp_f := 852;
        ELSIF x =- 1796 THEN
            exp_f := 854;
        ELSIF x =- 1795 THEN
            exp_f := 854;
        ELSIF x =- 1794 THEN
            exp_f := 854;
        ELSIF x =- 1793 THEN
            exp_f := 854;
        ELSIF x =- 1792 THEN
            exp_f := 854;
        ELSIF x =- 1791 THEN
            exp_f := 856;
        ELSIF x =- 1790 THEN
            exp_f := 856;
        ELSIF x =- 1789 THEN
            exp_f := 856;
        ELSIF x =- 1788 THEN
            exp_f := 856;
        ELSIF x =- 1787 THEN
            exp_f := 858;
        ELSIF x =- 1786 THEN
            exp_f := 858;
        ELSIF x =- 1785 THEN
            exp_f := 858;
        ELSIF x =- 1784 THEN
            exp_f := 858;
        ELSIF x =- 1783 THEN
            exp_f := 858;
        ELSIF x =- 1782 THEN
            exp_f := 860;
        ELSIF x =- 1781 THEN
            exp_f := 860;
        ELSIF x =- 1780 THEN
            exp_f := 860;
        ELSIF x =- 1779 THEN
            exp_f := 860;
        ELSIF x =- 1778 THEN
            exp_f := 860;
        ELSIF x =- 1777 THEN
            exp_f := 862;
        ELSIF x =- 1776 THEN
            exp_f := 862;
        ELSIF x =- 1775 THEN
            exp_f := 862;
        ELSIF x =- 1774 THEN
            exp_f := 862;
        ELSIF x =- 1773 THEN
            exp_f := 862;
        ELSIF x =- 1772 THEN
            exp_f := 864;
        ELSIF x =- 1771 THEN
            exp_f := 864;
        ELSIF x =- 1770 THEN
            exp_f := 864;
        ELSIF x =- 1769 THEN
            exp_f := 864;
        ELSIF x =- 1768 THEN
            exp_f := 864;
        ELSIF x =- 1767 THEN
            exp_f := 866;
        ELSIF x =- 1766 THEN
            exp_f := 866;
        ELSIF x =- 1765 THEN
            exp_f := 866;
        ELSIF x =- 1764 THEN
            exp_f := 866;
        ELSIF x =- 1763 THEN
            exp_f := 868;
        ELSIF x =- 1762 THEN
            exp_f := 868;
        ELSIF x =- 1761 THEN
            exp_f := 868;
        ELSIF x =- 1760 THEN
            exp_f := 868;
        ELSIF x =- 1759 THEN
            exp_f := 868;
        ELSIF x =- 1758 THEN
            exp_f := 870;
        ELSIF x =- 1757 THEN
            exp_f := 870;
        ELSIF x =- 1756 THEN
            exp_f := 870;
        ELSIF x =- 1755 THEN
            exp_f := 870;
        ELSIF x =- 1754 THEN
            exp_f := 870;
        ELSIF x =- 1753 THEN
            exp_f := 872;
        ELSIF x =- 1752 THEN
            exp_f := 872;
        ELSIF x =- 1751 THEN
            exp_f := 872;
        ELSIF x =- 1750 THEN
            exp_f := 872;
        ELSIF x =- 1749 THEN
            exp_f := 872;
        ELSIF x =- 1748 THEN
            exp_f := 874;
        ELSIF x =- 1747 THEN
            exp_f := 874;
        ELSIF x =- 1746 THEN
            exp_f := 874;
        ELSIF x =- 1745 THEN
            exp_f := 874;
        ELSIF x =- 1744 THEN
            exp_f := 874;
        ELSIF x =- 1743 THEN
            exp_f := 876;
        ELSIF x =- 1742 THEN
            exp_f := 876;
        ELSIF x =- 1741 THEN
            exp_f := 876;
        ELSIF x =- 1740 THEN
            exp_f := 876;
        ELSIF x =- 1739 THEN
            exp_f := 876;
        ELSIF x =- 1738 THEN
            exp_f := 878;
        ELSIF x =- 1737 THEN
            exp_f := 878;
        ELSIF x =- 1736 THEN
            exp_f := 878;
        ELSIF x =- 1735 THEN
            exp_f := 878;
        ELSIF x =- 1734 THEN
            exp_f := 880;
        ELSIF x =- 1733 THEN
            exp_f := 880;
        ELSIF x =- 1732 THEN
            exp_f := 880;
        ELSIF x =- 1731 THEN
            exp_f := 880;
        ELSIF x =- 1730 THEN
            exp_f := 880;
        ELSIF x =- 1729 THEN
            exp_f := 883;
        ELSIF x =- 1728 THEN
            exp_f := 883;
        ELSIF x =- 1727 THEN
            exp_f := 883;
        ELSIF x =- 1726 THEN
            exp_f := 883;
        ELSIF x =- 1725 THEN
            exp_f := 883;
        ELSIF x =- 1724 THEN
            exp_f := 885;
        ELSIF x =- 1723 THEN
            exp_f := 885;
        ELSIF x =- 1722 THEN
            exp_f := 885;
        ELSIF x =- 1721 THEN
            exp_f := 885;
        ELSIF x =- 1720 THEN
            exp_f := 885;
        ELSIF x =- 1719 THEN
            exp_f := 887;
        ELSIF x =- 1718 THEN
            exp_f := 887;
        ELSIF x =- 1717 THEN
            exp_f := 887;
        ELSIF x =- 1716 THEN
            exp_f := 887;
        ELSIF x =- 1715 THEN
            exp_f := 887;
        ELSIF x =- 1714 THEN
            exp_f := 889;
        ELSIF x =- 1713 THEN
            exp_f := 889;
        ELSIF x =- 1712 THEN
            exp_f := 889;
        ELSIF x =- 1711 THEN
            exp_f := 889;
        ELSIF x =- 1710 THEN
            exp_f := 889;
        ELSIF x =- 1709 THEN
            exp_f := 891;
        ELSIF x =- 1708 THEN
            exp_f := 891;
        ELSIF x =- 1707 THEN
            exp_f := 891;
        ELSIF x =- 1706 THEN
            exp_f := 891;
        ELSIF x =- 1705 THEN
            exp_f := 893;
        ELSIF x =- 1704 THEN
            exp_f := 893;
        ELSIF x =- 1703 THEN
            exp_f := 893;
        ELSIF x =- 1702 THEN
            exp_f := 893;
        ELSIF x =- 1701 THEN
            exp_f := 893;
        ELSIF x =- 1700 THEN
            exp_f := 895;
        ELSIF x =- 1699 THEN
            exp_f := 895;
        ELSIF x =- 1698 THEN
            exp_f := 895;
        ELSIF x =- 1697 THEN
            exp_f := 895;
        ELSIF x =- 1696 THEN
            exp_f := 895;
        ELSIF x =- 1695 THEN
            exp_f := 897;
        ELSIF x =- 1694 THEN
            exp_f := 897;
        ELSIF x =- 1693 THEN
            exp_f := 897;
        ELSIF x =- 1692 THEN
            exp_f := 897;
        ELSIF x =- 1691 THEN
            exp_f := 897;
        ELSIF x =- 1690 THEN
            exp_f := 899;
        ELSIF x =- 1689 THEN
            exp_f := 899;
        ELSIF x =- 1688 THEN
            exp_f := 899;
        ELSIF x =- 1687 THEN
            exp_f := 899;
        ELSIF x =- 1686 THEN
            exp_f := 899;
        ELSIF x =- 1685 THEN
            exp_f := 901;
        ELSIF x =- 1684 THEN
            exp_f := 901;
        ELSIF x =- 1683 THEN
            exp_f := 901;
        ELSIF x =- 1682 THEN
            exp_f := 901;
        ELSIF x =- 1681 THEN
            exp_f := 901;
        ELSIF x =- 1680 THEN
            exp_f := 903;
        ELSIF x =- 1679 THEN
            exp_f := 903;
        ELSIF x =- 1678 THEN
            exp_f := 903;
        ELSIF x =- 1677 THEN
            exp_f := 903;
        ELSIF x =- 1676 THEN
            exp_f := 905;
        ELSIF x =- 1675 THEN
            exp_f := 905;
        ELSIF x =- 1674 THEN
            exp_f := 905;
        ELSIF x =- 1673 THEN
            exp_f := 905;
        ELSIF x =- 1672 THEN
            exp_f := 905;
        ELSIF x =- 1671 THEN
            exp_f := 907;
        ELSIF x =- 1670 THEN
            exp_f := 907;
        ELSIF x =- 1669 THEN
            exp_f := 907;
        ELSIF x =- 1668 THEN
            exp_f := 907;
        ELSIF x =- 1667 THEN
            exp_f := 907;
        ELSIF x =- 1666 THEN
            exp_f := 909;
        ELSIF x =- 1665 THEN
            exp_f := 909;
        ELSIF x =- 1664 THEN
            exp_f := 909;
        ELSIF x =- 1663 THEN
            exp_f := 909;
        ELSIF x =- 1662 THEN
            exp_f := 909;
        ELSIF x =- 1661 THEN
            exp_f := 911;
        ELSIF x =- 1660 THEN
            exp_f := 911;
        ELSIF x =- 1659 THEN
            exp_f := 911;
        ELSIF x =- 1658 THEN
            exp_f := 911;
        ELSIF x =- 1657 THEN
            exp_f := 911;
        ELSIF x =- 1656 THEN
            exp_f := 914;
        ELSIF x =- 1655 THEN
            exp_f := 914;
        ELSIF x =- 1654 THEN
            exp_f := 914;
        ELSIF x =- 1653 THEN
            exp_f := 914;
        ELSIF x =- 1652 THEN
            exp_f := 914;
        ELSIF x =- 1651 THEN
            exp_f := 916;
        ELSIF x =- 1650 THEN
            exp_f := 916;
        ELSIF x =- 1649 THEN
            exp_f := 916;
        ELSIF x =- 1648 THEN
            exp_f := 916;
        ELSIF x =- 1647 THEN
            exp_f := 918;
        ELSIF x =- 1646 THEN
            exp_f := 918;
        ELSIF x =- 1645 THEN
            exp_f := 918;
        ELSIF x =- 1644 THEN
            exp_f := 918;
        ELSIF x =- 1643 THEN
            exp_f := 918;
        ELSIF x =- 1642 THEN
            exp_f := 920;
        ELSIF x =- 1641 THEN
            exp_f := 920;
        ELSIF x =- 1640 THEN
            exp_f := 920;
        ELSIF x =- 1639 THEN
            exp_f := 920;
        ELSIF x =- 1638 THEN
            exp_f := 920;
        ELSIF x =- 1637 THEN
            exp_f := 922;
        ELSIF x =- 1636 THEN
            exp_f := 922;
        ELSIF x =- 1635 THEN
            exp_f := 922;
        ELSIF x =- 1634 THEN
            exp_f := 922;
        ELSIF x =- 1633 THEN
            exp_f := 922;
        ELSIF x =- 1632 THEN
            exp_f := 924;
        ELSIF x =- 1631 THEN
            exp_f := 924;
        ELSIF x =- 1630 THEN
            exp_f := 924;
        ELSIF x =- 1629 THEN
            exp_f := 924;
        ELSIF x =- 1628 THEN
            exp_f := 924;
        ELSIF x =- 1627 THEN
            exp_f := 926;
        ELSIF x =- 1626 THEN
            exp_f := 926;
        ELSIF x =- 1625 THEN
            exp_f := 926;
        ELSIF x =- 1624 THEN
            exp_f := 926;
        ELSIF x =- 1623 THEN
            exp_f := 926;
        ELSIF x =- 1622 THEN
            exp_f := 928;
        ELSIF x =- 1621 THEN
            exp_f := 928;
        ELSIF x =- 1620 THEN
            exp_f := 928;
        ELSIF x =- 1619 THEN
            exp_f := 928;
        ELSIF x =- 1618 THEN
            exp_f := 930;
        ELSIF x =- 1617 THEN
            exp_f := 930;
        ELSIF x =- 1616 THEN
            exp_f := 930;
        ELSIF x =- 1615 THEN
            exp_f := 930;
        ELSIF x =- 1614 THEN
            exp_f := 930;
        ELSIF x =- 1613 THEN
            exp_f := 933;
        ELSIF x =- 1612 THEN
            exp_f := 933;
        ELSIF x =- 1611 THEN
            exp_f := 933;
        ELSIF x =- 1610 THEN
            exp_f := 933;
        ELSIF x =- 1609 THEN
            exp_f := 933;
        ELSIF x =- 1608 THEN
            exp_f := 935;
        ELSIF x =- 1607 THEN
            exp_f := 935;
        ELSIF x =- 1606 THEN
            exp_f := 935;
        ELSIF x =- 1605 THEN
            exp_f := 935;
        ELSIF x =- 1604 THEN
            exp_f := 935;
        ELSIF x =- 1603 THEN
            exp_f := 937;
        ELSIF x =- 1602 THEN
            exp_f := 937;
        ELSIF x =- 1601 THEN
            exp_f := 937;
        ELSIF x =- 1600 THEN
            exp_f := 937;
        ELSIF x =- 1599 THEN
            exp_f := 937;
        ELSIF x =- 1598 THEN
            exp_f := 939;
        ELSIF x =- 1597 THEN
            exp_f := 939;
        ELSIF x =- 1596 THEN
            exp_f := 939;
        ELSIF x =- 1595 THEN
            exp_f := 939;
        ELSIF x =- 1594 THEN
            exp_f := 939;
        ELSIF x =- 1593 THEN
            exp_f := 941;
        ELSIF x =- 1592 THEN
            exp_f := 941;
        ELSIF x =- 1591 THEN
            exp_f := 941;
        ELSIF x =- 1590 THEN
            exp_f := 941;
        ELSIF x =- 1589 THEN
            exp_f := 943;
        ELSIF x =- 1588 THEN
            exp_f := 943;
        ELSIF x =- 1587 THEN
            exp_f := 943;
        ELSIF x =- 1586 THEN
            exp_f := 943;
        ELSIF x =- 1585 THEN
            exp_f := 943;
        ELSIF x =- 1584 THEN
            exp_f := 945;
        ELSIF x =- 1583 THEN
            exp_f := 945;
        ELSIF x =- 1582 THEN
            exp_f := 945;
        ELSIF x =- 1581 THEN
            exp_f := 945;
        ELSIF x =- 1580 THEN
            exp_f := 945;
        ELSIF x =- 1579 THEN
            exp_f := 947;
        ELSIF x =- 1578 THEN
            exp_f := 947;
        ELSIF x =- 1577 THEN
            exp_f := 947;
        ELSIF x =- 1576 THEN
            exp_f := 947;
        ELSIF x =- 1575 THEN
            exp_f := 947;
        ELSIF x =- 1574 THEN
            exp_f := 950;
        ELSIF x =- 1573 THEN
            exp_f := 950;
        ELSIF x =- 1572 THEN
            exp_f := 950;
        ELSIF x =- 1571 THEN
            exp_f := 950;
        ELSIF x =- 1570 THEN
            exp_f := 950;
        ELSIF x =- 1569 THEN
            exp_f := 952;
        ELSIF x =- 1568 THEN
            exp_f := 952;
        ELSIF x =- 1567 THEN
            exp_f := 952;
        ELSIF x =- 1566 THEN
            exp_f := 952;
        ELSIF x =- 1565 THEN
            exp_f := 952;
        ELSIF x =- 1564 THEN
            exp_f := 954;
        ELSIF x =- 1563 THEN
            exp_f := 954;
        ELSIF x =- 1562 THEN
            exp_f := 954;
        ELSIF x =- 1561 THEN
            exp_f := 954;
        ELSIF x =- 1560 THEN
            exp_f := 956;
        ELSIF x =- 1559 THEN
            exp_f := 956;
        ELSIF x =- 1558 THEN
            exp_f := 956;
        ELSIF x =- 1557 THEN
            exp_f := 956;
        ELSIF x =- 1556 THEN
            exp_f := 956;
        ELSIF x =- 1555 THEN
            exp_f := 958;
        ELSIF x =- 1554 THEN
            exp_f := 958;
        ELSIF x =- 1553 THEN
            exp_f := 958;
        ELSIF x =- 1552 THEN
            exp_f := 958;
        ELSIF x =- 1551 THEN
            exp_f := 958;
        ELSIF x =- 1550 THEN
            exp_f := 960;
        ELSIF x =- 1549 THEN
            exp_f := 960;
        ELSIF x =- 1548 THEN
            exp_f := 960;
        ELSIF x =- 1547 THEN
            exp_f := 960;
        ELSIF x =- 1546 THEN
            exp_f := 960;
        ELSIF x =- 1545 THEN
            exp_f := 962;
        ELSIF x =- 1544 THEN
            exp_f := 962;
        ELSIF x =- 1543 THEN
            exp_f := 962;
        ELSIF x =- 1542 THEN
            exp_f := 962;
        ELSIF x =- 1541 THEN
            exp_f := 962;
        ELSIF x =- 1540 THEN
            exp_f := 965;
        ELSIF x =- 1539 THEN
            exp_f := 965;
        ELSIF x =- 1538 THEN
            exp_f := 965;
        ELSIF x =- 1537 THEN
            exp_f := 965;
        ELSIF x =- 1536 THEN
            exp_f := 965;
        ELSIF x =- 1535 THEN
            exp_f := 967;
        ELSIF x =- 1534 THEN
            exp_f := 967;
        ELSIF x =- 1533 THEN
            exp_f := 967;
        ELSIF x =- 1532 THEN
            exp_f := 969;
        ELSIF x =- 1531 THEN
            exp_f := 969;
        ELSIF x =- 1530 THEN
            exp_f := 969;
        ELSIF x =- 1529 THEN
            exp_f := 969;
        ELSIF x =- 1528 THEN
            exp_f := 971;
        ELSIF x =- 1527 THEN
            exp_f := 971;
        ELSIF x =- 1526 THEN
            exp_f := 971;
        ELSIF x =- 1525 THEN
            exp_f := 971;
        ELSIF x =- 1524 THEN
            exp_f := 971;
        ELSIF x =- 1523 THEN
            exp_f := 973;
        ELSIF x =- 1522 THEN
            exp_f := 973;
        ELSIF x =- 1521 THEN
            exp_f := 973;
        ELSIF x =- 1520 THEN
            exp_f := 973;
        ELSIF x =- 1519 THEN
            exp_f := 976;
        ELSIF x =- 1518 THEN
            exp_f := 976;
        ELSIF x =- 1517 THEN
            exp_f := 976;
        ELSIF x =- 1516 THEN
            exp_f := 976;
        ELSIF x =- 1515 THEN
            exp_f := 978;
        ELSIF x =- 1514 THEN
            exp_f := 978;
        ELSIF x =- 1513 THEN
            exp_f := 978;
        ELSIF x =- 1512 THEN
            exp_f := 978;
        ELSIF x =- 1511 THEN
            exp_f := 978;
        ELSIF x =- 1510 THEN
            exp_f := 980;
        ELSIF x =- 1509 THEN
            exp_f := 980;
        ELSIF x =- 1508 THEN
            exp_f := 980;
        ELSIF x =- 1507 THEN
            exp_f := 980;
        ELSIF x =- 1506 THEN
            exp_f := 982;
        ELSIF x =- 1505 THEN
            exp_f := 982;
        ELSIF x =- 1504 THEN
            exp_f := 982;
        ELSIF x =- 1503 THEN
            exp_f := 982;
        ELSIF x =- 1502 THEN
            exp_f := 982;
        ELSIF x =- 1501 THEN
            exp_f := 984;
        ELSIF x =- 1500 THEN
            exp_f := 984;
        ELSIF x =- 1499 THEN
            exp_f := 984;
        ELSIF x =- 1498 THEN
            exp_f := 984;
        ELSIF x =- 1497 THEN
            exp_f := 986;
        ELSIF x =- 1496 THEN
            exp_f := 986;
        ELSIF x =- 1495 THEN
            exp_f := 986;
        ELSIF x =- 1494 THEN
            exp_f := 986;
        ELSIF x =- 1493 THEN
            exp_f := 989;
        ELSIF x =- 1492 THEN
            exp_f := 989;
        ELSIF x =- 1491 THEN
            exp_f := 989;
        ELSIF x =- 1490 THEN
            exp_f := 989;
        ELSIF x =- 1489 THEN
            exp_f := 989;
        ELSIF x =- 1488 THEN
            exp_f := 991;
        ELSIF x =- 1487 THEN
            exp_f := 991;
        ELSIF x =- 1486 THEN
            exp_f := 991;
        ELSIF x =- 1485 THEN
            exp_f := 991;
        ELSIF x =- 1484 THEN
            exp_f := 993;
        ELSIF x =- 1483 THEN
            exp_f := 993;
        ELSIF x =- 1482 THEN
            exp_f := 993;
        ELSIF x =- 1481 THEN
            exp_f := 993;
        ELSIF x =- 1480 THEN
            exp_f := 993;
        ELSIF x =- 1479 THEN
            exp_f := 995;
        ELSIF x =- 1478 THEN
            exp_f := 995;
        ELSIF x =- 1477 THEN
            exp_f := 995;
        ELSIF x =- 1476 THEN
            exp_f := 995;
        ELSIF x =- 1475 THEN
            exp_f := 997;
        ELSIF x =- 1474 THEN
            exp_f := 997;
        ELSIF x =- 1473 THEN
            exp_f := 997;
        ELSIF x =- 1472 THEN
            exp_f := 997;
        ELSIF x =- 1471 THEN
            exp_f := 1000;
        ELSIF x =- 1470 THEN
            exp_f := 1000;
        ELSIF x =- 1469 THEN
            exp_f := 1000;
        ELSIF x =- 1468 THEN
            exp_f := 1000;
        ELSIF x =- 1467 THEN
            exp_f := 1000;
        ELSIF x =- 1466 THEN
            exp_f := 1002;
        ELSIF x =- 1465 THEN
            exp_f := 1002;
        ELSIF x =- 1464 THEN
            exp_f := 1002;
        ELSIF x =- 1463 THEN
            exp_f := 1002;
        ELSIF x =- 1462 THEN
            exp_f := 1004;
        ELSIF x =- 1461 THEN
            exp_f := 1004;
        ELSIF x =- 1460 THEN
            exp_f := 1004;
        ELSIF x =- 1459 THEN
            exp_f := 1004;
        ELSIF x =- 1458 THEN
            exp_f := 1004;
        ELSIF x =- 1457 THEN
            exp_f := 1006;
        ELSIF x =- 1456 THEN
            exp_f := 1006;
        ELSIF x =- 1455 THEN
            exp_f := 1006;
        ELSIF x =- 1454 THEN
            exp_f := 1006;
        ELSIF x =- 1453 THEN
            exp_f := 1009;
        ELSIF x =- 1452 THEN
            exp_f := 1009;
        ELSIF x =- 1451 THEN
            exp_f := 1009;
        ELSIF x =- 1450 THEN
            exp_f := 1009;
        ELSIF x =- 1449 THEN
            exp_f := 1011;
        ELSIF x =- 1448 THEN
            exp_f := 1011;
        ELSIF x =- 1447 THEN
            exp_f := 1011;
        ELSIF x =- 1446 THEN
            exp_f := 1011;
        ELSIF x =- 1445 THEN
            exp_f := 1011;
        ELSIF x =- 1444 THEN
            exp_f := 1013;
        ELSIF x =- 1443 THEN
            exp_f := 1013;
        ELSIF x =- 1442 THEN
            exp_f := 1013;
        ELSIF x =- 1441 THEN
            exp_f := 1013;
        ELSIF x =- 1440 THEN
            exp_f := 1015;
        ELSIF x =- 1439 THEN
            exp_f := 1015;
        ELSIF x =- 1438 THEN
            exp_f := 1015;
        ELSIF x =- 1437 THEN
            exp_f := 1015;
        ELSIF x =- 1436 THEN
            exp_f := 1015;
        ELSIF x =- 1435 THEN
            exp_f := 1018;
        ELSIF x =- 1434 THEN
            exp_f := 1018;
        ELSIF x =- 1433 THEN
            exp_f := 1018;
        ELSIF x =- 1432 THEN
            exp_f := 1018;
        ELSIF x =- 1431 THEN
            exp_f := 1020;
        ELSIF x =- 1430 THEN
            exp_f := 1020;
        ELSIF x =- 1429 THEN
            exp_f := 1020;
        ELSIF x =- 1428 THEN
            exp_f := 1020;
        ELSIF x =- 1427 THEN
            exp_f := 1020;
        ELSIF x =- 1426 THEN
            exp_f := 1022;
        ELSIF x =- 1425 THEN
            exp_f := 1022;
        ELSIF x =- 1424 THEN
            exp_f := 1022;
        ELSIF x =- 1423 THEN
            exp_f := 1022;
        ELSIF x =- 1422 THEN
            exp_f := 1024;
        ELSIF x =- 1421 THEN
            exp_f := 1024;
        ELSIF x =- 1420 THEN
            exp_f := 1024;
        ELSIF x =- 1419 THEN
            exp_f := 1024;
        ELSIF x =- 1418 THEN
            exp_f := 1027;
        ELSIF x =- 1417 THEN
            exp_f := 1027;
        ELSIF x =- 1416 THEN
            exp_f := 1027;
        ELSIF x =- 1415 THEN
            exp_f := 1027;
        ELSIF x =- 1414 THEN
            exp_f := 1027;
        ELSIF x =- 1413 THEN
            exp_f := 1029;
        ELSIF x =- 1412 THEN
            exp_f := 1029;
        ELSIF x =- 1411 THEN
            exp_f := 1029;
        ELSIF x =- 1410 THEN
            exp_f := 1029;
        ELSIF x =- 1409 THEN
            exp_f := 1031;
        ELSIF x =- 1408 THEN
            exp_f := 1031;
        ELSIF x =- 1407 THEN
            exp_f := 1031;
        ELSIF x =- 1406 THEN
            exp_f := 1031;
        ELSIF x =- 1405 THEN
            exp_f := 1031;
        ELSIF x =- 1404 THEN
            exp_f := 1033;
        ELSIF x =- 1403 THEN
            exp_f := 1033;
        ELSIF x =- 1402 THEN
            exp_f := 1033;
        ELSIF x =- 1401 THEN
            exp_f := 1033;
        ELSIF x =- 1400 THEN
            exp_f := 1036;
        ELSIF x =- 1399 THEN
            exp_f := 1036;
        ELSIF x =- 1398 THEN
            exp_f := 1036;
        ELSIF x =- 1397 THEN
            exp_f := 1036;
        ELSIF x =- 1396 THEN
            exp_f := 1038;
        ELSIF x =- 1395 THEN
            exp_f := 1038;
        ELSIF x =- 1394 THEN
            exp_f := 1038;
        ELSIF x =- 1393 THEN
            exp_f := 1038;
        ELSIF x =- 1392 THEN
            exp_f := 1038;
        ELSIF x =- 1391 THEN
            exp_f := 1040;
        ELSIF x =- 1390 THEN
            exp_f := 1040;
        ELSIF x =- 1389 THEN
            exp_f := 1040;
        ELSIF x =- 1388 THEN
            exp_f := 1040;
        ELSIF x =- 1387 THEN
            exp_f := 1042;
        ELSIF x =- 1386 THEN
            exp_f := 1042;
        ELSIF x =- 1385 THEN
            exp_f := 1042;
        ELSIF x =- 1384 THEN
            exp_f := 1042;
        ELSIF x =- 1383 THEN
            exp_f := 1042;
        ELSIF x =- 1382 THEN
            exp_f := 1045;
        ELSIF x =- 1381 THEN
            exp_f := 1045;
        ELSIF x =- 1380 THEN
            exp_f := 1045;
        ELSIF x =- 1379 THEN
            exp_f := 1045;
        ELSIF x =- 1378 THEN
            exp_f := 1047;
        ELSIF x =- 1377 THEN
            exp_f := 1047;
        ELSIF x =- 1376 THEN
            exp_f := 1047;
        ELSIF x =- 1375 THEN
            exp_f := 1047;
        ELSIF x =- 1374 THEN
            exp_f := 1049;
        ELSIF x =- 1373 THEN
            exp_f := 1049;
        ELSIF x =- 1372 THEN
            exp_f := 1049;
        ELSIF x =- 1371 THEN
            exp_f := 1049;
        ELSIF x =- 1370 THEN
            exp_f := 1049;
        ELSIF x =- 1369 THEN
            exp_f := 1052;
        ELSIF x =- 1368 THEN
            exp_f := 1052;
        ELSIF x =- 1367 THEN
            exp_f := 1052;
        ELSIF x =- 1366 THEN
            exp_f := 1052;
        ELSIF x =- 1365 THEN
            exp_f := 1054;
        ELSIF x =- 1364 THEN
            exp_f := 1054;
        ELSIF x =- 1363 THEN
            exp_f := 1054;
        ELSIF x =- 1362 THEN
            exp_f := 1054;
        ELSIF x =- 1361 THEN
            exp_f := 1054;
        ELSIF x =- 1360 THEN
            exp_f := 1056;
        ELSIF x =- 1359 THEN
            exp_f := 1056;
        ELSIF x =- 1358 THEN
            exp_f := 1056;
        ELSIF x =- 1357 THEN
            exp_f := 1056;
        ELSIF x =- 1356 THEN
            exp_f := 1058;
        ELSIF x =- 1355 THEN
            exp_f := 1058;
        ELSIF x =- 1354 THEN
            exp_f := 1058;
        ELSIF x =- 1353 THEN
            exp_f := 1058;
        ELSIF x =- 1352 THEN
            exp_f := 1061;
        ELSIF x =- 1351 THEN
            exp_f := 1061;
        ELSIF x =- 1350 THEN
            exp_f := 1061;
        ELSIF x =- 1349 THEN
            exp_f := 1061;
        ELSIF x =- 1348 THEN
            exp_f := 1061;
        ELSIF x =- 1347 THEN
            exp_f := 1063;
        ELSIF x =- 1346 THEN
            exp_f := 1063;
        ELSIF x =- 1345 THEN
            exp_f := 1063;
        ELSIF x =- 1344 THEN
            exp_f := 1063;
        ELSIF x =- 1343 THEN
            exp_f := 1065;
        ELSIF x =- 1342 THEN
            exp_f := 1065;
        ELSIF x =- 1341 THEN
            exp_f := 1065;
        ELSIF x =- 1340 THEN
            exp_f := 1065;
        ELSIF x =- 1339 THEN
            exp_f := 1065;
        ELSIF x =- 1338 THEN
            exp_f := 1068;
        ELSIF x =- 1337 THEN
            exp_f := 1068;
        ELSIF x =- 1336 THEN
            exp_f := 1068;
        ELSIF x =- 1335 THEN
            exp_f := 1068;
        ELSIF x =- 1334 THEN
            exp_f := 1070;
        ELSIF x =- 1333 THEN
            exp_f := 1070;
        ELSIF x =- 1332 THEN
            exp_f := 1070;
        ELSIF x =- 1331 THEN
            exp_f := 1070;
        ELSIF x =- 1330 THEN
            exp_f := 1072;
        ELSIF x =- 1329 THEN
            exp_f := 1072;
        ELSIF x =- 1328 THEN
            exp_f := 1072;
        ELSIF x =- 1327 THEN
            exp_f := 1072;
        ELSIF x =- 1326 THEN
            exp_f := 1072;
        ELSIF x =- 1325 THEN
            exp_f := 1075;
        ELSIF x =- 1324 THEN
            exp_f := 1075;
        ELSIF x =- 1323 THEN
            exp_f := 1075;
        ELSIF x =- 1322 THEN
            exp_f := 1075;
        ELSIF x =- 1321 THEN
            exp_f := 1077;
        ELSIF x =- 1320 THEN
            exp_f := 1077;
        ELSIF x =- 1319 THEN
            exp_f := 1077;
        ELSIF x =- 1318 THEN
            exp_f := 1077;
        ELSIF x =- 1317 THEN
            exp_f := 1077;
        ELSIF x =- 1316 THEN
            exp_f := 1079;
        ELSIF x =- 1315 THEN
            exp_f := 1079;
        ELSIF x =- 1314 THEN
            exp_f := 1079;
        ELSIF x =- 1313 THEN
            exp_f := 1079;
        ELSIF x =- 1312 THEN
            exp_f := 1082;
        ELSIF x =- 1311 THEN
            exp_f := 1082;
        ELSIF x =- 1310 THEN
            exp_f := 1082;
        ELSIF x =- 1309 THEN
            exp_f := 1082;
        ELSIF x =- 1308 THEN
            exp_f := 1084;
        ELSIF x =- 1307 THEN
            exp_f := 1084;
        ELSIF x =- 1306 THEN
            exp_f := 1084;
        ELSIF x =- 1305 THEN
            exp_f := 1084;
        ELSIF x =- 1304 THEN
            exp_f := 1084;
        ELSIF x =- 1303 THEN
            exp_f := 1086;
        ELSIF x =- 1302 THEN
            exp_f := 1086;
        ELSIF x =- 1301 THEN
            exp_f := 1086;
        ELSIF x =- 1300 THEN
            exp_f := 1086;
        ELSIF x =- 1299 THEN
            exp_f := 1089;
        ELSIF x =- 1298 THEN
            exp_f := 1089;
        ELSIF x =- 1297 THEN
            exp_f := 1089;
        ELSIF x =- 1296 THEN
            exp_f := 1089;
        ELSIF x =- 1295 THEN
            exp_f := 1089;
        ELSIF x =- 1294 THEN
            exp_f := 1091;
        ELSIF x =- 1293 THEN
            exp_f := 1091;
        ELSIF x =- 1292 THEN
            exp_f := 1091;
        ELSIF x =- 1291 THEN
            exp_f := 1091;
        ELSIF x =- 1290 THEN
            exp_f := 1093;
        ELSIF x =- 1289 THEN
            exp_f := 1093;
        ELSIF x =- 1288 THEN
            exp_f := 1093;
        ELSIF x =- 1287 THEN
            exp_f := 1093;
        ELSIF x =- 1286 THEN
            exp_f := 1096;
        ELSIF x =- 1285 THEN
            exp_f := 1096;
        ELSIF x =- 1284 THEN
            exp_f := 1096;
        ELSIF x =- 1283 THEN
            exp_f := 1096;
        ELSIF x =- 1282 THEN
            exp_f := 1096;
        ELSIF x =- 1281 THEN
            exp_f := 1098;
        ELSIF x =- 1280 THEN
            exp_f := 1098;
        ELSIF x =- 1279 THEN
            exp_f := 1098;
        ELSIF x =- 1278 THEN
            exp_f := 1098;
        ELSIF x =- 1277 THEN
            exp_f := 1100;
        ELSIF x =- 1276 THEN
            exp_f := 1100;
        ELSIF x =- 1275 THEN
            exp_f := 1100;
        ELSIF x =- 1274 THEN
            exp_f := 1100;
        ELSIF x =- 1273 THEN
            exp_f := 1100;
        ELSIF x =- 1272 THEN
            exp_f := 1103;
        ELSIF x =- 1271 THEN
            exp_f := 1103;
        ELSIF x =- 1270 THEN
            exp_f := 1103;
        ELSIF x =- 1269 THEN
            exp_f := 1103;
        ELSIF x =- 1268 THEN
            exp_f := 1105;
        ELSIF x =- 1267 THEN
            exp_f := 1105;
        ELSIF x =- 1266 THEN
            exp_f := 1105;
        ELSIF x =- 1265 THEN
            exp_f := 1105;
        ELSIF x =- 1264 THEN
            exp_f := 1107;
        ELSIF x =- 1263 THEN
            exp_f := 1107;
        ELSIF x =- 1262 THEN
            exp_f := 1107;
        ELSIF x =- 1261 THEN
            exp_f := 1107;
        ELSIF x =- 1260 THEN
            exp_f := 1107;
        ELSIF x =- 1259 THEN
            exp_f := 1110;
        ELSIF x =- 1258 THEN
            exp_f := 1110;
        ELSIF x =- 1257 THEN
            exp_f := 1110;
        ELSIF x =- 1256 THEN
            exp_f := 1110;
        ELSIF x =- 1255 THEN
            exp_f := 1112;
        ELSIF x =- 1254 THEN
            exp_f := 1112;
        ELSIF x =- 1253 THEN
            exp_f := 1112;
        ELSIF x =- 1252 THEN
            exp_f := 1112;
        ELSIF x =- 1251 THEN
            exp_f := 1112;
        ELSIF x =- 1250 THEN
            exp_f := 1115;
        ELSIF x =- 1249 THEN
            exp_f := 1115;
        ELSIF x =- 1248 THEN
            exp_f := 1115;
        ELSIF x =- 1247 THEN
            exp_f := 1115;
        ELSIF x =- 1246 THEN
            exp_f := 1117;
        ELSIF x =- 1245 THEN
            exp_f := 1117;
        ELSIF x =- 1244 THEN
            exp_f := 1117;
        ELSIF x =- 1243 THEN
            exp_f := 1117;
        ELSIF x =- 1242 THEN
            exp_f := 1119;
        ELSIF x =- 1241 THEN
            exp_f := 1119;
        ELSIF x =- 1240 THEN
            exp_f := 1119;
        ELSIF x =- 1239 THEN
            exp_f := 1119;
        ELSIF x =- 1238 THEN
            exp_f := 1119;
        ELSIF x =- 1237 THEN
            exp_f := 1122;
        ELSIF x =- 1236 THEN
            exp_f := 1122;
        ELSIF x =- 1235 THEN
            exp_f := 1122;
        ELSIF x =- 1234 THEN
            exp_f := 1122;
        ELSIF x =- 1233 THEN
            exp_f := 1124;
        ELSIF x =- 1232 THEN
            exp_f := 1124;
        ELSIF x =- 1231 THEN
            exp_f := 1124;
        ELSIF x =- 1230 THEN
            exp_f := 1124;
        ELSIF x =- 1229 THEN
            exp_f := 1124;
        ELSIF x =- 1228 THEN
            exp_f := 1127;
        ELSIF x =- 1227 THEN
            exp_f := 1127;
        ELSIF x =- 1226 THEN
            exp_f := 1127;
        ELSIF x =- 1225 THEN
            exp_f := 1127;
        ELSIF x =- 1224 THEN
            exp_f := 1129;
        ELSIF x =- 1223 THEN
            exp_f := 1129;
        ELSIF x =- 1222 THEN
            exp_f := 1129;
        ELSIF x =- 1221 THEN
            exp_f := 1129;
        ELSIF x =- 1220 THEN
            exp_f := 1129;
        ELSIF x =- 1219 THEN
            exp_f := 1131;
        ELSIF x =- 1218 THEN
            exp_f := 1131;
        ELSIF x =- 1217 THEN
            exp_f := 1131;
        ELSIF x =- 1216 THEN
            exp_f := 1131;
        ELSIF x =- 1215 THEN
            exp_f := 1134;
        ELSIF x =- 1214 THEN
            exp_f := 1134;
        ELSIF x =- 1213 THEN
            exp_f := 1134;
        ELSIF x =- 1212 THEN
            exp_f := 1134;
        ELSIF x =- 1211 THEN
            exp_f := 1136;
        ELSIF x =- 1210 THEN
            exp_f := 1136;
        ELSIF x =- 1209 THEN
            exp_f := 1136;
        ELSIF x =- 1208 THEN
            exp_f := 1136;
        ELSIF x =- 1207 THEN
            exp_f := 1136;
        ELSIF x =- 1206 THEN
            exp_f := 1139;
        ELSIF x =- 1205 THEN
            exp_f := 1139;
        ELSIF x =- 1204 THEN
            exp_f := 1139;
        ELSIF x =- 1203 THEN
            exp_f := 1139;
        ELSIF x =- 1202 THEN
            exp_f := 1141;
        ELSIF x =- 1201 THEN
            exp_f := 1141;
        ELSIF x =- 1200 THEN
            exp_f := 1141;
        ELSIF x =- 1199 THEN
            exp_f := 1141;
        ELSIF x =- 1198 THEN
            exp_f := 1141;
        ELSIF x =- 1197 THEN
            exp_f := 1144;
        ELSIF x =- 1196 THEN
            exp_f := 1144;
        ELSIF x =- 1195 THEN
            exp_f := 1144;
        ELSIF x =- 1194 THEN
            exp_f := 1144;
        ELSIF x =- 1193 THEN
            exp_f := 1146;
        ELSIF x =- 1192 THEN
            exp_f := 1146;
        ELSIF x =- 1191 THEN
            exp_f := 1146;
        ELSIF x =- 1190 THEN
            exp_f := 1146;
        ELSIF x =- 1189 THEN
            exp_f := 1148;
        ELSIF x =- 1188 THEN
            exp_f := 1148;
        ELSIF x =- 1187 THEN
            exp_f := 1148;
        ELSIF x =- 1186 THEN
            exp_f := 1148;
        ELSIF x =- 1185 THEN
            exp_f := 1148;
        ELSIF x =- 1184 THEN
            exp_f := 1151;
        ELSIF x =- 1183 THEN
            exp_f := 1151;
        ELSIF x =- 1182 THEN
            exp_f := 1151;
        ELSIF x =- 1181 THEN
            exp_f := 1151;
        ELSIF x =- 1180 THEN
            exp_f := 1153;
        ELSIF x =- 1179 THEN
            exp_f := 1153;
        ELSIF x =- 1178 THEN
            exp_f := 1153;
        ELSIF x =- 1177 THEN
            exp_f := 1153;
        ELSIF x =- 1176 THEN
            exp_f := 1153;
        ELSIF x =- 1175 THEN
            exp_f := 1156;
        ELSIF x =- 1174 THEN
            exp_f := 1156;
        ELSIF x =- 1173 THEN
            exp_f := 1156;
        ELSIF x =- 1172 THEN
            exp_f := 1156;
        ELSIF x =- 1171 THEN
            exp_f := 1158;
        ELSIF x =- 1170 THEN
            exp_f := 1158;
        ELSIF x =- 1169 THEN
            exp_f := 1158;
        ELSIF x =- 1168 THEN
            exp_f := 1158;
        ELSIF x =- 1167 THEN
            exp_f := 1161;
        ELSIF x =- 1166 THEN
            exp_f := 1161;
        ELSIF x =- 1165 THEN
            exp_f := 1161;
        ELSIF x =- 1164 THEN
            exp_f := 1161;
        ELSIF x =- 1163 THEN
            exp_f := 1161;
        ELSIF x =- 1162 THEN
            exp_f := 1163;
        ELSIF x =- 1161 THEN
            exp_f := 1163;
        ELSIF x =- 1160 THEN
            exp_f := 1163;
        ELSIF x =- 1159 THEN
            exp_f := 1163;
        ELSIF x =- 1158 THEN
            exp_f := 1166;
        ELSIF x =- 1157 THEN
            exp_f := 1166;
        ELSIF x =- 1156 THEN
            exp_f := 1166;
        ELSIF x =- 1155 THEN
            exp_f := 1166;
        ELSIF x =- 1154 THEN
            exp_f := 1166;
        ELSIF x =- 1153 THEN
            exp_f := 1168;
        ELSIF x =- 1152 THEN
            exp_f := 1168;
        ELSIF x =- 1151 THEN
            exp_f := 1168;
        ELSIF x =- 1150 THEN
            exp_f := 1168;
        ELSIF x =- 1149 THEN
            exp_f := 1170;
        ELSIF x =- 1148 THEN
            exp_f := 1170;
        ELSIF x =- 1147 THEN
            exp_f := 1170;
        ELSIF x =- 1146 THEN
            exp_f := 1170;
        ELSIF x =- 1145 THEN
            exp_f := 1173;
        ELSIF x =- 1144 THEN
            exp_f := 1173;
        ELSIF x =- 1143 THEN
            exp_f := 1173;
        ELSIF x =- 1142 THEN
            exp_f := 1173;
        ELSIF x =- 1141 THEN
            exp_f := 1173;
        ELSIF x =- 1140 THEN
            exp_f := 1175;
        ELSIF x =- 1139 THEN
            exp_f := 1175;
        ELSIF x =- 1138 THEN
            exp_f := 1175;
        ELSIF x =- 1137 THEN
            exp_f := 1175;
        ELSIF x =- 1136 THEN
            exp_f := 1178;
        ELSIF x =- 1135 THEN
            exp_f := 1178;
        ELSIF x =- 1134 THEN
            exp_f := 1178;
        ELSIF x =- 1133 THEN
            exp_f := 1178;
        ELSIF x =- 1132 THEN
            exp_f := 1178;
        ELSIF x =- 1131 THEN
            exp_f := 1180;
        ELSIF x =- 1130 THEN
            exp_f := 1180;
        ELSIF x =- 1129 THEN
            exp_f := 1180;
        ELSIF x =- 1128 THEN
            exp_f := 1180;
        ELSIF x =- 1127 THEN
            exp_f := 1183;
        ELSIF x =- 1126 THEN
            exp_f := 1183;
        ELSIF x =- 1125 THEN
            exp_f := 1183;
        ELSIF x =- 1124 THEN
            exp_f := 1183;
        ELSIF x =- 1123 THEN
            exp_f := 1185;
        ELSIF x =- 1122 THEN
            exp_f := 1185;
        ELSIF x =- 1121 THEN
            exp_f := 1185;
        ELSIF x =- 1120 THEN
            exp_f := 1185;
        ELSIF x =- 1119 THEN
            exp_f := 1185;
        ELSIF x =- 1118 THEN
            exp_f := 1188;
        ELSIF x =- 1117 THEN
            exp_f := 1188;
        ELSIF x =- 1116 THEN
            exp_f := 1188;
        ELSIF x =- 1115 THEN
            exp_f := 1188;
        ELSIF x =- 1114 THEN
            exp_f := 1190;
        ELSIF x =- 1113 THEN
            exp_f := 1190;
        ELSIF x =- 1112 THEN
            exp_f := 1190;
        ELSIF x =- 1111 THEN
            exp_f := 1190;
        ELSIF x =- 1110 THEN
            exp_f := 1190;
        ELSIF x =- 1109 THEN
            exp_f := 1193;
        ELSIF x =- 1108 THEN
            exp_f := 1193;
        ELSIF x =- 1107 THEN
            exp_f := 1193;
        ELSIF x =- 1106 THEN
            exp_f := 1193;
        ELSIF x =- 1105 THEN
            exp_f := 1195;
        ELSIF x =- 1104 THEN
            exp_f := 1195;
        ELSIF x =- 1103 THEN
            exp_f := 1195;
        ELSIF x =- 1102 THEN
            exp_f := 1195;
        ELSIF x =- 1101 THEN
            exp_f := 1198;
        ELSIF x =- 1100 THEN
            exp_f := 1198;
        ELSIF x =- 1099 THEN
            exp_f := 1198;
        ELSIF x =- 1098 THEN
            exp_f := 1198;
        ELSIF x =- 1097 THEN
            exp_f := 1198;
        ELSIF x =- 1096 THEN
            exp_f := 1200;
        ELSIF x =- 1095 THEN
            exp_f := 1200;
        ELSIF x =- 1094 THEN
            exp_f := 1200;
        ELSIF x =- 1093 THEN
            exp_f := 1200;
        ELSIF x =- 1092 THEN
            exp_f := 1203;
        ELSIF x =- 1091 THEN
            exp_f := 1203;
        ELSIF x =- 1090 THEN
            exp_f := 1203;
        ELSIF x =- 1089 THEN
            exp_f := 1203;
        ELSIF x =- 1088 THEN
            exp_f := 1203;
        ELSIF x =- 1087 THEN
            exp_f := 1205;
        ELSIF x =- 1086 THEN
            exp_f := 1205;
        ELSIF x =- 1085 THEN
            exp_f := 1205;
        ELSIF x =- 1084 THEN
            exp_f := 1205;
        ELSIF x =- 1083 THEN
            exp_f := 1208;
        ELSIF x =- 1082 THEN
            exp_f := 1208;
        ELSIF x =- 1081 THEN
            exp_f := 1208;
        ELSIF x =- 1080 THEN
            exp_f := 1208;
        ELSIF x =- 1079 THEN
            exp_f := 1210;
        ELSIF x =- 1078 THEN
            exp_f := 1210;
        ELSIF x =- 1077 THEN
            exp_f := 1210;
        ELSIF x =- 1076 THEN
            exp_f := 1210;
        ELSIF x =- 1075 THEN
            exp_f := 1210;
        ELSIF x =- 1074 THEN
            exp_f := 1213;
        ELSIF x =- 1073 THEN
            exp_f := 1213;
        ELSIF x =- 1072 THEN
            exp_f := 1213;
        ELSIF x =- 1071 THEN
            exp_f := 1213;
        ELSIF x =- 1070 THEN
            exp_f := 1216;
        ELSIF x =- 1069 THEN
            exp_f := 1216;
        ELSIF x =- 1068 THEN
            exp_f := 1216;
        ELSIF x =- 1067 THEN
            exp_f := 1216;
        ELSIF x =- 1066 THEN
            exp_f := 1216;
        ELSIF x =- 1065 THEN
            exp_f := 1218;
        ELSIF x =- 1064 THEN
            exp_f := 1218;
        ELSIF x =- 1063 THEN
            exp_f := 1218;
        ELSIF x =- 1062 THEN
            exp_f := 1218;
        ELSIF x =- 1061 THEN
            exp_f := 1221;
        ELSIF x =- 1060 THEN
            exp_f := 1221;
        ELSIF x =- 1059 THEN
            exp_f := 1221;
        ELSIF x =- 1058 THEN
            exp_f := 1221;
        ELSIF x =- 1057 THEN
            exp_f := 1223;
        ELSIF x =- 1056 THEN
            exp_f := 1223;
        ELSIF x =- 1055 THEN
            exp_f := 1223;
        ELSIF x =- 1054 THEN
            exp_f := 1223;
        ELSIF x =- 1053 THEN
            exp_f := 1223;
        ELSIF x =- 1052 THEN
            exp_f := 1226;
        ELSIF x =- 1051 THEN
            exp_f := 1226;
        ELSIF x =- 1050 THEN
            exp_f := 1226;
        ELSIF x =- 1049 THEN
            exp_f := 1226;
        ELSIF x =- 1048 THEN
            exp_f := 1228;
        ELSIF x =- 1047 THEN
            exp_f := 1228;
        ELSIF x =- 1046 THEN
            exp_f := 1228;
        ELSIF x =- 1045 THEN
            exp_f := 1228;
        ELSIF x =- 1044 THEN
            exp_f := 1228;
        ELSIF x =- 1043 THEN
            exp_f := 1231;
        ELSIF x =- 1042 THEN
            exp_f := 1231;
        ELSIF x =- 1041 THEN
            exp_f := 1231;
        ELSIF x =- 1040 THEN
            exp_f := 1231;
        ELSIF x =- 1039 THEN
            exp_f := 1233;
        ELSIF x =- 1038 THEN
            exp_f := 1233;
        ELSIF x =- 1037 THEN
            exp_f := 1233;
        ELSIF x =- 1036 THEN
            exp_f := 1233;
        ELSIF x =- 1035 THEN
            exp_f := 1236;
        ELSIF x =- 1034 THEN
            exp_f := 1236;
        ELSIF x =- 1033 THEN
            exp_f := 1236;
        ELSIF x =- 1032 THEN
            exp_f := 1236;
        ELSIF x =- 1031 THEN
            exp_f := 1236;
        ELSIF x =- 1030 THEN
            exp_f := 1239;
        ELSIF x =- 1029 THEN
            exp_f := 1239;
        ELSIF x =- 1028 THEN
            exp_f := 1239;
        ELSIF x =- 1027 THEN
            exp_f := 1239;
        ELSIF x =- 1026 THEN
            exp_f := 1241;
        ELSIF x =- 1025 THEN
            exp_f := 1241;
        ELSIF x =- 1024 THEN
            exp_f := 1241;
        ELSIF x =- 1023 THEN
            exp_f := 1241;
        ELSIF x =- 1022 THEN
            exp_f := 1241;
        ELSIF x =- 1021 THEN
            exp_f := 1244;
        ELSIF x =- 1020 THEN
            exp_f := 1244;
        ELSIF x =- 1019 THEN
            exp_f := 1244;
        ELSIF x =- 1018 THEN
            exp_f := 1244;
        ELSIF x =- 1017 THEN
            exp_f := 1246;
        ELSIF x =- 1016 THEN
            exp_f := 1246;
        ELSIF x =- 1015 THEN
            exp_f := 1246;
        ELSIF x =- 1014 THEN
            exp_f := 1246;
        ELSIF x =- 1013 THEN
            exp_f := 1249;
        ELSIF x =- 1012 THEN
            exp_f := 1249;
        ELSIF x =- 1011 THEN
            exp_f := 1249;
        ELSIF x =- 1010 THEN
            exp_f := 1249;
        ELSIF x =- 1009 THEN
            exp_f := 1252;
        ELSIF x =- 1008 THEN
            exp_f := 1252;
        ELSIF x =- 1007 THEN
            exp_f := 1252;
        ELSIF x =- 1006 THEN
            exp_f := 1252;
        ELSIF x =- 1005 THEN
            exp_f := 1254;
        ELSIF x =- 1004 THEN
            exp_f := 1254;
        ELSIF x =- 1003 THEN
            exp_f := 1254;
        ELSIF x =- 1002 THEN
            exp_f := 1254;
        ELSIF x =- 1001 THEN
            exp_f := 1257;
        ELSIF x =- 1000 THEN
            exp_f := 1257;
        ELSIF x =- 999 THEN
            exp_f := 1257;
        ELSIF x =- 998 THEN
            exp_f := 1257;
        ELSIF x =- 997 THEN
            exp_f := 1259;
        ELSIF x =- 996 THEN
            exp_f := 1259;
        ELSIF x =- 995 THEN
            exp_f := 1259;
        ELSIF x =- 994 THEN
            exp_f := 1259;
        ELSIF x =- 993 THEN
            exp_f := 1259;
        ELSIF x =- 992 THEN
            exp_f := 1262;
        ELSIF x =- 991 THEN
            exp_f := 1262;
        ELSIF x =- 990 THEN
            exp_f := 1262;
        ELSIF x =- 989 THEN
            exp_f := 1262;
        ELSIF x =- 988 THEN
            exp_f := 1265;
        ELSIF x =- 987 THEN
            exp_f := 1265;
        ELSIF x =- 986 THEN
            exp_f := 1265;
        ELSIF x =- 985 THEN
            exp_f := 1265;
        ELSIF x =- 984 THEN
            exp_f := 1267;
        ELSIF x =- 983 THEN
            exp_f := 1267;
        ELSIF x =- 982 THEN
            exp_f := 1267;
        ELSIF x =- 981 THEN
            exp_f := 1267;
        ELSIF x =- 980 THEN
            exp_f := 1270;
        ELSIF x =- 979 THEN
            exp_f := 1270;
        ELSIF x =- 978 THEN
            exp_f := 1270;
        ELSIF x =- 977 THEN
            exp_f := 1270;
        ELSIF x =- 976 THEN
            exp_f := 1272;
        ELSIF x =- 975 THEN
            exp_f := 1272;
        ELSIF x =- 974 THEN
            exp_f := 1272;
        ELSIF x =- 973 THEN
            exp_f := 1272;
        ELSIF x =- 972 THEN
            exp_f := 1275;
        ELSIF x =- 971 THEN
            exp_f := 1275;
        ELSIF x =- 970 THEN
            exp_f := 1275;
        ELSIF x =- 969 THEN
            exp_f := 1275;
        ELSIF x =- 968 THEN
            exp_f := 1278;
        ELSIF x =- 967 THEN
            exp_f := 1278;
        ELSIF x =- 966 THEN
            exp_f := 1278;
        ELSIF x =- 965 THEN
            exp_f := 1278;
        ELSIF x =- 964 THEN
            exp_f := 1280;
        ELSIF x =- 963 THEN
            exp_f := 1280;
        ELSIF x =- 962 THEN
            exp_f := 1280;
        ELSIF x =- 961 THEN
            exp_f := 1280;
        ELSIF x =- 960 THEN
            exp_f := 1280;
        ELSIF x =- 959 THEN
            exp_f := 1283;
        ELSIF x =- 958 THEN
            exp_f := 1283;
        ELSIF x =- 957 THEN
            exp_f := 1283;
        ELSIF x =- 956 THEN
            exp_f := 1283;
        ELSIF x =- 955 THEN
            exp_f := 1286;
        ELSIF x =- 954 THEN
            exp_f := 1286;
        ELSIF x =- 953 THEN
            exp_f := 1286;
        ELSIF x =- 952 THEN
            exp_f := 1286;
        ELSIF x =- 951 THEN
            exp_f := 1288;
        ELSIF x =- 950 THEN
            exp_f := 1288;
        ELSIF x =- 949 THEN
            exp_f := 1288;
        ELSIF x =- 948 THEN
            exp_f := 1288;
        ELSIF x =- 947 THEN
            exp_f := 1291;
        ELSIF x =- 946 THEN
            exp_f := 1291;
        ELSIF x =- 945 THEN
            exp_f := 1291;
        ELSIF x =- 944 THEN
            exp_f := 1291;
        ELSIF x =- 943 THEN
            exp_f := 1294;
        ELSIF x =- 942 THEN
            exp_f := 1294;
        ELSIF x =- 941 THEN
            exp_f := 1294;
        ELSIF x =- 940 THEN
            exp_f := 1294;
        ELSIF x =- 939 THEN
            exp_f := 1296;
        ELSIF x =- 938 THEN
            exp_f := 1296;
        ELSIF x =- 937 THEN
            exp_f := 1296;
        ELSIF x =- 936 THEN
            exp_f := 1296;
        ELSIF x =- 935 THEN
            exp_f := 1299;
        ELSIF x =- 934 THEN
            exp_f := 1299;
        ELSIF x =- 933 THEN
            exp_f := 1299;
        ELSIF x =- 932 THEN
            exp_f := 1299;
        ELSIF x =- 931 THEN
            exp_f := 1299;
        ELSIF x =- 930 THEN
            exp_f := 1302;
        ELSIF x =- 929 THEN
            exp_f := 1302;
        ELSIF x =- 928 THEN
            exp_f := 1302;
        ELSIF x =- 927 THEN
            exp_f := 1302;
        ELSIF x =- 926 THEN
            exp_f := 1304;
        ELSIF x =- 925 THEN
            exp_f := 1304;
        ELSIF x =- 924 THEN
            exp_f := 1304;
        ELSIF x =- 923 THEN
            exp_f := 1304;
        ELSIF x =- 922 THEN
            exp_f := 1307;
        ELSIF x =- 921 THEN
            exp_f := 1307;
        ELSIF x =- 920 THEN
            exp_f := 1307;
        ELSIF x =- 919 THEN
            exp_f := 1307;
        ELSIF x =- 918 THEN
            exp_f := 1310;
        ELSIF x =- 917 THEN
            exp_f := 1310;
        ELSIF x =- 916 THEN
            exp_f := 1310;
        ELSIF x =- 915 THEN
            exp_f := 1310;
        ELSIF x =- 914 THEN
            exp_f := 1312;
        ELSIF x =- 913 THEN
            exp_f := 1312;
        ELSIF x =- 912 THEN
            exp_f := 1312;
        ELSIF x =- 911 THEN
            exp_f := 1312;
        ELSIF x =- 910 THEN
            exp_f := 1315;
        ELSIF x =- 909 THEN
            exp_f := 1315;
        ELSIF x =- 908 THEN
            exp_f := 1315;
        ELSIF x =- 907 THEN
            exp_f := 1315;
        ELSIF x =- 906 THEN
            exp_f := 1318;
        ELSIF x =- 905 THEN
            exp_f := 1318;
        ELSIF x =- 904 THEN
            exp_f := 1318;
        ELSIF x =- 903 THEN
            exp_f := 1318;
        ELSIF x =- 902 THEN
            exp_f := 1318;
        ELSIF x =- 901 THEN
            exp_f := 1320;
        ELSIF x =- 900 THEN
            exp_f := 1320;
        ELSIF x =- 899 THEN
            exp_f := 1320;
        ELSIF x =- 898 THEN
            exp_f := 1320;
        ELSIF x =- 897 THEN
            exp_f := 1323;
        ELSIF x =- 896 THEN
            exp_f := 1323;
        ELSIF x =- 895 THEN
            exp_f := 1323;
        ELSIF x =- 894 THEN
            exp_f := 1323;
        ELSIF x =- 893 THEN
            exp_f := 1326;
        ELSIF x =- 892 THEN
            exp_f := 1326;
        ELSIF x =- 891 THEN
            exp_f := 1326;
        ELSIF x =- 890 THEN
            exp_f := 1326;
        ELSIF x =- 889 THEN
            exp_f := 1329;
        ELSIF x =- 888 THEN
            exp_f := 1329;
        ELSIF x =- 887 THEN
            exp_f := 1329;
        ELSIF x =- 886 THEN
            exp_f := 1329;
        ELSIF x =- 885 THEN
            exp_f := 1331;
        ELSIF x =- 884 THEN
            exp_f := 1331;
        ELSIF x =- 883 THEN
            exp_f := 1331;
        ELSIF x =- 882 THEN
            exp_f := 1331;
        ELSIF x =- 881 THEN
            exp_f := 1334;
        ELSIF x =- 880 THEN
            exp_f := 1334;
        ELSIF x =- 879 THEN
            exp_f := 1334;
        ELSIF x =- 878 THEN
            exp_f := 1334;
        ELSIF x =- 877 THEN
            exp_f := 1337;
        ELSIF x =- 876 THEN
            exp_f := 1337;
        ELSIF x =- 875 THEN
            exp_f := 1337;
        ELSIF x =- 874 THEN
            exp_f := 1337;
        ELSIF x =- 873 THEN
            exp_f := 1337;
        ELSIF x =- 872 THEN
            exp_f := 1339;
        ELSIF x =- 871 THEN
            exp_f := 1339;
        ELSIF x =- 870 THEN
            exp_f := 1339;
        ELSIF x =- 869 THEN
            exp_f := 1339;
        ELSIF x =- 868 THEN
            exp_f := 1342;
        ELSIF x =- 867 THEN
            exp_f := 1342;
        ELSIF x =- 866 THEN
            exp_f := 1342;
        ELSIF x =- 865 THEN
            exp_f := 1342;
        ELSIF x =- 864 THEN
            exp_f := 1345;
        ELSIF x =- 863 THEN
            exp_f := 1345;
        ELSIF x =- 862 THEN
            exp_f := 1345;
        ELSIF x =- 861 THEN
            exp_f := 1345;
        ELSIF x =- 860 THEN
            exp_f := 1348;
        ELSIF x =- 859 THEN
            exp_f := 1348;
        ELSIF x =- 858 THEN
            exp_f := 1348;
        ELSIF x =- 857 THEN
            exp_f := 1348;
        ELSIF x =- 856 THEN
            exp_f := 1350;
        ELSIF x =- 855 THEN
            exp_f := 1350;
        ELSIF x =- 854 THEN
            exp_f := 1350;
        ELSIF x =- 853 THEN
            exp_f := 1350;
        ELSIF x =- 852 THEN
            exp_f := 1353;
        ELSIF x =- 851 THEN
            exp_f := 1353;
        ELSIF x =- 850 THEN
            exp_f := 1353;
        ELSIF x =- 849 THEN
            exp_f := 1353;
        ELSIF x =- 848 THEN
            exp_f := 1356;
        ELSIF x =- 847 THEN
            exp_f := 1356;
        ELSIF x =- 846 THEN
            exp_f := 1356;
        ELSIF x =- 845 THEN
            exp_f := 1356;
        ELSIF x =- 844 THEN
            exp_f := 1359;
        ELSIF x =- 843 THEN
            exp_f := 1359;
        ELSIF x =- 842 THEN
            exp_f := 1359;
        ELSIF x =- 841 THEN
            exp_f := 1359;
        ELSIF x =- 840 THEN
            exp_f := 1359;
        ELSIF x =- 839 THEN
            exp_f := 1362;
        ELSIF x =- 838 THEN
            exp_f := 1362;
        ELSIF x =- 837 THEN
            exp_f := 1362;
        ELSIF x =- 836 THEN
            exp_f := 1362;
        ELSIF x =- 835 THEN
            exp_f := 1364;
        ELSIF x =- 834 THEN
            exp_f := 1364;
        ELSIF x =- 833 THEN
            exp_f := 1364;
        ELSIF x =- 832 THEN
            exp_f := 1364;
        ELSIF x =- 831 THEN
            exp_f := 1367;
        ELSIF x =- 830 THEN
            exp_f := 1367;
        ELSIF x =- 829 THEN
            exp_f := 1367;
        ELSIF x =- 828 THEN
            exp_f := 1367;
        ELSIF x =- 827 THEN
            exp_f := 1370;
        ELSIF x =- 826 THEN
            exp_f := 1370;
        ELSIF x =- 825 THEN
            exp_f := 1370;
        ELSIF x =- 824 THEN
            exp_f := 1370;
        ELSIF x =- 823 THEN
            exp_f := 1373;
        ELSIF x =- 822 THEN
            exp_f := 1373;
        ELSIF x =- 821 THEN
            exp_f := 1373;
        ELSIF x =- 820 THEN
            exp_f := 1373;
        ELSIF x =- 819 THEN
            exp_f := 1375;
        ELSIF x =- 818 THEN
            exp_f := 1375;
        ELSIF x =- 817 THEN
            exp_f := 1375;
        ELSIF x =- 816 THEN
            exp_f := 1375;
        ELSIF x =- 815 THEN
            exp_f := 1378;
        ELSIF x =- 814 THEN
            exp_f := 1378;
        ELSIF x =- 813 THEN
            exp_f := 1378;
        ELSIF x =- 812 THEN
            exp_f := 1378;
        ELSIF x =- 811 THEN
            exp_f := 1378;
        ELSIF x =- 810 THEN
            exp_f := 1381;
        ELSIF x =- 809 THEN
            exp_f := 1381;
        ELSIF x =- 808 THEN
            exp_f := 1381;
        ELSIF x =- 807 THEN
            exp_f := 1381;
        ELSIF x =- 806 THEN
            exp_f := 1384;
        ELSIF x =- 805 THEN
            exp_f := 1384;
        ELSIF x =- 804 THEN
            exp_f := 1384;
        ELSIF x =- 803 THEN
            exp_f := 1384;
        ELSIF x =- 802 THEN
            exp_f := 1387;
        ELSIF x =- 801 THEN
            exp_f := 1387;
        ELSIF x =- 800 THEN
            exp_f := 1387;
        ELSIF x =- 799 THEN
            exp_f := 1387;
        ELSIF x =- 798 THEN
            exp_f := 1389;
        ELSIF x =- 797 THEN
            exp_f := 1389;
        ELSIF x =- 796 THEN
            exp_f := 1389;
        ELSIF x =- 795 THEN
            exp_f := 1389;
        ELSIF x =- 794 THEN
            exp_f := 1392;
        ELSIF x =- 793 THEN
            exp_f := 1392;
        ELSIF x =- 792 THEN
            exp_f := 1392;
        ELSIF x =- 791 THEN
            exp_f := 1392;
        ELSIF x =- 790 THEN
            exp_f := 1395;
        ELSIF x =- 789 THEN
            exp_f := 1395;
        ELSIF x =- 788 THEN
            exp_f := 1395;
        ELSIF x =- 787 THEN
            exp_f := 1395;
        ELSIF x =- 786 THEN
            exp_f := 1398;
        ELSIF x =- 785 THEN
            exp_f := 1398;
        ELSIF x =- 784 THEN
            exp_f := 1398;
        ELSIF x =- 783 THEN
            exp_f := 1398;
        ELSIF x =- 782 THEN
            exp_f := 1398;
        ELSIF x =- 781 THEN
            exp_f := 1401;
        ELSIF x =- 780 THEN
            exp_f := 1401;
        ELSIF x =- 779 THEN
            exp_f := 1401;
        ELSIF x =- 778 THEN
            exp_f := 1401;
        ELSIF x =- 777 THEN
            exp_f := 1404;
        ELSIF x =- 776 THEN
            exp_f := 1404;
        ELSIF x =- 775 THEN
            exp_f := 1404;
        ELSIF x =- 774 THEN
            exp_f := 1404;
        ELSIF x =- 773 THEN
            exp_f := 1406;
        ELSIF x =- 772 THEN
            exp_f := 1406;
        ELSIF x =- 771 THEN
            exp_f := 1406;
        ELSIF x =- 770 THEN
            exp_f := 1406;
        ELSIF x =- 769 THEN
            exp_f := 1409;
        ELSIF x =- 768 THEN
            exp_f := 1409;
        ELSIF x =- 767 THEN
            exp_f := 1409;
        ELSIF x =- 766 THEN
            exp_f := 1409;
        ELSIF x =- 765 THEN
            exp_f := 1412;
        ELSIF x =- 764 THEN
            exp_f := 1412;
        ELSIF x =- 763 THEN
            exp_f := 1412;
        ELSIF x =- 762 THEN
            exp_f := 1412;
        ELSIF x =- 761 THEN
            exp_f := 1415;
        ELSIF x =- 760 THEN
            exp_f := 1415;
        ELSIF x =- 759 THEN
            exp_f := 1415;
        ELSIF x =- 758 THEN
            exp_f := 1415;
        ELSIF x =- 757 THEN
            exp_f := 1418;
        ELSIF x =- 756 THEN
            exp_f := 1418;
        ELSIF x =- 755 THEN
            exp_f := 1418;
        ELSIF x =- 754 THEN
            exp_f := 1418;
        ELSIF x =- 753 THEN
            exp_f := 1421;
        ELSIF x =- 752 THEN
            exp_f := 1421;
        ELSIF x =- 751 THEN
            exp_f := 1421;
        ELSIF x =- 750 THEN
            exp_f := 1421;
        ELSIF x =- 749 THEN
            exp_f := 1421;
        ELSIF x =- 748 THEN
            exp_f := 1424;
        ELSIF x =- 747 THEN
            exp_f := 1424;
        ELSIF x =- 746 THEN
            exp_f := 1424;
        ELSIF x =- 745 THEN
            exp_f := 1424;
        ELSIF x =- 744 THEN
            exp_f := 1426;
        ELSIF x =- 743 THEN
            exp_f := 1426;
        ELSIF x =- 742 THEN
            exp_f := 1426;
        ELSIF x =- 741 THEN
            exp_f := 1426;
        ELSIF x =- 740 THEN
            exp_f := 1429;
        ELSIF x =- 739 THEN
            exp_f := 1429;
        ELSIF x =- 738 THEN
            exp_f := 1429;
        ELSIF x =- 737 THEN
            exp_f := 1429;
        ELSIF x =- 736 THEN
            exp_f := 1432;
        ELSIF x =- 735 THEN
            exp_f := 1432;
        ELSIF x =- 734 THEN
            exp_f := 1432;
        ELSIF x =- 733 THEN
            exp_f := 1432;
        ELSIF x =- 732 THEN
            exp_f := 1435;
        ELSIF x =- 731 THEN
            exp_f := 1435;
        ELSIF x =- 730 THEN
            exp_f := 1435;
        ELSIF x =- 729 THEN
            exp_f := 1435;
        ELSIF x =- 728 THEN
            exp_f := 1438;
        ELSIF x =- 727 THEN
            exp_f := 1438;
        ELSIF x =- 726 THEN
            exp_f := 1438;
        ELSIF x =- 725 THEN
            exp_f := 1438;
        ELSIF x =- 724 THEN
            exp_f := 1441;
        ELSIF x =- 723 THEN
            exp_f := 1441;
        ELSIF x =- 722 THEN
            exp_f := 1441;
        ELSIF x =- 721 THEN
            exp_f := 1441;
        ELSIF x =- 720 THEN
            exp_f := 1441;
        ELSIF x =- 719 THEN
            exp_f := 1444;
        ELSIF x =- 718 THEN
            exp_f := 1444;
        ELSIF x =- 717 THEN
            exp_f := 1444;
        ELSIF x =- 716 THEN
            exp_f := 1444;
        ELSIF x =- 715 THEN
            exp_f := 1447;
        ELSIF x =- 714 THEN
            exp_f := 1447;
        ELSIF x =- 713 THEN
            exp_f := 1447;
        ELSIF x =- 712 THEN
            exp_f := 1447;
        ELSIF x =- 711 THEN
            exp_f := 1450;
        ELSIF x =- 710 THEN
            exp_f := 1450;
        ELSIF x =- 709 THEN
            exp_f := 1450;
        ELSIF x =- 708 THEN
            exp_f := 1450;
        ELSIF x =- 707 THEN
            exp_f := 1453;
        ELSIF x =- 706 THEN
            exp_f := 1453;
        ELSIF x =- 705 THEN
            exp_f := 1453;
        ELSIF x =- 704 THEN
            exp_f := 1453;
        ELSIF x =- 703 THEN
            exp_f := 1456;
        ELSIF x =- 702 THEN
            exp_f := 1456;
        ELSIF x =- 701 THEN
            exp_f := 1456;
        ELSIF x =- 700 THEN
            exp_f := 1456;
        ELSIF x =- 699 THEN
            exp_f := 1458;
        ELSIF x =- 698 THEN
            exp_f := 1458;
        ELSIF x =- 697 THEN
            exp_f := 1458;
        ELSIF x =- 696 THEN
            exp_f := 1458;
        ELSIF x =- 695 THEN
            exp_f := 1461;
        ELSIF x =- 694 THEN
            exp_f := 1461;
        ELSIF x =- 693 THEN
            exp_f := 1461;
        ELSIF x =- 692 THEN
            exp_f := 1461;
        ELSIF x =- 691 THEN
            exp_f := 1461;
        ELSIF x =- 690 THEN
            exp_f := 1464;
        ELSIF x =- 689 THEN
            exp_f := 1464;
        ELSIF x =- 688 THEN
            exp_f := 1464;
        ELSIF x =- 687 THEN
            exp_f := 1464;
        ELSIF x =- 686 THEN
            exp_f := 1467;
        ELSIF x =- 685 THEN
            exp_f := 1467;
        ELSIF x =- 684 THEN
            exp_f := 1467;
        ELSIF x =- 683 THEN
            exp_f := 1467;
        ELSIF x =- 682 THEN
            exp_f := 1470;
        ELSIF x =- 681 THEN
            exp_f := 1470;
        ELSIF x =- 680 THEN
            exp_f := 1470;
        ELSIF x =- 679 THEN
            exp_f := 1470;
        ELSIF x =- 678 THEN
            exp_f := 1473;
        ELSIF x =- 677 THEN
            exp_f := 1473;
        ELSIF x =- 676 THEN
            exp_f := 1473;
        ELSIF x =- 675 THEN
            exp_f := 1473;
        ELSIF x =- 674 THEN
            exp_f := 1476;
        ELSIF x =- 673 THEN
            exp_f := 1476;
        ELSIF x =- 672 THEN
            exp_f := 1476;
        ELSIF x =- 671 THEN
            exp_f := 1476;
        ELSIF x =- 670 THEN
            exp_f := 1479;
        ELSIF x =- 669 THEN
            exp_f := 1479;
        ELSIF x =- 668 THEN
            exp_f := 1479;
        ELSIF x =- 667 THEN
            exp_f := 1479;
        ELSIF x =- 666 THEN
            exp_f := 1482;
        ELSIF x =- 665 THEN
            exp_f := 1482;
        ELSIF x =- 664 THEN
            exp_f := 1482;
        ELSIF x =- 663 THEN
            exp_f := 1482;
        ELSIF x =- 662 THEN
            exp_f := 1482;
        ELSIF x =- 661 THEN
            exp_f := 1485;
        ELSIF x =- 660 THEN
            exp_f := 1485;
        ELSIF x =- 659 THEN
            exp_f := 1485;
        ELSIF x =- 658 THEN
            exp_f := 1485;
        ELSIF x =- 657 THEN
            exp_f := 1488;
        ELSIF x =- 656 THEN
            exp_f := 1488;
        ELSIF x =- 655 THEN
            exp_f := 1488;
        ELSIF x =- 654 THEN
            exp_f := 1488;
        ELSIF x =- 653 THEN
            exp_f := 1491;
        ELSIF x =- 652 THEN
            exp_f := 1491;
        ELSIF x =- 651 THEN
            exp_f := 1491;
        ELSIF x =- 650 THEN
            exp_f := 1491;
        ELSIF x =- 649 THEN
            exp_f := 1494;
        ELSIF x =- 648 THEN
            exp_f := 1494;
        ELSIF x =- 647 THEN
            exp_f := 1494;
        ELSIF x =- 646 THEN
            exp_f := 1494;
        ELSIF x =- 645 THEN
            exp_f := 1497;
        ELSIF x =- 644 THEN
            exp_f := 1497;
        ELSIF x =- 643 THEN
            exp_f := 1497;
        ELSIF x =- 642 THEN
            exp_f := 1497;
        ELSIF x =- 641 THEN
            exp_f := 1500;
        ELSIF x =- 640 THEN
            exp_f := 1500;
        ELSIF x =- 639 THEN
            exp_f := 1500;
        ELSIF x =- 638 THEN
            exp_f := 1500;
        ELSIF x =- 637 THEN
            exp_f := 1503;
        ELSIF x =- 636 THEN
            exp_f := 1503;
        ELSIF x =- 635 THEN
            exp_f := 1503;
        ELSIF x =- 634 THEN
            exp_f := 1503;
        ELSIF x =- 633 THEN
            exp_f := 1506;
        ELSIF x =- 632 THEN
            exp_f := 1506;
        ELSIF x =- 631 THEN
            exp_f := 1506;
        ELSIF x =- 630 THEN
            exp_f := 1506;
        ELSIF x =- 629 THEN
            exp_f := 1506;
        ELSIF x =- 628 THEN
            exp_f := 1509;
        ELSIF x =- 627 THEN
            exp_f := 1509;
        ELSIF x =- 626 THEN
            exp_f := 1509;
        ELSIF x =- 625 THEN
            exp_f := 1509;
        ELSIF x =- 624 THEN
            exp_f := 1512;
        ELSIF x =- 623 THEN
            exp_f := 1512;
        ELSIF x =- 622 THEN
            exp_f := 1512;
        ELSIF x =- 621 THEN
            exp_f := 1512;
        ELSIF x =- 620 THEN
            exp_f := 1515;
        ELSIF x =- 619 THEN
            exp_f := 1515;
        ELSIF x =- 618 THEN
            exp_f := 1515;
        ELSIF x =- 617 THEN
            exp_f := 1515;
        ELSIF x =- 616 THEN
            exp_f := 1518;
        ELSIF x =- 615 THEN
            exp_f := 1518;
        ELSIF x =- 614 THEN
            exp_f := 1518;
        ELSIF x =- 613 THEN
            exp_f := 1518;
        ELSIF x =- 612 THEN
            exp_f := 1521;
        ELSIF x =- 611 THEN
            exp_f := 1521;
        ELSIF x =- 610 THEN
            exp_f := 1521;
        ELSIF x =- 609 THEN
            exp_f := 1521;
        ELSIF x =- 608 THEN
            exp_f := 1524;
        ELSIF x =- 607 THEN
            exp_f := 1524;
        ELSIF x =- 606 THEN
            exp_f := 1524;
        ELSIF x =- 605 THEN
            exp_f := 1524;
        ELSIF x =- 604 THEN
            exp_f := 1527;
        ELSIF x =- 603 THEN
            exp_f := 1527;
        ELSIF x =- 602 THEN
            exp_f := 1527;
        ELSIF x =- 601 THEN
            exp_f := 1527;
        ELSIF x =- 600 THEN
            exp_f := 1527;
        ELSIF x =- 599 THEN
            exp_f := 1530;
        ELSIF x =- 598 THEN
            exp_f := 1530;
        ELSIF x =- 597 THEN
            exp_f := 1530;
        ELSIF x =- 596 THEN
            exp_f := 1530;
        ELSIF x =- 595 THEN
            exp_f := 1533;
        ELSIF x =- 594 THEN
            exp_f := 1533;
        ELSIF x =- 593 THEN
            exp_f := 1533;
        ELSIF x =- 592 THEN
            exp_f := 1533;
        ELSIF x =- 591 THEN
            exp_f := 1536;
        ELSIF x =- 590 THEN
            exp_f := 1536;
        ELSIF x =- 589 THEN
            exp_f := 1536;
        ELSIF x =- 588 THEN
            exp_f := 1536;
        ELSIF x =- 587 THEN
            exp_f := 1539;
        ELSIF x =- 586 THEN
            exp_f := 1539;
        ELSIF x =- 585 THEN
            exp_f := 1539;
        ELSIF x =- 584 THEN
            exp_f := 1539;
        ELSIF x =- 583 THEN
            exp_f := 1543;
        ELSIF x =- 582 THEN
            exp_f := 1543;
        ELSIF x =- 581 THEN
            exp_f := 1543;
        ELSIF x =- 580 THEN
            exp_f := 1543;
        ELSIF x =- 579 THEN
            exp_f := 1546;
        ELSIF x =- 578 THEN
            exp_f := 1546;
        ELSIF x =- 577 THEN
            exp_f := 1546;
        ELSIF x =- 576 THEN
            exp_f := 1546;
        ELSIF x =- 575 THEN
            exp_f := 1549;
        ELSIF x =- 574 THEN
            exp_f := 1549;
        ELSIF x =- 573 THEN
            exp_f := 1549;
        ELSIF x =- 572 THEN
            exp_f := 1549;
        ELSIF x =- 571 THEN
            exp_f := 1549;
        ELSIF x =- 570 THEN
            exp_f := 1552;
        ELSIF x =- 569 THEN
            exp_f := 1552;
        ELSIF x =- 568 THEN
            exp_f := 1552;
        ELSIF x =- 567 THEN
            exp_f := 1552;
        ELSIF x =- 566 THEN
            exp_f := 1555;
        ELSIF x =- 565 THEN
            exp_f := 1555;
        ELSIF x =- 564 THEN
            exp_f := 1555;
        ELSIF x =- 563 THEN
            exp_f := 1555;
        ELSIF x =- 562 THEN
            exp_f := 1558;
        ELSIF x =- 561 THEN
            exp_f := 1558;
        ELSIF x =- 560 THEN
            exp_f := 1558;
        ELSIF x =- 559 THEN
            exp_f := 1558;
        ELSIF x =- 558 THEN
            exp_f := 1561;
        ELSIF x =- 557 THEN
            exp_f := 1561;
        ELSIF x =- 556 THEN
            exp_f := 1561;
        ELSIF x =- 555 THEN
            exp_f := 1561;
        ELSIF x =- 554 THEN
            exp_f := 1564;
        ELSIF x =- 553 THEN
            exp_f := 1564;
        ELSIF x =- 552 THEN
            exp_f := 1564;
        ELSIF x =- 551 THEN
            exp_f := 1564;
        ELSIF x =- 550 THEN
            exp_f := 1567;
        ELSIF x =- 549 THEN
            exp_f := 1567;
        ELSIF x =- 548 THEN
            exp_f := 1567;
        ELSIF x =- 547 THEN
            exp_f := 1567;
        ELSIF x =- 546 THEN
            exp_f := 1570;
        ELSIF x =- 545 THEN
            exp_f := 1570;
        ELSIF x =- 544 THEN
            exp_f := 1570;
        ELSIF x =- 543 THEN
            exp_f := 1570;
        ELSIF x =- 542 THEN
            exp_f := 1570;
        ELSIF x =- 541 THEN
            exp_f := 1574;
        ELSIF x =- 540 THEN
            exp_f := 1574;
        ELSIF x =- 539 THEN
            exp_f := 1574;
        ELSIF x =- 538 THEN
            exp_f := 1574;
        ELSIF x =- 537 THEN
            exp_f := 1577;
        ELSIF x =- 536 THEN
            exp_f := 1577;
        ELSIF x =- 535 THEN
            exp_f := 1577;
        ELSIF x =- 534 THEN
            exp_f := 1577;
        ELSIF x =- 533 THEN
            exp_f := 1580;
        ELSIF x =- 532 THEN
            exp_f := 1580;
        ELSIF x =- 531 THEN
            exp_f := 1580;
        ELSIF x =- 530 THEN
            exp_f := 1580;
        ELSIF x =- 529 THEN
            exp_f := 1583;
        ELSIF x =- 528 THEN
            exp_f := 1583;
        ELSIF x =- 527 THEN
            exp_f := 1583;
        ELSIF x =- 526 THEN
            exp_f := 1583;
        ELSIF x =- 525 THEN
            exp_f := 1586;
        ELSIF x =- 524 THEN
            exp_f := 1586;
        ELSIF x =- 523 THEN
            exp_f := 1586;
        ELSIF x =- 522 THEN
            exp_f := 1586;
        ELSIF x =- 521 THEN
            exp_f := 1589;
        ELSIF x =- 520 THEN
            exp_f := 1589;
        ELSIF x =- 519 THEN
            exp_f := 1589;
        ELSIF x =- 518 THEN
            exp_f := 1589;
        ELSIF x =- 517 THEN
            exp_f := 1592;
        ELSIF x =- 516 THEN
            exp_f := 1592;
        ELSIF x =- 515 THEN
            exp_f := 1592;
        ELSIF x =- 514 THEN
            exp_f := 1592;
        ELSIF x =- 513 THEN
            exp_f := 1596;
        ELSIF x =- 512 THEN
            exp_f := 1596;
        ELSIF x =- 511 THEN
            exp_f := 1596;
        ELSIF x =- 510 THEN
            exp_f := 1596;
        ELSIF x =- 509 THEN
            exp_f := 1596;
        ELSIF x =- 508 THEN
            exp_f := 1596;
        ELSIF x =- 507 THEN
            exp_f := 1599;
        ELSIF x =- 506 THEN
            exp_f := 1599;
        ELSIF x =- 505 THEN
            exp_f := 1599;
        ELSIF x =- 504 THEN
            exp_f := 1599;
        ELSIF x =- 503 THEN
            exp_f := 1602;
        ELSIF x =- 502 THEN
            exp_f := 1602;
        ELSIF x =- 501 THEN
            exp_f := 1602;
        ELSIF x =- 500 THEN
            exp_f := 1602;
        ELSIF x =- 499 THEN
            exp_f := 1605;
        ELSIF x =- 498 THEN
            exp_f := 1605;
        ELSIF x =- 497 THEN
            exp_f := 1605;
        ELSIF x =- 496 THEN
            exp_f := 1605;
        ELSIF x =- 495 THEN
            exp_f := 1608;
        ELSIF x =- 494 THEN
            exp_f := 1608;
        ELSIF x =- 493 THEN
            exp_f := 1608;
        ELSIF x =- 492 THEN
            exp_f := 1608;
        ELSIF x =- 491 THEN
            exp_f := 1611;
        ELSIF x =- 490 THEN
            exp_f := 1611;
        ELSIF x =- 489 THEN
            exp_f := 1611;
        ELSIF x =- 488 THEN
            exp_f := 1611;
        ELSIF x =- 487 THEN
            exp_f := 1615;
        ELSIF x =- 486 THEN
            exp_f := 1615;
        ELSIF x =- 485 THEN
            exp_f := 1615;
        ELSIF x =- 484 THEN
            exp_f := 1615;
        ELSIF x =- 483 THEN
            exp_f := 1618;
        ELSIF x =- 482 THEN
            exp_f := 1618;
        ELSIF x =- 481 THEN
            exp_f := 1618;
        ELSIF x =- 480 THEN
            exp_f := 1618;
        ELSIF x =- 479 THEN
            exp_f := 1621;
        ELSIF x =- 478 THEN
            exp_f := 1621;
        ELSIF x =- 477 THEN
            exp_f := 1621;
        ELSIF x =- 476 THEN
            exp_f := 1621;
        ELSIF x =- 475 THEN
            exp_f := 1624;
        ELSIF x =- 474 THEN
            exp_f := 1624;
        ELSIF x =- 473 THEN
            exp_f := 1624;
        ELSIF x =- 472 THEN
            exp_f := 1624;
        ELSIF x =- 471 THEN
            exp_f := 1627;
        ELSIF x =- 470 THEN
            exp_f := 1627;
        ELSIF x =- 469 THEN
            exp_f := 1627;
        ELSIF x =- 468 THEN
            exp_f := 1627;
        ELSIF x =- 467 THEN
            exp_f := 1631;
        ELSIF x =- 466 THEN
            exp_f := 1631;
        ELSIF x =- 465 THEN
            exp_f := 1631;
        ELSIF x =- 464 THEN
            exp_f := 1631;
        ELSIF x =- 463 THEN
            exp_f := 1634;
        ELSIF x =- 462 THEN
            exp_f := 1634;
        ELSIF x =- 461 THEN
            exp_f := 1634;
        ELSIF x =- 460 THEN
            exp_f := 1634;
        ELSIF x =- 459 THEN
            exp_f := 1637;
        ELSIF x =- 458 THEN
            exp_f := 1637;
        ELSIF x =- 457 THEN
            exp_f := 1637;
        ELSIF x =- 456 THEN
            exp_f := 1637;
        ELSIF x =- 455 THEN
            exp_f := 1640;
        ELSIF x =- 454 THEN
            exp_f := 1640;
        ELSIF x =- 453 THEN
            exp_f := 1640;
        ELSIF x =- 452 THEN
            exp_f := 1640;
        ELSIF x =- 451 THEN
            exp_f := 1644;
        ELSIF x =- 450 THEN
            exp_f := 1644;
        ELSIF x =- 449 THEN
            exp_f := 1644;
        ELSIF x =- 448 THEN
            exp_f := 1644;
        ELSIF x =- 447 THEN
            exp_f := 1647;
        ELSIF x =- 446 THEN
            exp_f := 1647;
        ELSIF x =- 445 THEN
            exp_f := 1647;
        ELSIF x =- 444 THEN
            exp_f := 1647;
        ELSIF x =- 443 THEN
            exp_f := 1650;
        ELSIF x =- 442 THEN
            exp_f := 1650;
        ELSIF x =- 441 THEN
            exp_f := 1650;
        ELSIF x =- 440 THEN
            exp_f := 1650;
        ELSIF x =- 439 THEN
            exp_f := 1653;
        ELSIF x =- 438 THEN
            exp_f := 1653;
        ELSIF x =- 437 THEN
            exp_f := 1653;
        ELSIF x =- 436 THEN
            exp_f := 1653;
        ELSIF x =- 435 THEN
            exp_f := 1657;
        ELSIF x =- 434 THEN
            exp_f := 1657;
        ELSIF x =- 433 THEN
            exp_f := 1657;
        ELSIF x =- 432 THEN
            exp_f := 1657;
        ELSIF x =- 431 THEN
            exp_f := 1660;
        ELSIF x =- 430 THEN
            exp_f := 1660;
        ELSIF x =- 429 THEN
            exp_f := 1660;
        ELSIF x =- 428 THEN
            exp_f := 1660;
        ELSIF x =- 427 THEN
            exp_f := 1663;
        ELSIF x =- 426 THEN
            exp_f := 1663;
        ELSIF x =- 425 THEN
            exp_f := 1663;
        ELSIF x =- 424 THEN
            exp_f := 1663;
        ELSIF x =- 423 THEN
            exp_f := 1667;
        ELSIF x =- 422 THEN
            exp_f := 1667;
        ELSIF x =- 421 THEN
            exp_f := 1667;
        ELSIF x =- 420 THEN
            exp_f := 1667;
        ELSIF x =- 419 THEN
            exp_f := 1670;
        ELSIF x =- 418 THEN
            exp_f := 1670;
        ELSIF x =- 417 THEN
            exp_f := 1670;
        ELSIF x =- 416 THEN
            exp_f := 1670;
        ELSIF x =- 415 THEN
            exp_f := 1673;
        ELSIF x =- 414 THEN
            exp_f := 1673;
        ELSIF x =- 413 THEN
            exp_f := 1673;
        ELSIF x =- 412 THEN
            exp_f := 1673;
        ELSIF x =- 411 THEN
            exp_f := 1676;
        ELSIF x =- 410 THEN
            exp_f := 1676;
        ELSIF x =- 409 THEN
            exp_f := 1676;
        ELSIF x =- 408 THEN
            exp_f := 1676;
        ELSIF x =- 407 THEN
            exp_f := 1680;
        ELSIF x =- 406 THEN
            exp_f := 1680;
        ELSIF x =- 405 THEN
            exp_f := 1680;
        ELSIF x =- 404 THEN
            exp_f := 1680;
        ELSIF x =- 403 THEN
            exp_f := 1683;
        ELSIF x =- 402 THEN
            exp_f := 1683;
        ELSIF x =- 401 THEN
            exp_f := 1683;
        ELSIF x =- 400 THEN
            exp_f := 1683;
        ELSIF x =- 399 THEN
            exp_f := 1686;
        ELSIF x =- 398 THEN
            exp_f := 1686;
        ELSIF x =- 397 THEN
            exp_f := 1686;
        ELSIF x =- 396 THEN
            exp_f := 1686;
        ELSIF x =- 395 THEN
            exp_f := 1690;
        ELSIF x =- 394 THEN
            exp_f := 1690;
        ELSIF x =- 393 THEN
            exp_f := 1690;
        ELSIF x =- 392 THEN
            exp_f := 1690;
        ELSIF x =- 391 THEN
            exp_f := 1693;
        ELSIF x =- 390 THEN
            exp_f := 1693;
        ELSIF x =- 389 THEN
            exp_f := 1693;
        ELSIF x =- 388 THEN
            exp_f := 1693;
        ELSIF x =- 387 THEN
            exp_f := 1696;
        ELSIF x =- 386 THEN
            exp_f := 1696;
        ELSIF x =- 385 THEN
            exp_f := 1696;
        ELSIF x =- 384 THEN
            exp_f := 1696;
        ELSIF x =- 383 THEN
            exp_f := 1700;
        ELSIF x =- 382 THEN
            exp_f := 1700;
        ELSIF x =- 381 THEN
            exp_f := 1700;
        ELSIF x =- 380 THEN
            exp_f := 1700;
        ELSIF x =- 379 THEN
            exp_f := 1703;
        ELSIF x =- 378 THEN
            exp_f := 1703;
        ELSIF x =- 377 THEN
            exp_f := 1703;
        ELSIF x =- 376 THEN
            exp_f := 1703;
        ELSIF x =- 375 THEN
            exp_f := 1706;
        ELSIF x =- 374 THEN
            exp_f := 1706;
        ELSIF x =- 373 THEN
            exp_f := 1706;
        ELSIF x =- 372 THEN
            exp_f := 1706;
        ELSIF x =- 371 THEN
            exp_f := 1710;
        ELSIF x =- 370 THEN
            exp_f := 1710;
        ELSIF x =- 369 THEN
            exp_f := 1710;
        ELSIF x =- 368 THEN
            exp_f := 1710;
        ELSIF x =- 367 THEN
            exp_f := 1713;
        ELSIF x =- 366 THEN
            exp_f := 1713;
        ELSIF x =- 365 THEN
            exp_f := 1713;
        ELSIF x =- 364 THEN
            exp_f := 1713;
        ELSIF x =- 363 THEN
            exp_f := 1717;
        ELSIF x =- 362 THEN
            exp_f := 1717;
        ELSIF x =- 361 THEN
            exp_f := 1717;
        ELSIF x =- 360 THEN
            exp_f := 1717;
        ELSIF x =- 359 THEN
            exp_f := 1720;
        ELSIF x =- 358 THEN
            exp_f := 1720;
        ELSIF x =- 357 THEN
            exp_f := 1720;
        ELSIF x =- 356 THEN
            exp_f := 1720;
        ELSIF x =- 355 THEN
            exp_f := 1723;
        ELSIF x =- 354 THEN
            exp_f := 1723;
        ELSIF x =- 353 THEN
            exp_f := 1723;
        ELSIF x =- 352 THEN
            exp_f := 1723;
        ELSIF x =- 351 THEN
            exp_f := 1727;
        ELSIF x =- 350 THEN
            exp_f := 1727;
        ELSIF x =- 349 THEN
            exp_f := 1727;
        ELSIF x =- 348 THEN
            exp_f := 1727;
        ELSIF x =- 347 THEN
            exp_f := 1730;
        ELSIF x =- 346 THEN
            exp_f := 1730;
        ELSIF x =- 345 THEN
            exp_f := 1730;
        ELSIF x =- 344 THEN
            exp_f := 1730;
        ELSIF x =- 343 THEN
            exp_f := 1734;
        ELSIF x =- 342 THEN
            exp_f := 1734;
        ELSIF x =- 341 THEN
            exp_f := 1734;
        ELSIF x =- 340 THEN
            exp_f := 1734;
        ELSIF x =- 339 THEN
            exp_f := 1737;
        ELSIF x =- 338 THEN
            exp_f := 1737;
        ELSIF x =- 337 THEN
            exp_f := 1737;
        ELSIF x =- 336 THEN
            exp_f := 1737;
        ELSIF x =- 335 THEN
            exp_f := 1740;
        ELSIF x =- 334 THEN
            exp_f := 1740;
        ELSIF x =- 333 THEN
            exp_f := 1740;
        ELSIF x =- 332 THEN
            exp_f := 1740;
        ELSIF x =- 331 THEN
            exp_f := 1744;
        ELSIF x =- 330 THEN
            exp_f := 1744;
        ELSIF x =- 329 THEN
            exp_f := 1744;
        ELSIF x =- 328 THEN
            exp_f := 1744;
        ELSIF x =- 327 THEN
            exp_f := 1747;
        ELSIF x =- 326 THEN
            exp_f := 1747;
        ELSIF x =- 325 THEN
            exp_f := 1747;
        ELSIF x =- 324 THEN
            exp_f := 1747;
        ELSIF x =- 323 THEN
            exp_f := 1751;
        ELSIF x =- 322 THEN
            exp_f := 1751;
        ELSIF x =- 321 THEN
            exp_f := 1751;
        ELSIF x =- 320 THEN
            exp_f := 1751;
        ELSIF x =- 319 THEN
            exp_f := 1754;
        ELSIF x =- 318 THEN
            exp_f := 1754;
        ELSIF x =- 317 THEN
            exp_f := 1754;
        ELSIF x =- 316 THEN
            exp_f := 1754;
        ELSIF x =- 315 THEN
            exp_f := 1758;
        ELSIF x =- 314 THEN
            exp_f := 1758;
        ELSIF x =- 313 THEN
            exp_f := 1758;
        ELSIF x =- 312 THEN
            exp_f := 1758;
        ELSIF x =- 311 THEN
            exp_f := 1761;
        ELSIF x =- 310 THEN
            exp_f := 1761;
        ELSIF x =- 309 THEN
            exp_f := 1761;
        ELSIF x =- 308 THEN
            exp_f := 1761;
        ELSIF x =- 307 THEN
            exp_f := 1765;
        ELSIF x =- 306 THEN
            exp_f := 1765;
        ELSIF x =- 305 THEN
            exp_f := 1765;
        ELSIF x =- 304 THEN
            exp_f := 1765;
        ELSIF x =- 303 THEN
            exp_f := 1768;
        ELSIF x =- 302 THEN
            exp_f := 1768;
        ELSIF x =- 301 THEN
            exp_f := 1768;
        ELSIF x =- 300 THEN
            exp_f := 1768;
        ELSIF x =- 299 THEN
            exp_f := 1771;
        ELSIF x =- 298 THEN
            exp_f := 1771;
        ELSIF x =- 297 THEN
            exp_f := 1771;
        ELSIF x =- 296 THEN
            exp_f := 1771;
        ELSIF x =- 295 THEN
            exp_f := 1775;
        ELSIF x =- 294 THEN
            exp_f := 1775;
        ELSIF x =- 293 THEN
            exp_f := 1775;
        ELSIF x =- 292 THEN
            exp_f := 1775;
        ELSIF x =- 291 THEN
            exp_f := 1778;
        ELSIF x =- 290 THEN
            exp_f := 1778;
        ELSIF x =- 289 THEN
            exp_f := 1778;
        ELSIF x =- 288 THEN
            exp_f := 1778;
        ELSIF x =- 287 THEN
            exp_f := 1782;
        ELSIF x =- 286 THEN
            exp_f := 1782;
        ELSIF x =- 285 THEN
            exp_f := 1782;
        ELSIF x =- 284 THEN
            exp_f := 1782;
        ELSIF x =- 283 THEN
            exp_f := 1785;
        ELSIF x =- 282 THEN
            exp_f := 1785;
        ELSIF x =- 281 THEN
            exp_f := 1785;
        ELSIF x =- 280 THEN
            exp_f := 1785;
        ELSIF x =- 279 THEN
            exp_f := 1789;
        ELSIF x =- 278 THEN
            exp_f := 1789;
        ELSIF x =- 277 THEN
            exp_f := 1789;
        ELSIF x =- 276 THEN
            exp_f := 1789;
        ELSIF x =- 275 THEN
            exp_f := 1792;
        ELSIF x =- 274 THEN
            exp_f := 1792;
        ELSIF x =- 273 THEN
            exp_f := 1792;
        ELSIF x =- 272 THEN
            exp_f := 1792;
        ELSIF x =- 271 THEN
            exp_f := 1796;
        ELSIF x =- 270 THEN
            exp_f := 1796;
        ELSIF x =- 269 THEN
            exp_f := 1796;
        ELSIF x =- 268 THEN
            exp_f := 1796;
        ELSIF x =- 267 THEN
            exp_f := 1799;
        ELSIF x =- 266 THEN
            exp_f := 1799;
        ELSIF x =- 265 THEN
            exp_f := 1799;
        ELSIF x =- 264 THEN
            exp_f := 1799;
        ELSIF x =- 263 THEN
            exp_f := 1803;
        ELSIF x =- 262 THEN
            exp_f := 1803;
        ELSIF x =- 261 THEN
            exp_f := 1803;
        ELSIF x =- 260 THEN
            exp_f := 1803;
        ELSIF x =- 259 THEN
            exp_f := 1807;
        ELSIF x =- 258 THEN
            exp_f := 1807;
        ELSIF x =- 257 THEN
            exp_f := 1807;
        ELSIF x =- 256 THEN
            exp_f := 1807;
        ELSIF x =- 255 THEN
            exp_f := 1810;
        ELSIF x =- 254 THEN
            exp_f := 1810;
        ELSIF x =- 253 THEN
            exp_f := 1810;
        ELSIF x =- 252 THEN
            exp_f := 1810;
        ELSIF x =- 251 THEN
            exp_f := 1814;
        ELSIF x =- 250 THEN
            exp_f := 1814;
        ELSIF x =- 249 THEN
            exp_f := 1814;
        ELSIF x =- 248 THEN
            exp_f := 1814;
        ELSIF x =- 247 THEN
            exp_f := 1817;
        ELSIF x =- 246 THEN
            exp_f := 1817;
        ELSIF x =- 245 THEN
            exp_f := 1817;
        ELSIF x =- 244 THEN
            exp_f := 1817;
        ELSIF x =- 243 THEN
            exp_f := 1821;
        ELSIF x =- 242 THEN
            exp_f := 1821;
        ELSIF x =- 241 THEN
            exp_f := 1821;
        ELSIF x =- 240 THEN
            exp_f := 1821;
        ELSIF x =- 239 THEN
            exp_f := 1824;
        ELSIF x =- 238 THEN
            exp_f := 1824;
        ELSIF x =- 237 THEN
            exp_f := 1824;
        ELSIF x =- 236 THEN
            exp_f := 1824;
        ELSIF x =- 235 THEN
            exp_f := 1828;
        ELSIF x =- 234 THEN
            exp_f := 1828;
        ELSIF x =- 233 THEN
            exp_f := 1828;
        ELSIF x =- 232 THEN
            exp_f := 1828;
        ELSIF x =- 231 THEN
            exp_f := 1832;
        ELSIF x =- 230 THEN
            exp_f := 1832;
        ELSIF x =- 229 THEN
            exp_f := 1832;
        ELSIF x =- 228 THEN
            exp_f := 1832;
        ELSIF x =- 227 THEN
            exp_f := 1835;
        ELSIF x =- 226 THEN
            exp_f := 1835;
        ELSIF x =- 225 THEN
            exp_f := 1835;
        ELSIF x =- 224 THEN
            exp_f := 1835;
        ELSIF x =- 223 THEN
            exp_f := 1839;
        ELSIF x =- 222 THEN
            exp_f := 1839;
        ELSIF x =- 221 THEN
            exp_f := 1839;
        ELSIF x =- 220 THEN
            exp_f := 1839;
        ELSIF x =- 219 THEN
            exp_f := 1842;
        ELSIF x =- 218 THEN
            exp_f := 1842;
        ELSIF x =- 217 THEN
            exp_f := 1842;
        ELSIF x =- 216 THEN
            exp_f := 1842;
        ELSIF x =- 215 THEN
            exp_f := 1846;
        ELSIF x =- 214 THEN
            exp_f := 1846;
        ELSIF x =- 213 THEN
            exp_f := 1846;
        ELSIF x =- 212 THEN
            exp_f := 1846;
        ELSIF x =- 211 THEN
            exp_f := 1850;
        ELSIF x =- 210 THEN
            exp_f := 1850;
        ELSIF x =- 209 THEN
            exp_f := 1850;
        ELSIF x =- 208 THEN
            exp_f := 1850;
        ELSIF x =- 207 THEN
            exp_f := 1853;
        ELSIF x =- 206 THEN
            exp_f := 1853;
        ELSIF x =- 205 THEN
            exp_f := 1853;
        ELSIF x =- 204 THEN
            exp_f := 1853;
        ELSIF x =- 203 THEN
            exp_f := 1857;
        ELSIF x =- 202 THEN
            exp_f := 1857;
        ELSIF x =- 201 THEN
            exp_f := 1857;
        ELSIF x =- 200 THEN
            exp_f := 1857;
        ELSIF x =- 199 THEN
            exp_f := 1860;
        ELSIF x =- 198 THEN
            exp_f := 1860;
        ELSIF x =- 197 THEN
            exp_f := 1860;
        ELSIF x =- 196 THEN
            exp_f := 1860;
        ELSIF x =- 195 THEN
            exp_f := 1864;
        ELSIF x =- 194 THEN
            exp_f := 1864;
        ELSIF x =- 193 THEN
            exp_f := 1864;
        ELSIF x =- 192 THEN
            exp_f := 1864;
        ELSIF x =- 191 THEN
            exp_f := 1868;
        ELSIF x =- 190 THEN
            exp_f := 1868;
        ELSIF x =- 189 THEN
            exp_f := 1868;
        ELSIF x =- 188 THEN
            exp_f := 1868;
        ELSIF x =- 187 THEN
            exp_f := 1871;
        ELSIF x =- 186 THEN
            exp_f := 1871;
        ELSIF x =- 185 THEN
            exp_f := 1871;
        ELSIF x =- 184 THEN
            exp_f := 1871;
        ELSIF x =- 183 THEN
            exp_f := 1875;
        ELSIF x =- 182 THEN
            exp_f := 1875;
        ELSIF x =- 181 THEN
            exp_f := 1875;
        ELSIF x =- 180 THEN
            exp_f := 1875;
        ELSIF x =- 179 THEN
            exp_f := 1879;
        ELSIF x =- 178 THEN
            exp_f := 1879;
        ELSIF x =- 177 THEN
            exp_f := 1879;
        ELSIF x =- 176 THEN
            exp_f := 1879;
        ELSIF x =- 175 THEN
            exp_f := 1882;
        ELSIF x =- 174 THEN
            exp_f := 1882;
        ELSIF x =- 173 THEN
            exp_f := 1882;
        ELSIF x =- 172 THEN
            exp_f := 1882;
        ELSIF x =- 171 THEN
            exp_f := 1886;
        ELSIF x =- 170 THEN
            exp_f := 1886;
        ELSIF x =- 169 THEN
            exp_f := 1886;
        ELSIF x =- 168 THEN
            exp_f := 1886;
        ELSIF x =- 167 THEN
            exp_f := 1890;
        ELSIF x =- 166 THEN
            exp_f := 1890;
        ELSIF x =- 165 THEN
            exp_f := 1890;
        ELSIF x =- 164 THEN
            exp_f := 1890;
        ELSIF x =- 163 THEN
            exp_f := 1894;
        ELSIF x =- 162 THEN
            exp_f := 1894;
        ELSIF x =- 161 THEN
            exp_f := 1894;
        ELSIF x =- 160 THEN
            exp_f := 1894;
        ELSIF x =- 159 THEN
            exp_f := 1897;
        ELSIF x =- 158 THEN
            exp_f := 1897;
        ELSIF x =- 157 THEN
            exp_f := 1897;
        ELSIF x =- 156 THEN
            exp_f := 1897;
        ELSIF x =- 155 THEN
            exp_f := 1901;
        ELSIF x =- 154 THEN
            exp_f := 1901;
        ELSIF x =- 153 THEN
            exp_f := 1901;
        ELSIF x =- 152 THEN
            exp_f := 1901;
        ELSIF x =- 151 THEN
            exp_f := 1905;
        ELSIF x =- 150 THEN
            exp_f := 1905;
        ELSIF x =- 149 THEN
            exp_f := 1905;
        ELSIF x =- 148 THEN
            exp_f := 1905;
        ELSIF x =- 147 THEN
            exp_f := 1908;
        ELSIF x =- 146 THEN
            exp_f := 1908;
        ELSIF x =- 145 THEN
            exp_f := 1908;
        ELSIF x =- 144 THEN
            exp_f := 1908;
        ELSIF x =- 143 THEN
            exp_f := 1912;
        ELSIF x =- 142 THEN
            exp_f := 1912;
        ELSIF x =- 141 THEN
            exp_f := 1912;
        ELSIF x =- 140 THEN
            exp_f := 1912;
        ELSIF x =- 139 THEN
            exp_f := 1916;
        ELSIF x =- 138 THEN
            exp_f := 1916;
        ELSIF x =- 137 THEN
            exp_f := 1916;
        ELSIF x =- 136 THEN
            exp_f := 1916;
        ELSIF x =- 135 THEN
            exp_f := 1920;
        ELSIF x =- 134 THEN
            exp_f := 1920;
        ELSIF x =- 133 THEN
            exp_f := 1920;
        ELSIF x =- 132 THEN
            exp_f := 1920;
        ELSIF x =- 131 THEN
            exp_f := 1923;
        ELSIF x =- 130 THEN
            exp_f := 1923;
        ELSIF x =- 129 THEN
            exp_f := 1923;
        ELSIF x =- 128 THEN
            exp_f := 1923;
        ELSIF x =- 127 THEN
            exp_f := 1927;
        ELSIF x =- 126 THEN
            exp_f := 1927;
        ELSIF x =- 125 THEN
            exp_f := 1927;
        ELSIF x =- 124 THEN
            exp_f := 1927;
        ELSIF x =- 123 THEN
            exp_f := 1931;
        ELSIF x =- 122 THEN
            exp_f := 1931;
        ELSIF x =- 121 THEN
            exp_f := 1931;
        ELSIF x =- 120 THEN
            exp_f := 1931;
        ELSIF x =- 119 THEN
            exp_f := 1935;
        ELSIF x =- 118 THEN
            exp_f := 1935;
        ELSIF x =- 117 THEN
            exp_f := 1935;
        ELSIF x =- 116 THEN
            exp_f := 1935;
        ELSIF x =- 115 THEN
            exp_f := 1938;
        ELSIF x =- 114 THEN
            exp_f := 1938;
        ELSIF x =- 113 THEN
            exp_f := 1938;
        ELSIF x =- 112 THEN
            exp_f := 1938;
        ELSIF x =- 111 THEN
            exp_f := 1942;
        ELSIF x =- 110 THEN
            exp_f := 1942;
        ELSIF x =- 109 THEN
            exp_f := 1942;
        ELSIF x =- 108 THEN
            exp_f := 1942;
        ELSIF x =- 107 THEN
            exp_f := 1946;
        ELSIF x =- 106 THEN
            exp_f := 1946;
        ELSIF x =- 105 THEN
            exp_f := 1946;
        ELSIF x =- 104 THEN
            exp_f := 1946;
        ELSIF x =- 103 THEN
            exp_f := 1950;
        ELSIF x =- 102 THEN
            exp_f := 1950;
        ELSIF x =- 101 THEN
            exp_f := 1950;
        ELSIF x =- 100 THEN
            exp_f := 1950;
        ELSIF x =- 99 THEN
            exp_f := 1954;
        ELSIF x =- 98 THEN
            exp_f := 1954;
        ELSIF x =- 97 THEN
            exp_f := 1954;
        ELSIF x =- 96 THEN
            exp_f := 1954;
        ELSIF x =- 95 THEN
            exp_f := 1958;
        ELSIF x =- 94 THEN
            exp_f := 1958;
        ELSIF x =- 93 THEN
            exp_f := 1958;
        ELSIF x =- 92 THEN
            exp_f := 1958;
        ELSIF x =- 91 THEN
            exp_f := 1961;
        ELSIF x =- 90 THEN
            exp_f := 1961;
        ELSIF x =- 89 THEN
            exp_f := 1961;
        ELSIF x =- 88 THEN
            exp_f := 1961;
        ELSIF x =- 87 THEN
            exp_f := 1965;
        ELSIF x =- 86 THEN
            exp_f := 1965;
        ELSIF x =- 85 THEN
            exp_f := 1965;
        ELSIF x =- 84 THEN
            exp_f := 1965;
        ELSIF x =- 83 THEN
            exp_f := 1969;
        ELSIF x =- 82 THEN
            exp_f := 1969;
        ELSIF x =- 81 THEN
            exp_f := 1969;
        ELSIF x =- 80 THEN
            exp_f := 1969;
        ELSIF x =- 79 THEN
            exp_f := 1973;
        ELSIF x =- 78 THEN
            exp_f := 1973;
        ELSIF x =- 77 THEN
            exp_f := 1973;
        ELSIF x =- 76 THEN
            exp_f := 1973;
        ELSIF x =- 75 THEN
            exp_f := 1977;
        ELSIF x =- 74 THEN
            exp_f := 1977;
        ELSIF x =- 73 THEN
            exp_f := 1977;
        ELSIF x =- 72 THEN
            exp_f := 1977;
        ELSIF x =- 71 THEN
            exp_f := 1981;
        ELSIF x =- 70 THEN
            exp_f := 1981;
        ELSIF x =- 69 THEN
            exp_f := 1981;
        ELSIF x =- 68 THEN
            exp_f := 1981;
        ELSIF x =- 67 THEN
            exp_f := 1984;
        ELSIF x =- 66 THEN
            exp_f := 1984;
        ELSIF x =- 65 THEN
            exp_f := 1984;
        ELSIF x =- 64 THEN
            exp_f := 1984;
        ELSIF x =- 63 THEN
            exp_f := 1988;
        ELSIF x =- 62 THEN
            exp_f := 1988;
        ELSIF x =- 61 THEN
            exp_f := 1988;
        ELSIF x =- 60 THEN
            exp_f := 1988;
        ELSIF x =- 59 THEN
            exp_f := 1992;
        ELSIF x =- 58 THEN
            exp_f := 1992;
        ELSIF x =- 57 THEN
            exp_f := 1992;
        ELSIF x =- 56 THEN
            exp_f := 1992;
        ELSIF x =- 55 THEN
            exp_f := 1996;
        ELSIF x =- 54 THEN
            exp_f := 1996;
        ELSIF x =- 53 THEN
            exp_f := 1996;
        ELSIF x =- 52 THEN
            exp_f := 1996;
        ELSIF x =- 51 THEN
            exp_f := 2000;
        ELSIF x =- 50 THEN
            exp_f := 2000;
        ELSIF x =- 49 THEN
            exp_f := 2000;
        ELSIF x =- 48 THEN
            exp_f := 2000;
        ELSIF x =- 47 THEN
            exp_f := 2004;
        ELSIF x =- 46 THEN
            exp_f := 2004;
        ELSIF x =- 45 THEN
            exp_f := 2004;
        ELSIF x =- 44 THEN
            exp_f := 2004;
        ELSIF x =- 43 THEN
            exp_f := 2008;
        ELSIF x =- 42 THEN
            exp_f := 2008;
        ELSIF x =- 41 THEN
            exp_f := 2008;
        ELSIF x =- 40 THEN
            exp_f := 2008;
        ELSIF x =- 39 THEN
            exp_f := 2012;
        ELSIF x =- 38 THEN
            exp_f := 2012;
        ELSIF x =- 37 THEN
            exp_f := 2012;
        ELSIF x =- 36 THEN
            exp_f := 2012;
        ELSIF x =- 35 THEN
            exp_f := 2016;
        ELSIF x =- 34 THEN
            exp_f := 2016;
        ELSIF x =- 33 THEN
            exp_f := 2016;
        ELSIF x =- 32 THEN
            exp_f := 2016;
        ELSIF x =- 31 THEN
            exp_f := 2020;
        ELSIF x =- 30 THEN
            exp_f := 2020;
        ELSIF x =- 29 THEN
            exp_f := 2020;
        ELSIF x =- 28 THEN
            exp_f := 2020;
        ELSIF x =- 27 THEN
            exp_f := 2024;
        ELSIF x =- 26 THEN
            exp_f := 2024;
        ELSIF x =- 25 THEN
            exp_f := 2024;
        ELSIF x =- 24 THEN
            exp_f := 2024;
        ELSIF x =- 23 THEN
            exp_f := 2028;
        ELSIF x =- 22 THEN
            exp_f := 2028;
        ELSIF x =- 21 THEN
            exp_f := 2028;
        ELSIF x =- 20 THEN
            exp_f := 2028;
        ELSIF x =- 19 THEN
            exp_f := 2032;
        ELSIF x =- 18 THEN
            exp_f := 2032;
        ELSIF x =- 17 THEN
            exp_f := 2032;
        ELSIF x =- 16 THEN
            exp_f := 2032;
        ELSIF x =- 15 THEN
            exp_f := 2036;
        ELSIF x =- 14 THEN
            exp_f := 2036;
        ELSIF x =- 13 THEN
            exp_f := 2036;
        ELSIF x =- 12 THEN
            exp_f := 2036;
        ELSIF x =- 11 THEN
            exp_f := 2040;
        ELSIF x =- 10 THEN
            exp_f := 2040;
        ELSIF x =- 9 THEN
            exp_f := 2040;
        ELSIF x =- 8 THEN
            exp_f := 2040;
        ELSIF x =- 7 THEN
            exp_f := 2044;
        ELSIF x =- 6 THEN
            exp_f := 2044;
        ELSIF x =- 5 THEN
            exp_f := 2044;
        ELSIF x =- 4 THEN
            exp_f := 2044;
        ELSIF x =- 3 THEN
            exp_f := 2048;
        ELSIF x =- 2 THEN
            exp_f := 2048;
        ELSIF x =- 1 THEN
            exp_f := 2048;
        ELSIF x = 0 THEN
            exp_f := 2048;
        ELSIF x >= 1 THEN
            exp_f := 2048;
        END IF;
        RETURN exp_f;
    END;
END PACKAGE BODY exp_pkg;