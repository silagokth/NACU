-------------------------------------------------------
--! @file sigmoid_pkg.vhd
--! @brief Look up package for sigmoid (matlab generated)
--! @details 
--! @author Guido Baccelli
--! @version 1.0
--! @date 23/08/2019
--! @bug NONE
--! @todo NONE
--! @copyright  GNU Public License [GPL-3.0].
-------------------------------------------------------
---------------- Copyright (c) notice -----------------------------------------
--
-- The VHDL code, the logic and concepts described in this file constitute
-- the intellectual property of the authors listed below, who are affiliated
-- to KTH(Kungliga Tekniska Högskolan), School of ICT, Kista.
-- Any unauthorised use, copy or distribution is strictly prohibited.
-- Any authorised use, copy or distribution should carry this copyright notice
-- unaltered.
-------------------------------------------------------------------------------
-- Title      : Look up package for sigmoid (matlab generated)
-- Project    : SiLago
-------------------------------------------------------------------------------
-- File       : sigmoid_pkg.vhd
-- Author     : Guido Baccelli
-- Company    : KTH
-- Created    : 23/08/2019
-- Last update: 23/08/2019
-- Platform   : SiLago
-- Standard   : VHDL'08
-- Supervisor : Dimitrios Stathis
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Contact    : Dimitrios Stathis <stathis@kth.se>
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author                  Description
-- 23/08/2019  1.0      Guido Baccelli          Created
-------------------------------------------------------------------------------

--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#
--                                                                         #
--This file is part of SiLago.                                             #
--                                                                         #
--    SiLago platform source code is distributed freely: you can           #
--    redistribute it and/or modify it under the terms of the GNU          #
--    General Public License as published by the Free Software Foundation, #
--    either version 3 of the License, or (at your option) any             #
--    later version.                                                       #
--                                                                         #
--    SiLago is distributed in the hope that it will be useful,            #
--    but WITHOUT ANY WARRANTY; without even the implied warranty of       #
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the        #
--    GNU General Public License for more details.                         #
--                                                                         #
--    You should have received a copy of the GNU General Public License    #
--    along with SiLago.  If not, see <https://www.gnu.org/licenses/>.     #
--                                                                         #
--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#

--! Standard ieee library
LIBRARY ieee;
--! Default working library
LIBRARY work;
--! Standard logic package
USE ieee.std_logic_1164.ALL;
--! Standard numeric package for signed and unsigned
USE ieee.numeric_std.ALL;

--! @brief Package file with Sigmoid behavior model for testbench
--! @details The only content is the 'sigmoid_fp11' function that emulates behavior of Sigmoid operation inside 'NACU'
PACKAGE sigmoid_pkg IS

    FUNCTION sigmoid_fp11(
        x : INTEGER
    ) RETURN INTEGER;

END PACKAGE sigmoid_pkg;

--! @brief Contains body of function 'sigmoid_fp11'
--! @details The function 'sigmoid_fp11' (and the testbench) interpret input and output data words
--! as integer values instead of fixed-point values. This makes the model easier to describe.
--! The function describes the Sigmoid by assigning the corresponding output to each possible
--! input value representable on Q4.11.
PACKAGE BODY sigmoid_pkg IS
    FUNCTION sigmoid_fp11(
        x : INTEGER)
        RETURN INTEGER IS
        VARIABLE sigmoid_f : INTEGER;
    BEGIN
        IF x <= - 16896 THEN
            sigmoid_f := 0;
        ELSIF x =- 16895 THEN
            sigmoid_f := 1;
        ELSIF x =- 16894 THEN
            sigmoid_f := 1;
        ELSIF x =- 16893 THEN
            sigmoid_f := 1;
        ELSIF x =- 16892 THEN
            sigmoid_f := 1;
        ELSIF x =- 16891 THEN
            sigmoid_f := 1;
        ELSIF x =- 16890 THEN
            sigmoid_f := 1;
        ELSIF x =- 16889 THEN
            sigmoid_f := 1;
        ELSIF x =- 16888 THEN
            sigmoid_f := 1;
        ELSIF x =- 16887 THEN
            sigmoid_f := 1;
        ELSIF x =- 16886 THEN
            sigmoid_f := 1;
        ELSIF x =- 16885 THEN
            sigmoid_f := 1;
        ELSIF x =- 16884 THEN
            sigmoid_f := 1;
        ELSIF x =- 16883 THEN
            sigmoid_f := 1;
        ELSIF x =- 16882 THEN
            sigmoid_f := 1;
        ELSIF x =- 16881 THEN
            sigmoid_f := 1;
        ELSIF x =- 16880 THEN
            sigmoid_f := 1;
        ELSIF x =- 16879 THEN
            sigmoid_f := 1;
        ELSIF x =- 16878 THEN
            sigmoid_f := 1;
        ELSIF x =- 16877 THEN
            sigmoid_f := 1;
        ELSIF x =- 16876 THEN
            sigmoid_f := 1;
        ELSIF x =- 16875 THEN
            sigmoid_f := 1;
        ELSIF x =- 16874 THEN
            sigmoid_f := 1;
        ELSIF x =- 16873 THEN
            sigmoid_f := 1;
        ELSIF x =- 16872 THEN
            sigmoid_f := 1;
        ELSIF x =- 16871 THEN
            sigmoid_f := 1;
        ELSIF x =- 16870 THEN
            sigmoid_f := 1;
        ELSIF x =- 16869 THEN
            sigmoid_f := 1;
        ELSIF x =- 16868 THEN
            sigmoid_f := 1;
        ELSIF x =- 16867 THEN
            sigmoid_f := 1;
        ELSIF x =- 16866 THEN
            sigmoid_f := 1;
        ELSIF x =- 16865 THEN
            sigmoid_f := 1;
        ELSIF x =- 16864 THEN
            sigmoid_f := 1;
        ELSIF x =- 16863 THEN
            sigmoid_f := 1;
        ELSIF x =- 16862 THEN
            sigmoid_f := 1;
        ELSIF x =- 16861 THEN
            sigmoid_f := 1;
        ELSIF x =- 16860 THEN
            sigmoid_f := 1;
        ELSIF x =- 16859 THEN
            sigmoid_f := 1;
        ELSIF x =- 16858 THEN
            sigmoid_f := 1;
        ELSIF x =- 16857 THEN
            sigmoid_f := 1;
        ELSIF x =- 16856 THEN
            sigmoid_f := 1;
        ELSIF x =- 16855 THEN
            sigmoid_f := 1;
        ELSIF x =- 16854 THEN
            sigmoid_f := 1;
        ELSIF x =- 16853 THEN
            sigmoid_f := 1;
        ELSIF x =- 16852 THEN
            sigmoid_f := 1;
        ELSIF x =- 16851 THEN
            sigmoid_f := 1;
        ELSIF x =- 16850 THEN
            sigmoid_f := 1;
        ELSIF x =- 16849 THEN
            sigmoid_f := 1;
        ELSIF x =- 16848 THEN
            sigmoid_f := 1;
        ELSIF x =- 16847 THEN
            sigmoid_f := 1;
        ELSIF x =- 16846 THEN
            sigmoid_f := 1;
        ELSIF x =- 16845 THEN
            sigmoid_f := 1;
        ELSIF x =- 16844 THEN
            sigmoid_f := 1;
        ELSIF x =- 16843 THEN
            sigmoid_f := 1;
        ELSIF x =- 16842 THEN
            sigmoid_f := 1;
        ELSIF x =- 16841 THEN
            sigmoid_f := 1;
        ELSIF x =- 16840 THEN
            sigmoid_f := 1;
        ELSIF x =- 16839 THEN
            sigmoid_f := 1;
        ELSIF x =- 16838 THEN
            sigmoid_f := 1;
        ELSIF x =- 16837 THEN
            sigmoid_f := 1;
        ELSIF x =- 16836 THEN
            sigmoid_f := 1;
        ELSIF x =- 16835 THEN
            sigmoid_f := 1;
        ELSIF x =- 16834 THEN
            sigmoid_f := 1;
        ELSIF x =- 16833 THEN
            sigmoid_f := 1;
        ELSIF x =- 16832 THEN
            sigmoid_f := 1;
        ELSIF x =- 16831 THEN
            sigmoid_f := 1;
        ELSIF x =- 16830 THEN
            sigmoid_f := 1;
        ELSIF x =- 16829 THEN
            sigmoid_f := 1;
        ELSIF x =- 16828 THEN
            sigmoid_f := 1;
        ELSIF x =- 16827 THEN
            sigmoid_f := 1;
        ELSIF x =- 16826 THEN
            sigmoid_f := 1;
        ELSIF x =- 16825 THEN
            sigmoid_f := 1;
        ELSIF x =- 16824 THEN
            sigmoid_f := 1;
        ELSIF x =- 16823 THEN
            sigmoid_f := 1;
        ELSIF x =- 16822 THEN
            sigmoid_f := 1;
        ELSIF x =- 16821 THEN
            sigmoid_f := 1;
        ELSIF x =- 16820 THEN
            sigmoid_f := 1;
        ELSIF x =- 16819 THEN
            sigmoid_f := 1;
        ELSIF x =- 16818 THEN
            sigmoid_f := 1;
        ELSIF x =- 16817 THEN
            sigmoid_f := 1;
        ELSIF x =- 16816 THEN
            sigmoid_f := 1;
        ELSIF x =- 16815 THEN
            sigmoid_f := 1;
        ELSIF x =- 16814 THEN
            sigmoid_f := 1;
        ELSIF x =- 16813 THEN
            sigmoid_f := 1;
        ELSIF x =- 16812 THEN
            sigmoid_f := 1;
        ELSIF x =- 16811 THEN
            sigmoid_f := 1;
        ELSIF x =- 16810 THEN
            sigmoid_f := 1;
        ELSIF x =- 16809 THEN
            sigmoid_f := 1;
        ELSIF x =- 16808 THEN
            sigmoid_f := 1;
        ELSIF x =- 16807 THEN
            sigmoid_f := 1;
        ELSIF x =- 16806 THEN
            sigmoid_f := 1;
        ELSIF x =- 16805 THEN
            sigmoid_f := 1;
        ELSIF x =- 16804 THEN
            sigmoid_f := 1;
        ELSIF x =- 16803 THEN
            sigmoid_f := 1;
        ELSIF x =- 16802 THEN
            sigmoid_f := 1;
        ELSIF x =- 16801 THEN
            sigmoid_f := 1;
        ELSIF x =- 16800 THEN
            sigmoid_f := 1;
        ELSIF x =- 16799 THEN
            sigmoid_f := 1;
        ELSIF x =- 16798 THEN
            sigmoid_f := 1;
        ELSIF x =- 16797 THEN
            sigmoid_f := 1;
        ELSIF x =- 16796 THEN
            sigmoid_f := 1;
        ELSIF x =- 16795 THEN
            sigmoid_f := 1;
        ELSIF x =- 16794 THEN
            sigmoid_f := 1;
        ELSIF x =- 16793 THEN
            sigmoid_f := 1;
        ELSIF x =- 16792 THEN
            sigmoid_f := 1;
        ELSIF x =- 16791 THEN
            sigmoid_f := 1;
        ELSIF x =- 16790 THEN
            sigmoid_f := 1;
        ELSIF x =- 16789 THEN
            sigmoid_f := 1;
        ELSIF x =- 16788 THEN
            sigmoid_f := 1;
        ELSIF x =- 16787 THEN
            sigmoid_f := 1;
        ELSIF x =- 16786 THEN
            sigmoid_f := 1;
        ELSIF x =- 16785 THEN
            sigmoid_f := 1;
        ELSIF x =- 16784 THEN
            sigmoid_f := 1;
        ELSIF x =- 16783 THEN
            sigmoid_f := 1;
        ELSIF x =- 16782 THEN
            sigmoid_f := 1;
        ELSIF x =- 16781 THEN
            sigmoid_f := 1;
        ELSIF x =- 16780 THEN
            sigmoid_f := 1;
        ELSIF x =- 16779 THEN
            sigmoid_f := 1;
        ELSIF x =- 16778 THEN
            sigmoid_f := 1;
        ELSIF x =- 16777 THEN
            sigmoid_f := 1;
        ELSIF x =- 16776 THEN
            sigmoid_f := 1;
        ELSIF x =- 16775 THEN
            sigmoid_f := 1;
        ELSIF x =- 16774 THEN
            sigmoid_f := 1;
        ELSIF x =- 16773 THEN
            sigmoid_f := 1;
        ELSIF x =- 16772 THEN
            sigmoid_f := 1;
        ELSIF x =- 16771 THEN
            sigmoid_f := 1;
        ELSIF x =- 16770 THEN
            sigmoid_f := 1;
        ELSIF x =- 16769 THEN
            sigmoid_f := 1;
        ELSIF x =- 16768 THEN
            sigmoid_f := 1;
        ELSIF x =- 16767 THEN
            sigmoid_f := 1;
        ELSIF x =- 16766 THEN
            sigmoid_f := 1;
        ELSIF x =- 16765 THEN
            sigmoid_f := 1;
        ELSIF x =- 16764 THEN
            sigmoid_f := 1;
        ELSIF x =- 16763 THEN
            sigmoid_f := 1;
        ELSIF x =- 16762 THEN
            sigmoid_f := 1;
        ELSIF x =- 16761 THEN
            sigmoid_f := 1;
        ELSIF x =- 16760 THEN
            sigmoid_f := 1;
        ELSIF x =- 16759 THEN
            sigmoid_f := 1;
        ELSIF x =- 16758 THEN
            sigmoid_f := 1;
        ELSIF x =- 16757 THEN
            sigmoid_f := 1;
        ELSIF x =- 16756 THEN
            sigmoid_f := 1;
        ELSIF x =- 16755 THEN
            sigmoid_f := 1;
        ELSIF x =- 16754 THEN
            sigmoid_f := 1;
        ELSIF x =- 16753 THEN
            sigmoid_f := 1;
        ELSIF x =- 16752 THEN
            sigmoid_f := 1;
        ELSIF x =- 16751 THEN
            sigmoid_f := 1;
        ELSIF x =- 16750 THEN
            sigmoid_f := 1;
        ELSIF x =- 16749 THEN
            sigmoid_f := 1;
        ELSIF x =- 16748 THEN
            sigmoid_f := 1;
        ELSIF x =- 16747 THEN
            sigmoid_f := 1;
        ELSIF x =- 16746 THEN
            sigmoid_f := 1;
        ELSIF x =- 16745 THEN
            sigmoid_f := 1;
        ELSIF x =- 16744 THEN
            sigmoid_f := 1;
        ELSIF x =- 16743 THEN
            sigmoid_f := 1;
        ELSIF x =- 16742 THEN
            sigmoid_f := 1;
        ELSIF x =- 16741 THEN
            sigmoid_f := 1;
        ELSIF x =- 16740 THEN
            sigmoid_f := 1;
        ELSIF x =- 16739 THEN
            sigmoid_f := 1;
        ELSIF x =- 16738 THEN
            sigmoid_f := 1;
        ELSIF x =- 16737 THEN
            sigmoid_f := 1;
        ELSIF x =- 16736 THEN
            sigmoid_f := 1;
        ELSIF x =- 16735 THEN
            sigmoid_f := 1;
        ELSIF x =- 16734 THEN
            sigmoid_f := 1;
        ELSIF x =- 16733 THEN
            sigmoid_f := 1;
        ELSIF x =- 16732 THEN
            sigmoid_f := 1;
        ELSIF x =- 16731 THEN
            sigmoid_f := 1;
        ELSIF x =- 16730 THEN
            sigmoid_f := 1;
        ELSIF x =- 16729 THEN
            sigmoid_f := 1;
        ELSIF x =- 16728 THEN
            sigmoid_f := 1;
        ELSIF x =- 16727 THEN
            sigmoid_f := 1;
        ELSIF x =- 16726 THEN
            sigmoid_f := 1;
        ELSIF x =- 16725 THEN
            sigmoid_f := 1;
        ELSIF x =- 16724 THEN
            sigmoid_f := 1;
        ELSIF x =- 16723 THEN
            sigmoid_f := 1;
        ELSIF x =- 16722 THEN
            sigmoid_f := 1;
        ELSIF x =- 16721 THEN
            sigmoid_f := 1;
        ELSIF x =- 16720 THEN
            sigmoid_f := 1;
        ELSIF x =- 16719 THEN
            sigmoid_f := 1;
        ELSIF x =- 16718 THEN
            sigmoid_f := 1;
        ELSIF x =- 16717 THEN
            sigmoid_f := 1;
        ELSIF x =- 16716 THEN
            sigmoid_f := 1;
        ELSIF x =- 16715 THEN
            sigmoid_f := 1;
        ELSIF x =- 16714 THEN
            sigmoid_f := 1;
        ELSIF x =- 16713 THEN
            sigmoid_f := 1;
        ELSIF x =- 16712 THEN
            sigmoid_f := 1;
        ELSIF x =- 16711 THEN
            sigmoid_f := 1;
        ELSIF x =- 16710 THEN
            sigmoid_f := 1;
        ELSIF x =- 16709 THEN
            sigmoid_f := 1;
        ELSIF x =- 16708 THEN
            sigmoid_f := 1;
        ELSIF x =- 16707 THEN
            sigmoid_f := 1;
        ELSIF x =- 16706 THEN
            sigmoid_f := 1;
        ELSIF x =- 16705 THEN
            sigmoid_f := 1;
        ELSIF x =- 16704 THEN
            sigmoid_f := 1;
        ELSIF x =- 16703 THEN
            sigmoid_f := 1;
        ELSIF x =- 16702 THEN
            sigmoid_f := 1;
        ELSIF x =- 16701 THEN
            sigmoid_f := 1;
        ELSIF x =- 16700 THEN
            sigmoid_f := 1;
        ELSIF x =- 16699 THEN
            sigmoid_f := 1;
        ELSIF x =- 16698 THEN
            sigmoid_f := 1;
        ELSIF x =- 16697 THEN
            sigmoid_f := 1;
        ELSIF x =- 16696 THEN
            sigmoid_f := 1;
        ELSIF x =- 16695 THEN
            sigmoid_f := 1;
        ELSIF x =- 16694 THEN
            sigmoid_f := 1;
        ELSIF x =- 16693 THEN
            sigmoid_f := 1;
        ELSIF x =- 16692 THEN
            sigmoid_f := 1;
        ELSIF x =- 16691 THEN
            sigmoid_f := 1;
        ELSIF x =- 16690 THEN
            sigmoid_f := 1;
        ELSIF x =- 16689 THEN
            sigmoid_f := 1;
        ELSIF x =- 16688 THEN
            sigmoid_f := 1;
        ELSIF x =- 16687 THEN
            sigmoid_f := 1;
        ELSIF x =- 16686 THEN
            sigmoid_f := 1;
        ELSIF x =- 16685 THEN
            sigmoid_f := 1;
        ELSIF x =- 16684 THEN
            sigmoid_f := 1;
        ELSIF x =- 16683 THEN
            sigmoid_f := 1;
        ELSIF x =- 16682 THEN
            sigmoid_f := 1;
        ELSIF x =- 16681 THEN
            sigmoid_f := 1;
        ELSIF x =- 16680 THEN
            sigmoid_f := 1;
        ELSIF x =- 16679 THEN
            sigmoid_f := 1;
        ELSIF x =- 16678 THEN
            sigmoid_f := 1;
        ELSIF x =- 16677 THEN
            sigmoid_f := 1;
        ELSIF x =- 16676 THEN
            sigmoid_f := 1;
        ELSIF x =- 16675 THEN
            sigmoid_f := 1;
        ELSIF x =- 16674 THEN
            sigmoid_f := 1;
        ELSIF x =- 16673 THEN
            sigmoid_f := 1;
        ELSIF x =- 16672 THEN
            sigmoid_f := 1;
        ELSIF x =- 16671 THEN
            sigmoid_f := 1;
        ELSIF x =- 16670 THEN
            sigmoid_f := 1;
        ELSIF x =- 16669 THEN
            sigmoid_f := 1;
        ELSIF x =- 16668 THEN
            sigmoid_f := 1;
        ELSIF x =- 16667 THEN
            sigmoid_f := 1;
        ELSIF x =- 16666 THEN
            sigmoid_f := 1;
        ELSIF x =- 16665 THEN
            sigmoid_f := 1;
        ELSIF x =- 16664 THEN
            sigmoid_f := 1;
        ELSIF x =- 16663 THEN
            sigmoid_f := 1;
        ELSIF x =- 16662 THEN
            sigmoid_f := 1;
        ELSIF x =- 16661 THEN
            sigmoid_f := 1;
        ELSIF x =- 16660 THEN
            sigmoid_f := 1;
        ELSIF x =- 16659 THEN
            sigmoid_f := 1;
        ELSIF x =- 16658 THEN
            sigmoid_f := 1;
        ELSIF x =- 16657 THEN
            sigmoid_f := 1;
        ELSIF x =- 16656 THEN
            sigmoid_f := 1;
        ELSIF x =- 16655 THEN
            sigmoid_f := 1;
        ELSIF x =- 16654 THEN
            sigmoid_f := 1;
        ELSIF x =- 16653 THEN
            sigmoid_f := 1;
        ELSIF x =- 16652 THEN
            sigmoid_f := 1;
        ELSIF x =- 16651 THEN
            sigmoid_f := 1;
        ELSIF x =- 16650 THEN
            sigmoid_f := 1;
        ELSIF x =- 16649 THEN
            sigmoid_f := 1;
        ELSIF x =- 16648 THEN
            sigmoid_f := 1;
        ELSIF x =- 16647 THEN
            sigmoid_f := 1;
        ELSIF x =- 16646 THEN
            sigmoid_f := 1;
        ELSIF x =- 16645 THEN
            sigmoid_f := 1;
        ELSIF x =- 16644 THEN
            sigmoid_f := 1;
        ELSIF x =- 16643 THEN
            sigmoid_f := 1;
        ELSIF x =- 16642 THEN
            sigmoid_f := 1;
        ELSIF x =- 16641 THEN
            sigmoid_f := 1;
        ELSIF x =- 16640 THEN
            sigmoid_f := 1;
        ELSIF x =- 16639 THEN
            sigmoid_f := 1;
        ELSIF x =- 16638 THEN
            sigmoid_f := 1;
        ELSIF x =- 16637 THEN
            sigmoid_f := 1;
        ELSIF x =- 16636 THEN
            sigmoid_f := 1;
        ELSIF x =- 16635 THEN
            sigmoid_f := 1;
        ELSIF x =- 16634 THEN
            sigmoid_f := 1;
        ELSIF x =- 16633 THEN
            sigmoid_f := 1;
        ELSIF x =- 16632 THEN
            sigmoid_f := 1;
        ELSIF x =- 16631 THEN
            sigmoid_f := 1;
        ELSIF x =- 16630 THEN
            sigmoid_f := 1;
        ELSIF x =- 16629 THEN
            sigmoid_f := 1;
        ELSIF x =- 16628 THEN
            sigmoid_f := 1;
        ELSIF x =- 16627 THEN
            sigmoid_f := 1;
        ELSIF x =- 16626 THEN
            sigmoid_f := 1;
        ELSIF x =- 16625 THEN
            sigmoid_f := 1;
        ELSIF x =- 16624 THEN
            sigmoid_f := 1;
        ELSIF x =- 16623 THEN
            sigmoid_f := 1;
        ELSIF x =- 16622 THEN
            sigmoid_f := 1;
        ELSIF x =- 16621 THEN
            sigmoid_f := 1;
        ELSIF x =- 16620 THEN
            sigmoid_f := 1;
        ELSIF x =- 16619 THEN
            sigmoid_f := 1;
        ELSIF x =- 16618 THEN
            sigmoid_f := 1;
        ELSIF x =- 16617 THEN
            sigmoid_f := 1;
        ELSIF x =- 16616 THEN
            sigmoid_f := 1;
        ELSIF x =- 16615 THEN
            sigmoid_f := 1;
        ELSIF x =- 16614 THEN
            sigmoid_f := 1;
        ELSIF x =- 16613 THEN
            sigmoid_f := 1;
        ELSIF x =- 16612 THEN
            sigmoid_f := 1;
        ELSIF x =- 16611 THEN
            sigmoid_f := 1;
        ELSIF x =- 16610 THEN
            sigmoid_f := 1;
        ELSIF x =- 16609 THEN
            sigmoid_f := 1;
        ELSIF x =- 16608 THEN
            sigmoid_f := 1;
        ELSIF x =- 16607 THEN
            sigmoid_f := 1;
        ELSIF x =- 16606 THEN
            sigmoid_f := 1;
        ELSIF x =- 16605 THEN
            sigmoid_f := 1;
        ELSIF x =- 16604 THEN
            sigmoid_f := 1;
        ELSIF x =- 16603 THEN
            sigmoid_f := 1;
        ELSIF x =- 16602 THEN
            sigmoid_f := 1;
        ELSIF x =- 16601 THEN
            sigmoid_f := 1;
        ELSIF x =- 16600 THEN
            sigmoid_f := 1;
        ELSIF x =- 16599 THEN
            sigmoid_f := 1;
        ELSIF x =- 16598 THEN
            sigmoid_f := 1;
        ELSIF x =- 16597 THEN
            sigmoid_f := 1;
        ELSIF x =- 16596 THEN
            sigmoid_f := 1;
        ELSIF x =- 16595 THEN
            sigmoid_f := 1;
        ELSIF x =- 16594 THEN
            sigmoid_f := 1;
        ELSIF x =- 16593 THEN
            sigmoid_f := 1;
        ELSIF x =- 16592 THEN
            sigmoid_f := 1;
        ELSIF x =- 16591 THEN
            sigmoid_f := 1;
        ELSIF x =- 16590 THEN
            sigmoid_f := 1;
        ELSIF x =- 16589 THEN
            sigmoid_f := 1;
        ELSIF x =- 16588 THEN
            sigmoid_f := 1;
        ELSIF x =- 16587 THEN
            sigmoid_f := 1;
        ELSIF x =- 16586 THEN
            sigmoid_f := 1;
        ELSIF x =- 16585 THEN
            sigmoid_f := 1;
        ELSIF x =- 16584 THEN
            sigmoid_f := 1;
        ELSIF x =- 16583 THEN
            sigmoid_f := 1;
        ELSIF x =- 16582 THEN
            sigmoid_f := 1;
        ELSIF x =- 16581 THEN
            sigmoid_f := 1;
        ELSIF x =- 16580 THEN
            sigmoid_f := 1;
        ELSIF x =- 16579 THEN
            sigmoid_f := 1;
        ELSIF x =- 16578 THEN
            sigmoid_f := 1;
        ELSIF x =- 16577 THEN
            sigmoid_f := 1;
        ELSIF x =- 16576 THEN
            sigmoid_f := 1;
        ELSIF x =- 16575 THEN
            sigmoid_f := 1;
        ELSIF x =- 16574 THEN
            sigmoid_f := 1;
        ELSIF x =- 16573 THEN
            sigmoid_f := 1;
        ELSIF x =- 16572 THEN
            sigmoid_f := 1;
        ELSIF x =- 16571 THEN
            sigmoid_f := 1;
        ELSIF x =- 16570 THEN
            sigmoid_f := 1;
        ELSIF x =- 16569 THEN
            sigmoid_f := 1;
        ELSIF x =- 16568 THEN
            sigmoid_f := 1;
        ELSIF x =- 16567 THEN
            sigmoid_f := 1;
        ELSIF x =- 16566 THEN
            sigmoid_f := 1;
        ELSIF x =- 16565 THEN
            sigmoid_f := 1;
        ELSIF x =- 16564 THEN
            sigmoid_f := 1;
        ELSIF x =- 16563 THEN
            sigmoid_f := 1;
        ELSIF x =- 16562 THEN
            sigmoid_f := 1;
        ELSIF x =- 16561 THEN
            sigmoid_f := 1;
        ELSIF x =- 16560 THEN
            sigmoid_f := 1;
        ELSIF x =- 16559 THEN
            sigmoid_f := 1;
        ELSIF x =- 16558 THEN
            sigmoid_f := 1;
        ELSIF x =- 16557 THEN
            sigmoid_f := 1;
        ELSIF x =- 16556 THEN
            sigmoid_f := 1;
        ELSIF x =- 16555 THEN
            sigmoid_f := 1;
        ELSIF x =- 16554 THEN
            sigmoid_f := 1;
        ELSIF x =- 16553 THEN
            sigmoid_f := 1;
        ELSIF x =- 16552 THEN
            sigmoid_f := 1;
        ELSIF x =- 16551 THEN
            sigmoid_f := 1;
        ELSIF x =- 16550 THEN
            sigmoid_f := 1;
        ELSIF x =- 16549 THEN
            sigmoid_f := 1;
        ELSIF x =- 16548 THEN
            sigmoid_f := 1;
        ELSIF x =- 16547 THEN
            sigmoid_f := 1;
        ELSIF x =- 16546 THEN
            sigmoid_f := 1;
        ELSIF x =- 16545 THEN
            sigmoid_f := 1;
        ELSIF x =- 16544 THEN
            sigmoid_f := 1;
        ELSIF x =- 16543 THEN
            sigmoid_f := 1;
        ELSIF x =- 16542 THEN
            sigmoid_f := 1;
        ELSIF x =- 16541 THEN
            sigmoid_f := 1;
        ELSIF x =- 16540 THEN
            sigmoid_f := 1;
        ELSIF x =- 16539 THEN
            sigmoid_f := 1;
        ELSIF x =- 16538 THEN
            sigmoid_f := 1;
        ELSIF x =- 16537 THEN
            sigmoid_f := 1;
        ELSIF x =- 16536 THEN
            sigmoid_f := 1;
        ELSIF x =- 16535 THEN
            sigmoid_f := 1;
        ELSIF x =- 16534 THEN
            sigmoid_f := 1;
        ELSIF x =- 16533 THEN
            sigmoid_f := 1;
        ELSIF x =- 16532 THEN
            sigmoid_f := 1;
        ELSIF x =- 16531 THEN
            sigmoid_f := 1;
        ELSIF x =- 16530 THEN
            sigmoid_f := 1;
        ELSIF x =- 16529 THEN
            sigmoid_f := 1;
        ELSIF x =- 16528 THEN
            sigmoid_f := 1;
        ELSIF x =- 16527 THEN
            sigmoid_f := 1;
        ELSIF x =- 16526 THEN
            sigmoid_f := 1;
        ELSIF x =- 16525 THEN
            sigmoid_f := 1;
        ELSIF x =- 16524 THEN
            sigmoid_f := 1;
        ELSIF x =- 16523 THEN
            sigmoid_f := 1;
        ELSIF x =- 16522 THEN
            sigmoid_f := 1;
        ELSIF x =- 16521 THEN
            sigmoid_f := 1;
        ELSIF x =- 16520 THEN
            sigmoid_f := 1;
        ELSIF x =- 16519 THEN
            sigmoid_f := 1;
        ELSIF x =- 16518 THEN
            sigmoid_f := 1;
        ELSIF x =- 16517 THEN
            sigmoid_f := 1;
        ELSIF x =- 16516 THEN
            sigmoid_f := 1;
        ELSIF x =- 16515 THEN
            sigmoid_f := 1;
        ELSIF x =- 16514 THEN
            sigmoid_f := 1;
        ELSIF x =- 16513 THEN
            sigmoid_f := 1;
        ELSIF x =- 16512 THEN
            sigmoid_f := 1;
        ELSIF x =- 16511 THEN
            sigmoid_f := 1;
        ELSIF x =- 16510 THEN
            sigmoid_f := 1;
        ELSIF x =- 16509 THEN
            sigmoid_f := 1;
        ELSIF x =- 16508 THEN
            sigmoid_f := 1;
        ELSIF x =- 16507 THEN
            sigmoid_f := 1;
        ELSIF x =- 16506 THEN
            sigmoid_f := 1;
        ELSIF x =- 16505 THEN
            sigmoid_f := 1;
        ELSIF x =- 16504 THEN
            sigmoid_f := 1;
        ELSIF x =- 16503 THEN
            sigmoid_f := 1;
        ELSIF x =- 16502 THEN
            sigmoid_f := 1;
        ELSIF x =- 16501 THEN
            sigmoid_f := 1;
        ELSIF x =- 16500 THEN
            sigmoid_f := 1;
        ELSIF x =- 16499 THEN
            sigmoid_f := 1;
        ELSIF x =- 16498 THEN
            sigmoid_f := 1;
        ELSIF x =- 16497 THEN
            sigmoid_f := 1;
        ELSIF x =- 16496 THEN
            sigmoid_f := 1;
        ELSIF x =- 16495 THEN
            sigmoid_f := 1;
        ELSIF x =- 16494 THEN
            sigmoid_f := 1;
        ELSIF x =- 16493 THEN
            sigmoid_f := 1;
        ELSIF x =- 16492 THEN
            sigmoid_f := 1;
        ELSIF x =- 16491 THEN
            sigmoid_f := 1;
        ELSIF x =- 16490 THEN
            sigmoid_f := 1;
        ELSIF x =- 16489 THEN
            sigmoid_f := 1;
        ELSIF x =- 16488 THEN
            sigmoid_f := 1;
        ELSIF x =- 16487 THEN
            sigmoid_f := 1;
        ELSIF x =- 16486 THEN
            sigmoid_f := 1;
        ELSIF x =- 16485 THEN
            sigmoid_f := 1;
        ELSIF x =- 16484 THEN
            sigmoid_f := 1;
        ELSIF x =- 16483 THEN
            sigmoid_f := 1;
        ELSIF x =- 16482 THEN
            sigmoid_f := 1;
        ELSIF x =- 16481 THEN
            sigmoid_f := 1;
        ELSIF x =- 16480 THEN
            sigmoid_f := 1;
        ELSIF x =- 16479 THEN
            sigmoid_f := 1;
        ELSIF x =- 16478 THEN
            sigmoid_f := 1;
        ELSIF x =- 16477 THEN
            sigmoid_f := 1;
        ELSIF x =- 16476 THEN
            sigmoid_f := 1;
        ELSIF x =- 16475 THEN
            sigmoid_f := 1;
        ELSIF x =- 16474 THEN
            sigmoid_f := 1;
        ELSIF x =- 16473 THEN
            sigmoid_f := 1;
        ELSIF x =- 16472 THEN
            sigmoid_f := 1;
        ELSIF x =- 16471 THEN
            sigmoid_f := 1;
        ELSIF x =- 16470 THEN
            sigmoid_f := 1;
        ELSIF x =- 16469 THEN
            sigmoid_f := 1;
        ELSIF x =- 16468 THEN
            sigmoid_f := 1;
        ELSIF x =- 16467 THEN
            sigmoid_f := 1;
        ELSIF x =- 16466 THEN
            sigmoid_f := 1;
        ELSIF x =- 16465 THEN
            sigmoid_f := 1;
        ELSIF x =- 16464 THEN
            sigmoid_f := 1;
        ELSIF x =- 16463 THEN
            sigmoid_f := 1;
        ELSIF x =- 16462 THEN
            sigmoid_f := 1;
        ELSIF x =- 16461 THEN
            sigmoid_f := 1;
        ELSIF x =- 16460 THEN
            sigmoid_f := 1;
        ELSIF x =- 16459 THEN
            sigmoid_f := 1;
        ELSIF x =- 16458 THEN
            sigmoid_f := 1;
        ELSIF x =- 16457 THEN
            sigmoid_f := 1;
        ELSIF x =- 16456 THEN
            sigmoid_f := 1;
        ELSIF x =- 16455 THEN
            sigmoid_f := 1;
        ELSIF x =- 16454 THEN
            sigmoid_f := 1;
        ELSIF x =- 16453 THEN
            sigmoid_f := 1;
        ELSIF x =- 16452 THEN
            sigmoid_f := 1;
        ELSIF x =- 16451 THEN
            sigmoid_f := 1;
        ELSIF x =- 16450 THEN
            sigmoid_f := 1;
        ELSIF x =- 16449 THEN
            sigmoid_f := 1;
        ELSIF x =- 16448 THEN
            sigmoid_f := 1;
        ELSIF x =- 16447 THEN
            sigmoid_f := 1;
        ELSIF x =- 16446 THEN
            sigmoid_f := 1;
        ELSIF x =- 16445 THEN
            sigmoid_f := 1;
        ELSIF x =- 16444 THEN
            sigmoid_f := 1;
        ELSIF x =- 16443 THEN
            sigmoid_f := 1;
        ELSIF x =- 16442 THEN
            sigmoid_f := 1;
        ELSIF x =- 16441 THEN
            sigmoid_f := 1;
        ELSIF x =- 16440 THEN
            sigmoid_f := 1;
        ELSIF x =- 16439 THEN
            sigmoid_f := 1;
        ELSIF x =- 16438 THEN
            sigmoid_f := 1;
        ELSIF x =- 16437 THEN
            sigmoid_f := 1;
        ELSIF x =- 16436 THEN
            sigmoid_f := 1;
        ELSIF x =- 16435 THEN
            sigmoid_f := 1;
        ELSIF x =- 16434 THEN
            sigmoid_f := 1;
        ELSIF x =- 16433 THEN
            sigmoid_f := 1;
        ELSIF x =- 16432 THEN
            sigmoid_f := 1;
        ELSIF x =- 16431 THEN
            sigmoid_f := 1;
        ELSIF x =- 16430 THEN
            sigmoid_f := 1;
        ELSIF x =- 16429 THEN
            sigmoid_f := 1;
        ELSIF x =- 16428 THEN
            sigmoid_f := 1;
        ELSIF x =- 16427 THEN
            sigmoid_f := 1;
        ELSIF x =- 16426 THEN
            sigmoid_f := 1;
        ELSIF x =- 16425 THEN
            sigmoid_f := 1;
        ELSIF x =- 16424 THEN
            sigmoid_f := 1;
        ELSIF x =- 16423 THEN
            sigmoid_f := 1;
        ELSIF x =- 16422 THEN
            sigmoid_f := 1;
        ELSIF x =- 16421 THEN
            sigmoid_f := 1;
        ELSIF x =- 16420 THEN
            sigmoid_f := 1;
        ELSIF x =- 16419 THEN
            sigmoid_f := 1;
        ELSIF x =- 16418 THEN
            sigmoid_f := 1;
        ELSIF x =- 16417 THEN
            sigmoid_f := 1;
        ELSIF x =- 16416 THEN
            sigmoid_f := 1;
        ELSIF x =- 16415 THEN
            sigmoid_f := 1;
        ELSIF x =- 16414 THEN
            sigmoid_f := 1;
        ELSIF x =- 16413 THEN
            sigmoid_f := 1;
        ELSIF x =- 16412 THEN
            sigmoid_f := 1;
        ELSIF x =- 16411 THEN
            sigmoid_f := 1;
        ELSIF x =- 16410 THEN
            sigmoid_f := 1;
        ELSIF x =- 16409 THEN
            sigmoid_f := 1;
        ELSIF x =- 16408 THEN
            sigmoid_f := 1;
        ELSIF x =- 16407 THEN
            sigmoid_f := 1;
        ELSIF x =- 16406 THEN
            sigmoid_f := 1;
        ELSIF x =- 16405 THEN
            sigmoid_f := 1;
        ELSIF x =- 16404 THEN
            sigmoid_f := 1;
        ELSIF x =- 16403 THEN
            sigmoid_f := 1;
        ELSIF x =- 16402 THEN
            sigmoid_f := 1;
        ELSIF x =- 16401 THEN
            sigmoid_f := 1;
        ELSIF x =- 16400 THEN
            sigmoid_f := 1;
        ELSIF x =- 16399 THEN
            sigmoid_f := 1;
        ELSIF x =- 16398 THEN
            sigmoid_f := 1;
        ELSIF x =- 16397 THEN
            sigmoid_f := 1;
        ELSIF x =- 16396 THEN
            sigmoid_f := 1;
        ELSIF x =- 16395 THEN
            sigmoid_f := 1;
        ELSIF x =- 16394 THEN
            sigmoid_f := 1;
        ELSIF x =- 16393 THEN
            sigmoid_f := 1;
        ELSIF x =- 16392 THEN
            sigmoid_f := 1;
        ELSIF x =- 16391 THEN
            sigmoid_f := 1;
        ELSIF x =- 16390 THEN
            sigmoid_f := 1;
        ELSIF x =- 16389 THEN
            sigmoid_f := 1;
        ELSIF x =- 16388 THEN
            sigmoid_f := 1;
        ELSIF x =- 16387 THEN
            sigmoid_f := 1;
        ELSIF x =- 16386 THEN
            sigmoid_f := 1;
        ELSIF x =- 16385 THEN
            sigmoid_f := 1;
        ELSIF x =- 16384 THEN
            sigmoid_f := 1;
        ELSIF x =- 16383 THEN
            sigmoid_f := 1;
        ELSIF x =- 16382 THEN
            sigmoid_f := 1;
        ELSIF x =- 16381 THEN
            sigmoid_f := 1;
        ELSIF x =- 16380 THEN
            sigmoid_f := 1;
        ELSIF x =- 16379 THEN
            sigmoid_f := 1;
        ELSIF x =- 16378 THEN
            sigmoid_f := 1;
        ELSIF x =- 16377 THEN
            sigmoid_f := 1;
        ELSIF x =- 16376 THEN
            sigmoid_f := 1;
        ELSIF x =- 16375 THEN
            sigmoid_f := 1;
        ELSIF x =- 16374 THEN
            sigmoid_f := 1;
        ELSIF x =- 16373 THEN
            sigmoid_f := 1;
        ELSIF x =- 16372 THEN
            sigmoid_f := 1;
        ELSIF x =- 16371 THEN
            sigmoid_f := 1;
        ELSIF x =- 16370 THEN
            sigmoid_f := 1;
        ELSIF x =- 16369 THEN
            sigmoid_f := 1;
        ELSIF x =- 16368 THEN
            sigmoid_f := 1;
        ELSIF x =- 16367 THEN
            sigmoid_f := 1;
        ELSIF x =- 16366 THEN
            sigmoid_f := 1;
        ELSIF x =- 16365 THEN
            sigmoid_f := 1;
        ELSIF x =- 16364 THEN
            sigmoid_f := 1;
        ELSIF x =- 16363 THEN
            sigmoid_f := 1;
        ELSIF x =- 16362 THEN
            sigmoid_f := 1;
        ELSIF x =- 16361 THEN
            sigmoid_f := 1;
        ELSIF x =- 16360 THEN
            sigmoid_f := 1;
        ELSIF x =- 16359 THEN
            sigmoid_f := 1;
        ELSIF x =- 16358 THEN
            sigmoid_f := 1;
        ELSIF x =- 16357 THEN
            sigmoid_f := 1;
        ELSIF x =- 16356 THEN
            sigmoid_f := 1;
        ELSIF x =- 16355 THEN
            sigmoid_f := 1;
        ELSIF x =- 16354 THEN
            sigmoid_f := 1;
        ELSIF x =- 16353 THEN
            sigmoid_f := 1;
        ELSIF x =- 16352 THEN
            sigmoid_f := 1;
        ELSIF x =- 16351 THEN
            sigmoid_f := 1;
        ELSIF x =- 16350 THEN
            sigmoid_f := 1;
        ELSIF x =- 16349 THEN
            sigmoid_f := 1;
        ELSIF x =- 16348 THEN
            sigmoid_f := 1;
        ELSIF x =- 16347 THEN
            sigmoid_f := 1;
        ELSIF x =- 16346 THEN
            sigmoid_f := 1;
        ELSIF x =- 16345 THEN
            sigmoid_f := 1;
        ELSIF x =- 16344 THEN
            sigmoid_f := 1;
        ELSIF x =- 16343 THEN
            sigmoid_f := 1;
        ELSIF x =- 16342 THEN
            sigmoid_f := 1;
        ELSIF x =- 16341 THEN
            sigmoid_f := 1;
        ELSIF x =- 16340 THEN
            sigmoid_f := 1;
        ELSIF x =- 16339 THEN
            sigmoid_f := 1;
        ELSIF x =- 16338 THEN
            sigmoid_f := 1;
        ELSIF x =- 16337 THEN
            sigmoid_f := 1;
        ELSIF x =- 16336 THEN
            sigmoid_f := 1;
        ELSIF x =- 16335 THEN
            sigmoid_f := 1;
        ELSIF x =- 16334 THEN
            sigmoid_f := 1;
        ELSIF x =- 16333 THEN
            sigmoid_f := 1;
        ELSIF x =- 16332 THEN
            sigmoid_f := 1;
        ELSIF x =- 16331 THEN
            sigmoid_f := 1;
        ELSIF x =- 16330 THEN
            sigmoid_f := 1;
        ELSIF x =- 16329 THEN
            sigmoid_f := 1;
        ELSIF x =- 16328 THEN
            sigmoid_f := 1;
        ELSIF x =- 16327 THEN
            sigmoid_f := 1;
        ELSIF x =- 16326 THEN
            sigmoid_f := 1;
        ELSIF x =- 16325 THEN
            sigmoid_f := 1;
        ELSIF x =- 16324 THEN
            sigmoid_f := 1;
        ELSIF x =- 16323 THEN
            sigmoid_f := 1;
        ELSIF x =- 16322 THEN
            sigmoid_f := 1;
        ELSIF x =- 16321 THEN
            sigmoid_f := 1;
        ELSIF x =- 16320 THEN
            sigmoid_f := 1;
        ELSIF x =- 16319 THEN
            sigmoid_f := 1;
        ELSIF x =- 16318 THEN
            sigmoid_f := 1;
        ELSIF x =- 16317 THEN
            sigmoid_f := 1;
        ELSIF x =- 16316 THEN
            sigmoid_f := 1;
        ELSIF x =- 16315 THEN
            sigmoid_f := 1;
        ELSIF x =- 16314 THEN
            sigmoid_f := 1;
        ELSIF x =- 16313 THEN
            sigmoid_f := 1;
        ELSIF x =- 16312 THEN
            sigmoid_f := 1;
        ELSIF x =- 16311 THEN
            sigmoid_f := 1;
        ELSIF x =- 16310 THEN
            sigmoid_f := 1;
        ELSIF x =- 16309 THEN
            sigmoid_f := 1;
        ELSIF x =- 16308 THEN
            sigmoid_f := 1;
        ELSIF x =- 16307 THEN
            sigmoid_f := 1;
        ELSIF x =- 16306 THEN
            sigmoid_f := 1;
        ELSIF x =- 16305 THEN
            sigmoid_f := 1;
        ELSIF x =- 16304 THEN
            sigmoid_f := 1;
        ELSIF x =- 16303 THEN
            sigmoid_f := 1;
        ELSIF x =- 16302 THEN
            sigmoid_f := 1;
        ELSIF x =- 16301 THEN
            sigmoid_f := 1;
        ELSIF x =- 16300 THEN
            sigmoid_f := 1;
        ELSIF x =- 16299 THEN
            sigmoid_f := 1;
        ELSIF x =- 16298 THEN
            sigmoid_f := 1;
        ELSIF x =- 16297 THEN
            sigmoid_f := 1;
        ELSIF x =- 16296 THEN
            sigmoid_f := 1;
        ELSIF x =- 16295 THEN
            sigmoid_f := 1;
        ELSIF x =- 16294 THEN
            sigmoid_f := 1;
        ELSIF x =- 16293 THEN
            sigmoid_f := 1;
        ELSIF x =- 16292 THEN
            sigmoid_f := 1;
        ELSIF x =- 16291 THEN
            sigmoid_f := 1;
        ELSIF x =- 16290 THEN
            sigmoid_f := 1;
        ELSIF x =- 16289 THEN
            sigmoid_f := 1;
        ELSIF x =- 16288 THEN
            sigmoid_f := 1;
        ELSIF x =- 16287 THEN
            sigmoid_f := 1;
        ELSIF x =- 16286 THEN
            sigmoid_f := 1;
        ELSIF x =- 16285 THEN
            sigmoid_f := 1;
        ELSIF x =- 16284 THEN
            sigmoid_f := 1;
        ELSIF x =- 16283 THEN
            sigmoid_f := 1;
        ELSIF x =- 16282 THEN
            sigmoid_f := 1;
        ELSIF x =- 16281 THEN
            sigmoid_f := 1;
        ELSIF x =- 16280 THEN
            sigmoid_f := 1;
        ELSIF x =- 16279 THEN
            sigmoid_f := 1;
        ELSIF x =- 16278 THEN
            sigmoid_f := 1;
        ELSIF x =- 16277 THEN
            sigmoid_f := 1;
        ELSIF x =- 16276 THEN
            sigmoid_f := 1;
        ELSIF x =- 16275 THEN
            sigmoid_f := 1;
        ELSIF x =- 16274 THEN
            sigmoid_f := 1;
        ELSIF x =- 16273 THEN
            sigmoid_f := 1;
        ELSIF x =- 16272 THEN
            sigmoid_f := 1;
        ELSIF x =- 16271 THEN
            sigmoid_f := 1;
        ELSIF x =- 16270 THEN
            sigmoid_f := 1;
        ELSIF x =- 16269 THEN
            sigmoid_f := 1;
        ELSIF x =- 16268 THEN
            sigmoid_f := 1;
        ELSIF x =- 16267 THEN
            sigmoid_f := 1;
        ELSIF x =- 16266 THEN
            sigmoid_f := 1;
        ELSIF x =- 16265 THEN
            sigmoid_f := 1;
        ELSIF x =- 16264 THEN
            sigmoid_f := 1;
        ELSIF x =- 16263 THEN
            sigmoid_f := 1;
        ELSIF x =- 16262 THEN
            sigmoid_f := 1;
        ELSIF x =- 16261 THEN
            sigmoid_f := 1;
        ELSIF x =- 16260 THEN
            sigmoid_f := 1;
        ELSIF x =- 16259 THEN
            sigmoid_f := 1;
        ELSIF x =- 16258 THEN
            sigmoid_f := 1;
        ELSIF x =- 16257 THEN
            sigmoid_f := 1;
        ELSIF x =- 16256 THEN
            sigmoid_f := 1;
        ELSIF x =- 16255 THEN
            sigmoid_f := 1;
        ELSIF x =- 16254 THEN
            sigmoid_f := 1;
        ELSIF x =- 16253 THEN
            sigmoid_f := 1;
        ELSIF x =- 16252 THEN
            sigmoid_f := 1;
        ELSIF x =- 16251 THEN
            sigmoid_f := 1;
        ELSIF x =- 16250 THEN
            sigmoid_f := 1;
        ELSIF x =- 16249 THEN
            sigmoid_f := 1;
        ELSIF x =- 16248 THEN
            sigmoid_f := 1;
        ELSIF x =- 16247 THEN
            sigmoid_f := 1;
        ELSIF x =- 16246 THEN
            sigmoid_f := 1;
        ELSIF x =- 16245 THEN
            sigmoid_f := 1;
        ELSIF x =- 16244 THEN
            sigmoid_f := 1;
        ELSIF x =- 16243 THEN
            sigmoid_f := 1;
        ELSIF x =- 16242 THEN
            sigmoid_f := 1;
        ELSIF x =- 16241 THEN
            sigmoid_f := 1;
        ELSIF x =- 16240 THEN
            sigmoid_f := 1;
        ELSIF x =- 16239 THEN
            sigmoid_f := 1;
        ELSIF x =- 16238 THEN
            sigmoid_f := 1;
        ELSIF x =- 16237 THEN
            sigmoid_f := 1;
        ELSIF x =- 16236 THEN
            sigmoid_f := 1;
        ELSIF x =- 16235 THEN
            sigmoid_f := 1;
        ELSIF x =- 16234 THEN
            sigmoid_f := 1;
        ELSIF x =- 16233 THEN
            sigmoid_f := 1;
        ELSIF x =- 16232 THEN
            sigmoid_f := 1;
        ELSIF x =- 16231 THEN
            sigmoid_f := 1;
        ELSIF x =- 16230 THEN
            sigmoid_f := 1;
        ELSIF x =- 16229 THEN
            sigmoid_f := 1;
        ELSIF x =- 16228 THEN
            sigmoid_f := 1;
        ELSIF x =- 16227 THEN
            sigmoid_f := 1;
        ELSIF x =- 16226 THEN
            sigmoid_f := 1;
        ELSIF x =- 16225 THEN
            sigmoid_f := 1;
        ELSIF x =- 16224 THEN
            sigmoid_f := 1;
        ELSIF x =- 16223 THEN
            sigmoid_f := 1;
        ELSIF x =- 16222 THEN
            sigmoid_f := 1;
        ELSIF x =- 16221 THEN
            sigmoid_f := 1;
        ELSIF x =- 16220 THEN
            sigmoid_f := 1;
        ELSIF x =- 16219 THEN
            sigmoid_f := 1;
        ELSIF x =- 16218 THEN
            sigmoid_f := 1;
        ELSIF x =- 16217 THEN
            sigmoid_f := 1;
        ELSIF x =- 16216 THEN
            sigmoid_f := 1;
        ELSIF x =- 16215 THEN
            sigmoid_f := 1;
        ELSIF x =- 16214 THEN
            sigmoid_f := 1;
        ELSIF x =- 16213 THEN
            sigmoid_f := 1;
        ELSIF x =- 16212 THEN
            sigmoid_f := 1;
        ELSIF x =- 16211 THEN
            sigmoid_f := 1;
        ELSIF x =- 16210 THEN
            sigmoid_f := 1;
        ELSIF x =- 16209 THEN
            sigmoid_f := 1;
        ELSIF x =- 16208 THEN
            sigmoid_f := 1;
        ELSIF x =- 16207 THEN
            sigmoid_f := 1;
        ELSIF x =- 16206 THEN
            sigmoid_f := 1;
        ELSIF x =- 16205 THEN
            sigmoid_f := 1;
        ELSIF x =- 16204 THEN
            sigmoid_f := 1;
        ELSIF x =- 16203 THEN
            sigmoid_f := 1;
        ELSIF x =- 16202 THEN
            sigmoid_f := 1;
        ELSIF x =- 16201 THEN
            sigmoid_f := 1;
        ELSIF x =- 16200 THEN
            sigmoid_f := 1;
        ELSIF x =- 16199 THEN
            sigmoid_f := 1;
        ELSIF x =- 16198 THEN
            sigmoid_f := 1;
        ELSIF x =- 16197 THEN
            sigmoid_f := 1;
        ELSIF x =- 16196 THEN
            sigmoid_f := 1;
        ELSIF x =- 16195 THEN
            sigmoid_f := 1;
        ELSIF x =- 16194 THEN
            sigmoid_f := 1;
        ELSIF x =- 16193 THEN
            sigmoid_f := 1;
        ELSIF x =- 16192 THEN
            sigmoid_f := 1;
        ELSIF x =- 16191 THEN
            sigmoid_f := 1;
        ELSIF x =- 16190 THEN
            sigmoid_f := 1;
        ELSIF x =- 16189 THEN
            sigmoid_f := 1;
        ELSIF x =- 16188 THEN
            sigmoid_f := 1;
        ELSIF x =- 16187 THEN
            sigmoid_f := 1;
        ELSIF x =- 16186 THEN
            sigmoid_f := 1;
        ELSIF x =- 16185 THEN
            sigmoid_f := 1;
        ELSIF x =- 16184 THEN
            sigmoid_f := 1;
        ELSIF x =- 16183 THEN
            sigmoid_f := 1;
        ELSIF x =- 16182 THEN
            sigmoid_f := 1;
        ELSIF x =- 16181 THEN
            sigmoid_f := 1;
        ELSIF x =- 16180 THEN
            sigmoid_f := 1;
        ELSIF x =- 16179 THEN
            sigmoid_f := 1;
        ELSIF x =- 16178 THEN
            sigmoid_f := 1;
        ELSIF x =- 16177 THEN
            sigmoid_f := 1;
        ELSIF x =- 16176 THEN
            sigmoid_f := 1;
        ELSIF x =- 16175 THEN
            sigmoid_f := 1;
        ELSIF x =- 16174 THEN
            sigmoid_f := 1;
        ELSIF x =- 16173 THEN
            sigmoid_f := 1;
        ELSIF x =- 16172 THEN
            sigmoid_f := 1;
        ELSIF x =- 16171 THEN
            sigmoid_f := 1;
        ELSIF x =- 16170 THEN
            sigmoid_f := 1;
        ELSIF x =- 16169 THEN
            sigmoid_f := 1;
        ELSIF x =- 16168 THEN
            sigmoid_f := 1;
        ELSIF x =- 16167 THEN
            sigmoid_f := 1;
        ELSIF x =- 16166 THEN
            sigmoid_f := 1;
        ELSIF x =- 16165 THEN
            sigmoid_f := 1;
        ELSIF x =- 16164 THEN
            sigmoid_f := 1;
        ELSIF x =- 16163 THEN
            sigmoid_f := 1;
        ELSIF x =- 16162 THEN
            sigmoid_f := 1;
        ELSIF x =- 16161 THEN
            sigmoid_f := 1;
        ELSIF x =- 16160 THEN
            sigmoid_f := 1;
        ELSIF x =- 16159 THEN
            sigmoid_f := 1;
        ELSIF x =- 16158 THEN
            sigmoid_f := 1;
        ELSIF x =- 16157 THEN
            sigmoid_f := 1;
        ELSIF x =- 16156 THEN
            sigmoid_f := 1;
        ELSIF x =- 16155 THEN
            sigmoid_f := 1;
        ELSIF x =- 16154 THEN
            sigmoid_f := 1;
        ELSIF x =- 16153 THEN
            sigmoid_f := 1;
        ELSIF x =- 16152 THEN
            sigmoid_f := 1;
        ELSIF x =- 16151 THEN
            sigmoid_f := 1;
        ELSIF x =- 16150 THEN
            sigmoid_f := 1;
        ELSIF x =- 16149 THEN
            sigmoid_f := 1;
        ELSIF x =- 16148 THEN
            sigmoid_f := 1;
        ELSIF x =- 16147 THEN
            sigmoid_f := 1;
        ELSIF x =- 16146 THEN
            sigmoid_f := 1;
        ELSIF x =- 16145 THEN
            sigmoid_f := 1;
        ELSIF x =- 16144 THEN
            sigmoid_f := 1;
        ELSIF x =- 16143 THEN
            sigmoid_f := 1;
        ELSIF x =- 16142 THEN
            sigmoid_f := 1;
        ELSIF x =- 16141 THEN
            sigmoid_f := 1;
        ELSIF x =- 16140 THEN
            sigmoid_f := 1;
        ELSIF x =- 16139 THEN
            sigmoid_f := 1;
        ELSIF x =- 16138 THEN
            sigmoid_f := 1;
        ELSIF x =- 16137 THEN
            sigmoid_f := 1;
        ELSIF x =- 16136 THEN
            sigmoid_f := 1;
        ELSIF x =- 16135 THEN
            sigmoid_f := 1;
        ELSIF x =- 16134 THEN
            sigmoid_f := 1;
        ELSIF x =- 16133 THEN
            sigmoid_f := 1;
        ELSIF x =- 16132 THEN
            sigmoid_f := 1;
        ELSIF x =- 16131 THEN
            sigmoid_f := 1;
        ELSIF x =- 16130 THEN
            sigmoid_f := 1;
        ELSIF x =- 16129 THEN
            sigmoid_f := 1;
        ELSIF x =- 16128 THEN
            sigmoid_f := 1;
        ELSIF x =- 16127 THEN
            sigmoid_f := 1;
        ELSIF x =- 16126 THEN
            sigmoid_f := 1;
        ELSIF x =- 16125 THEN
            sigmoid_f := 1;
        ELSIF x =- 16124 THEN
            sigmoid_f := 1;
        ELSIF x =- 16123 THEN
            sigmoid_f := 1;
        ELSIF x =- 16122 THEN
            sigmoid_f := 1;
        ELSIF x =- 16121 THEN
            sigmoid_f := 1;
        ELSIF x =- 16120 THEN
            sigmoid_f := 1;
        ELSIF x =- 16119 THEN
            sigmoid_f := 1;
        ELSIF x =- 16118 THEN
            sigmoid_f := 1;
        ELSIF x =- 16117 THEN
            sigmoid_f := 1;
        ELSIF x =- 16116 THEN
            sigmoid_f := 1;
        ELSIF x =- 16115 THEN
            sigmoid_f := 1;
        ELSIF x =- 16114 THEN
            sigmoid_f := 1;
        ELSIF x =- 16113 THEN
            sigmoid_f := 1;
        ELSIF x =- 16112 THEN
            sigmoid_f := 1;
        ELSIF x =- 16111 THEN
            sigmoid_f := 1;
        ELSIF x =- 16110 THEN
            sigmoid_f := 1;
        ELSIF x =- 16109 THEN
            sigmoid_f := 1;
        ELSIF x =- 16108 THEN
            sigmoid_f := 1;
        ELSIF x =- 16107 THEN
            sigmoid_f := 1;
        ELSIF x =- 16106 THEN
            sigmoid_f := 1;
        ELSIF x =- 16105 THEN
            sigmoid_f := 1;
        ELSIF x =- 16104 THEN
            sigmoid_f := 1;
        ELSIF x =- 16103 THEN
            sigmoid_f := 1;
        ELSIF x =- 16102 THEN
            sigmoid_f := 1;
        ELSIF x =- 16101 THEN
            sigmoid_f := 1;
        ELSIF x =- 16100 THEN
            sigmoid_f := 1;
        ELSIF x =- 16099 THEN
            sigmoid_f := 1;
        ELSIF x =- 16098 THEN
            sigmoid_f := 1;
        ELSIF x =- 16097 THEN
            sigmoid_f := 1;
        ELSIF x =- 16096 THEN
            sigmoid_f := 1;
        ELSIF x =- 16095 THEN
            sigmoid_f := 1;
        ELSIF x =- 16094 THEN
            sigmoid_f := 1;
        ELSIF x =- 16093 THEN
            sigmoid_f := 1;
        ELSIF x =- 16092 THEN
            sigmoid_f := 1;
        ELSIF x =- 16091 THEN
            sigmoid_f := 1;
        ELSIF x =- 16090 THEN
            sigmoid_f := 1;
        ELSIF x =- 16089 THEN
            sigmoid_f := 1;
        ELSIF x =- 16088 THEN
            sigmoid_f := 1;
        ELSIF x =- 16087 THEN
            sigmoid_f := 1;
        ELSIF x =- 16086 THEN
            sigmoid_f := 1;
        ELSIF x =- 16085 THEN
            sigmoid_f := 1;
        ELSIF x =- 16084 THEN
            sigmoid_f := 1;
        ELSIF x =- 16083 THEN
            sigmoid_f := 1;
        ELSIF x =- 16082 THEN
            sigmoid_f := 1;
        ELSIF x =- 16081 THEN
            sigmoid_f := 1;
        ELSIF x =- 16080 THEN
            sigmoid_f := 1;
        ELSIF x =- 16079 THEN
            sigmoid_f := 1;
        ELSIF x =- 16078 THEN
            sigmoid_f := 1;
        ELSIF x =- 16077 THEN
            sigmoid_f := 1;
        ELSIF x =- 16076 THEN
            sigmoid_f := 1;
        ELSIF x =- 16075 THEN
            sigmoid_f := 1;
        ELSIF x =- 16074 THEN
            sigmoid_f := 1;
        ELSIF x =- 16073 THEN
            sigmoid_f := 1;
        ELSIF x =- 16072 THEN
            sigmoid_f := 1;
        ELSIF x =- 16071 THEN
            sigmoid_f := 1;
        ELSIF x =- 16070 THEN
            sigmoid_f := 1;
        ELSIF x =- 16069 THEN
            sigmoid_f := 1;
        ELSIF x =- 16068 THEN
            sigmoid_f := 1;
        ELSIF x =- 16067 THEN
            sigmoid_f := 1;
        ELSIF x =- 16066 THEN
            sigmoid_f := 1;
        ELSIF x =- 16065 THEN
            sigmoid_f := 1;
        ELSIF x =- 16064 THEN
            sigmoid_f := 1;
        ELSIF x =- 16063 THEN
            sigmoid_f := 1;
        ELSIF x =- 16062 THEN
            sigmoid_f := 1;
        ELSIF x =- 16061 THEN
            sigmoid_f := 1;
        ELSIF x =- 16060 THEN
            sigmoid_f := 1;
        ELSIF x =- 16059 THEN
            sigmoid_f := 1;
        ELSIF x =- 16058 THEN
            sigmoid_f := 1;
        ELSIF x =- 16057 THEN
            sigmoid_f := 1;
        ELSIF x =- 16056 THEN
            sigmoid_f := 1;
        ELSIF x =- 16055 THEN
            sigmoid_f := 1;
        ELSIF x =- 16054 THEN
            sigmoid_f := 1;
        ELSIF x =- 16053 THEN
            sigmoid_f := 1;
        ELSIF x =- 16052 THEN
            sigmoid_f := 1;
        ELSIF x =- 16051 THEN
            sigmoid_f := 1;
        ELSIF x =- 16050 THEN
            sigmoid_f := 1;
        ELSIF x =- 16049 THEN
            sigmoid_f := 1;
        ELSIF x =- 16048 THEN
            sigmoid_f := 1;
        ELSIF x =- 16047 THEN
            sigmoid_f := 1;
        ELSIF x =- 16046 THEN
            sigmoid_f := 1;
        ELSIF x =- 16045 THEN
            sigmoid_f := 1;
        ELSIF x =- 16044 THEN
            sigmoid_f := 1;
        ELSIF x =- 16043 THEN
            sigmoid_f := 1;
        ELSIF x =- 16042 THEN
            sigmoid_f := 1;
        ELSIF x =- 16041 THEN
            sigmoid_f := 1;
        ELSIF x =- 16040 THEN
            sigmoid_f := 1;
        ELSIF x =- 16039 THEN
            sigmoid_f := 1;
        ELSIF x =- 16038 THEN
            sigmoid_f := 1;
        ELSIF x =- 16037 THEN
            sigmoid_f := 1;
        ELSIF x =- 16036 THEN
            sigmoid_f := 1;
        ELSIF x =- 16035 THEN
            sigmoid_f := 1;
        ELSIF x =- 16034 THEN
            sigmoid_f := 1;
        ELSIF x =- 16033 THEN
            sigmoid_f := 1;
        ELSIF x =- 16032 THEN
            sigmoid_f := 1;
        ELSIF x =- 16031 THEN
            sigmoid_f := 1;
        ELSIF x =- 16030 THEN
            sigmoid_f := 1;
        ELSIF x =- 16029 THEN
            sigmoid_f := 1;
        ELSIF x =- 16028 THEN
            sigmoid_f := 1;
        ELSIF x =- 16027 THEN
            sigmoid_f := 1;
        ELSIF x =- 16026 THEN
            sigmoid_f := 1;
        ELSIF x =- 16025 THEN
            sigmoid_f := 1;
        ELSIF x =- 16024 THEN
            sigmoid_f := 1;
        ELSIF x =- 16023 THEN
            sigmoid_f := 1;
        ELSIF x =- 16022 THEN
            sigmoid_f := 1;
        ELSIF x =- 16021 THEN
            sigmoid_f := 1;
        ELSIF x =- 16020 THEN
            sigmoid_f := 1;
        ELSIF x =- 16019 THEN
            sigmoid_f := 1;
        ELSIF x =- 16018 THEN
            sigmoid_f := 1;
        ELSIF x =- 16017 THEN
            sigmoid_f := 1;
        ELSIF x =- 16016 THEN
            sigmoid_f := 1;
        ELSIF x =- 16015 THEN
            sigmoid_f := 1;
        ELSIF x =- 16014 THEN
            sigmoid_f := 1;
        ELSIF x =- 16013 THEN
            sigmoid_f := 1;
        ELSIF x =- 16012 THEN
            sigmoid_f := 1;
        ELSIF x =- 16011 THEN
            sigmoid_f := 1;
        ELSIF x =- 16010 THEN
            sigmoid_f := 1;
        ELSIF x =- 16009 THEN
            sigmoid_f := 1;
        ELSIF x =- 16008 THEN
            sigmoid_f := 1;
        ELSIF x =- 16007 THEN
            sigmoid_f := 1;
        ELSIF x =- 16006 THEN
            sigmoid_f := 1;
        ELSIF x =- 16005 THEN
            sigmoid_f := 1;
        ELSIF x =- 16004 THEN
            sigmoid_f := 1;
        ELSIF x =- 16003 THEN
            sigmoid_f := 1;
        ELSIF x =- 16002 THEN
            sigmoid_f := 1;
        ELSIF x =- 16001 THEN
            sigmoid_f := 1;
        ELSIF x =- 16000 THEN
            sigmoid_f := 1;
        ELSIF x =- 15999 THEN
            sigmoid_f := 1;
        ELSIF x =- 15998 THEN
            sigmoid_f := 1;
        ELSIF x =- 15997 THEN
            sigmoid_f := 1;
        ELSIF x =- 15996 THEN
            sigmoid_f := 1;
        ELSIF x =- 15995 THEN
            sigmoid_f := 1;
        ELSIF x =- 15994 THEN
            sigmoid_f := 1;
        ELSIF x =- 15993 THEN
            sigmoid_f := 1;
        ELSIF x =- 15992 THEN
            sigmoid_f := 1;
        ELSIF x =- 15991 THEN
            sigmoid_f := 1;
        ELSIF x =- 15990 THEN
            sigmoid_f := 1;
        ELSIF x =- 15989 THEN
            sigmoid_f := 1;
        ELSIF x =- 15988 THEN
            sigmoid_f := 1;
        ELSIF x =- 15987 THEN
            sigmoid_f := 1;
        ELSIF x =- 15986 THEN
            sigmoid_f := 1;
        ELSIF x =- 15985 THEN
            sigmoid_f := 1;
        ELSIF x =- 15984 THEN
            sigmoid_f := 1;
        ELSIF x =- 15983 THEN
            sigmoid_f := 1;
        ELSIF x =- 15982 THEN
            sigmoid_f := 1;
        ELSIF x =- 15981 THEN
            sigmoid_f := 1;
        ELSIF x =- 15980 THEN
            sigmoid_f := 1;
        ELSIF x =- 15979 THEN
            sigmoid_f := 1;
        ELSIF x =- 15978 THEN
            sigmoid_f := 1;
        ELSIF x =- 15977 THEN
            sigmoid_f := 1;
        ELSIF x =- 15976 THEN
            sigmoid_f := 1;
        ELSIF x =- 15975 THEN
            sigmoid_f := 1;
        ELSIF x =- 15974 THEN
            sigmoid_f := 1;
        ELSIF x =- 15973 THEN
            sigmoid_f := 1;
        ELSIF x =- 15972 THEN
            sigmoid_f := 1;
        ELSIF x =- 15971 THEN
            sigmoid_f := 1;
        ELSIF x =- 15970 THEN
            sigmoid_f := 1;
        ELSIF x =- 15969 THEN
            sigmoid_f := 1;
        ELSIF x =- 15968 THEN
            sigmoid_f := 1;
        ELSIF x =- 15967 THEN
            sigmoid_f := 1;
        ELSIF x =- 15966 THEN
            sigmoid_f := 1;
        ELSIF x =- 15965 THEN
            sigmoid_f := 1;
        ELSIF x =- 15964 THEN
            sigmoid_f := 1;
        ELSIF x =- 15963 THEN
            sigmoid_f := 1;
        ELSIF x =- 15962 THEN
            sigmoid_f := 1;
        ELSIF x =- 15961 THEN
            sigmoid_f := 1;
        ELSIF x =- 15960 THEN
            sigmoid_f := 1;
        ELSIF x =- 15959 THEN
            sigmoid_f := 1;
        ELSIF x =- 15958 THEN
            sigmoid_f := 1;
        ELSIF x =- 15957 THEN
            sigmoid_f := 1;
        ELSIF x =- 15956 THEN
            sigmoid_f := 1;
        ELSIF x =- 15955 THEN
            sigmoid_f := 1;
        ELSIF x =- 15954 THEN
            sigmoid_f := 1;
        ELSIF x =- 15953 THEN
            sigmoid_f := 1;
        ELSIF x =- 15952 THEN
            sigmoid_f := 1;
        ELSIF x =- 15951 THEN
            sigmoid_f := 1;
        ELSIF x =- 15950 THEN
            sigmoid_f := 1;
        ELSIF x =- 15949 THEN
            sigmoid_f := 1;
        ELSIF x =- 15948 THEN
            sigmoid_f := 1;
        ELSIF x =- 15947 THEN
            sigmoid_f := 1;
        ELSIF x =- 15946 THEN
            sigmoid_f := 1;
        ELSIF x =- 15945 THEN
            sigmoid_f := 1;
        ELSIF x =- 15944 THEN
            sigmoid_f := 1;
        ELSIF x =- 15943 THEN
            sigmoid_f := 1;
        ELSIF x =- 15942 THEN
            sigmoid_f := 1;
        ELSIF x =- 15941 THEN
            sigmoid_f := 1;
        ELSIF x =- 15940 THEN
            sigmoid_f := 1;
        ELSIF x =- 15939 THEN
            sigmoid_f := 1;
        ELSIF x =- 15938 THEN
            sigmoid_f := 1;
        ELSIF x =- 15937 THEN
            sigmoid_f := 1;
        ELSIF x =- 15936 THEN
            sigmoid_f := 1;
        ELSIF x =- 15935 THEN
            sigmoid_f := 1;
        ELSIF x =- 15934 THEN
            sigmoid_f := 1;
        ELSIF x =- 15933 THEN
            sigmoid_f := 1;
        ELSIF x =- 15932 THEN
            sigmoid_f := 1;
        ELSIF x =- 15931 THEN
            sigmoid_f := 1;
        ELSIF x =- 15930 THEN
            sigmoid_f := 1;
        ELSIF x =- 15929 THEN
            sigmoid_f := 1;
        ELSIF x =- 15928 THEN
            sigmoid_f := 1;
        ELSIF x =- 15927 THEN
            sigmoid_f := 1;
        ELSIF x =- 15926 THEN
            sigmoid_f := 1;
        ELSIF x =- 15925 THEN
            sigmoid_f := 1;
        ELSIF x =- 15924 THEN
            sigmoid_f := 1;
        ELSIF x =- 15923 THEN
            sigmoid_f := 1;
        ELSIF x =- 15922 THEN
            sigmoid_f := 1;
        ELSIF x =- 15921 THEN
            sigmoid_f := 1;
        ELSIF x =- 15920 THEN
            sigmoid_f := 1;
        ELSIF x =- 15919 THEN
            sigmoid_f := 1;
        ELSIF x =- 15918 THEN
            sigmoid_f := 1;
        ELSIF x =- 15917 THEN
            sigmoid_f := 1;
        ELSIF x =- 15916 THEN
            sigmoid_f := 1;
        ELSIF x =- 15915 THEN
            sigmoid_f := 1;
        ELSIF x =- 15914 THEN
            sigmoid_f := 1;
        ELSIF x =- 15913 THEN
            sigmoid_f := 1;
        ELSIF x =- 15912 THEN
            sigmoid_f := 1;
        ELSIF x =- 15911 THEN
            sigmoid_f := 1;
        ELSIF x =- 15910 THEN
            sigmoid_f := 1;
        ELSIF x =- 15909 THEN
            sigmoid_f := 1;
        ELSIF x =- 15908 THEN
            sigmoid_f := 1;
        ELSIF x =- 15907 THEN
            sigmoid_f := 1;
        ELSIF x =- 15906 THEN
            sigmoid_f := 1;
        ELSIF x =- 15905 THEN
            sigmoid_f := 1;
        ELSIF x =- 15904 THEN
            sigmoid_f := 1;
        ELSIF x =- 15903 THEN
            sigmoid_f := 1;
        ELSIF x =- 15902 THEN
            sigmoid_f := 1;
        ELSIF x =- 15901 THEN
            sigmoid_f := 1;
        ELSIF x =- 15900 THEN
            sigmoid_f := 1;
        ELSIF x =- 15899 THEN
            sigmoid_f := 1;
        ELSIF x =- 15898 THEN
            sigmoid_f := 1;
        ELSIF x =- 15897 THEN
            sigmoid_f := 1;
        ELSIF x =- 15896 THEN
            sigmoid_f := 1;
        ELSIF x =- 15895 THEN
            sigmoid_f := 1;
        ELSIF x =- 15894 THEN
            sigmoid_f := 1;
        ELSIF x =- 15893 THEN
            sigmoid_f := 1;
        ELSIF x =- 15892 THEN
            sigmoid_f := 1;
        ELSIF x =- 15891 THEN
            sigmoid_f := 1;
        ELSIF x =- 15890 THEN
            sigmoid_f := 1;
        ELSIF x =- 15889 THEN
            sigmoid_f := 1;
        ELSIF x =- 15888 THEN
            sigmoid_f := 1;
        ELSIF x =- 15887 THEN
            sigmoid_f := 1;
        ELSIF x =- 15886 THEN
            sigmoid_f := 1;
        ELSIF x =- 15885 THEN
            sigmoid_f := 1;
        ELSIF x =- 15884 THEN
            sigmoid_f := 1;
        ELSIF x =- 15883 THEN
            sigmoid_f := 1;
        ELSIF x =- 15882 THEN
            sigmoid_f := 1;
        ELSIF x =- 15881 THEN
            sigmoid_f := 1;
        ELSIF x =- 15880 THEN
            sigmoid_f := 1;
        ELSIF x =- 15879 THEN
            sigmoid_f := 1;
        ELSIF x =- 15878 THEN
            sigmoid_f := 1;
        ELSIF x =- 15877 THEN
            sigmoid_f := 1;
        ELSIF x =- 15876 THEN
            sigmoid_f := 1;
        ELSIF x =- 15875 THEN
            sigmoid_f := 1;
        ELSIF x =- 15874 THEN
            sigmoid_f := 1;
        ELSIF x =- 15873 THEN
            sigmoid_f := 1;
        ELSIF x =- 15872 THEN
            sigmoid_f := 1;
        ELSIF x =- 15871 THEN
            sigmoid_f := 1;
        ELSIF x =- 15870 THEN
            sigmoid_f := 1;
        ELSIF x =- 15869 THEN
            sigmoid_f := 1;
        ELSIF x =- 15868 THEN
            sigmoid_f := 1;
        ELSIF x =- 15867 THEN
            sigmoid_f := 1;
        ELSIF x =- 15866 THEN
            sigmoid_f := 1;
        ELSIF x =- 15865 THEN
            sigmoid_f := 1;
        ELSIF x =- 15864 THEN
            sigmoid_f := 1;
        ELSIF x =- 15863 THEN
            sigmoid_f := 1;
        ELSIF x =- 15862 THEN
            sigmoid_f := 1;
        ELSIF x =- 15861 THEN
            sigmoid_f := 1;
        ELSIF x =- 15860 THEN
            sigmoid_f := 1;
        ELSIF x =- 15859 THEN
            sigmoid_f := 1;
        ELSIF x =- 15858 THEN
            sigmoid_f := 1;
        ELSIF x =- 15857 THEN
            sigmoid_f := 1;
        ELSIF x =- 15856 THEN
            sigmoid_f := 1;
        ELSIF x =- 15855 THEN
            sigmoid_f := 1;
        ELSIF x =- 15854 THEN
            sigmoid_f := 1;
        ELSIF x =- 15853 THEN
            sigmoid_f := 1;
        ELSIF x =- 15852 THEN
            sigmoid_f := 1;
        ELSIF x =- 15851 THEN
            sigmoid_f := 1;
        ELSIF x =- 15850 THEN
            sigmoid_f := 1;
        ELSIF x =- 15849 THEN
            sigmoid_f := 1;
        ELSIF x =- 15848 THEN
            sigmoid_f := 1;
        ELSIF x =- 15847 THEN
            sigmoid_f := 1;
        ELSIF x =- 15846 THEN
            sigmoid_f := 1;
        ELSIF x =- 15845 THEN
            sigmoid_f := 1;
        ELSIF x =- 15844 THEN
            sigmoid_f := 1;
        ELSIF x =- 15843 THEN
            sigmoid_f := 1;
        ELSIF x =- 15842 THEN
            sigmoid_f := 1;
        ELSIF x =- 15841 THEN
            sigmoid_f := 1;
        ELSIF x =- 15840 THEN
            sigmoid_f := 1;
        ELSIF x =- 15839 THEN
            sigmoid_f := 1;
        ELSIF x =- 15838 THEN
            sigmoid_f := 1;
        ELSIF x =- 15837 THEN
            sigmoid_f := 1;
        ELSIF x =- 15836 THEN
            sigmoid_f := 1;
        ELSIF x =- 15835 THEN
            sigmoid_f := 1;
        ELSIF x =- 15834 THEN
            sigmoid_f := 1;
        ELSIF x =- 15833 THEN
            sigmoid_f := 1;
        ELSIF x =- 15832 THEN
            sigmoid_f := 1;
        ELSIF x =- 15831 THEN
            sigmoid_f := 1;
        ELSIF x =- 15830 THEN
            sigmoid_f := 1;
        ELSIF x =- 15829 THEN
            sigmoid_f := 1;
        ELSIF x =- 15828 THEN
            sigmoid_f := 1;
        ELSIF x =- 15827 THEN
            sigmoid_f := 1;
        ELSIF x =- 15826 THEN
            sigmoid_f := 1;
        ELSIF x =- 15825 THEN
            sigmoid_f := 1;
        ELSIF x =- 15824 THEN
            sigmoid_f := 1;
        ELSIF x =- 15823 THEN
            sigmoid_f := 1;
        ELSIF x =- 15822 THEN
            sigmoid_f := 1;
        ELSIF x =- 15821 THEN
            sigmoid_f := 1;
        ELSIF x =- 15820 THEN
            sigmoid_f := 1;
        ELSIF x =- 15819 THEN
            sigmoid_f := 1;
        ELSIF x =- 15818 THEN
            sigmoid_f := 1;
        ELSIF x =- 15817 THEN
            sigmoid_f := 1;
        ELSIF x =- 15816 THEN
            sigmoid_f := 1;
        ELSIF x =- 15815 THEN
            sigmoid_f := 1;
        ELSIF x =- 15814 THEN
            sigmoid_f := 1;
        ELSIF x =- 15813 THEN
            sigmoid_f := 1;
        ELSIF x =- 15812 THEN
            sigmoid_f := 1;
        ELSIF x =- 15811 THEN
            sigmoid_f := 1;
        ELSIF x =- 15810 THEN
            sigmoid_f := 1;
        ELSIF x =- 15809 THEN
            sigmoid_f := 1;
        ELSIF x =- 15808 THEN
            sigmoid_f := 1;
        ELSIF x =- 15807 THEN
            sigmoid_f := 1;
        ELSIF x =- 15806 THEN
            sigmoid_f := 1;
        ELSIF x =- 15805 THEN
            sigmoid_f := 1;
        ELSIF x =- 15804 THEN
            sigmoid_f := 1;
        ELSIF x =- 15803 THEN
            sigmoid_f := 1;
        ELSIF x =- 15802 THEN
            sigmoid_f := 1;
        ELSIF x =- 15801 THEN
            sigmoid_f := 1;
        ELSIF x =- 15800 THEN
            sigmoid_f := 1;
        ELSIF x =- 15799 THEN
            sigmoid_f := 1;
        ELSIF x =- 15798 THEN
            sigmoid_f := 1;
        ELSIF x =- 15797 THEN
            sigmoid_f := 1;
        ELSIF x =- 15796 THEN
            sigmoid_f := 1;
        ELSIF x =- 15795 THEN
            sigmoid_f := 1;
        ELSIF x =- 15794 THEN
            sigmoid_f := 1;
        ELSIF x =- 15793 THEN
            sigmoid_f := 1;
        ELSIF x =- 15792 THEN
            sigmoid_f := 1;
        ELSIF x =- 15791 THEN
            sigmoid_f := 1;
        ELSIF x =- 15790 THEN
            sigmoid_f := 1;
        ELSIF x =- 15789 THEN
            sigmoid_f := 1;
        ELSIF x =- 15788 THEN
            sigmoid_f := 1;
        ELSIF x =- 15787 THEN
            sigmoid_f := 1;
        ELSIF x =- 15786 THEN
            sigmoid_f := 1;
        ELSIF x =- 15785 THEN
            sigmoid_f := 1;
        ELSIF x =- 15784 THEN
            sigmoid_f := 1;
        ELSIF x =- 15783 THEN
            sigmoid_f := 1;
        ELSIF x =- 15782 THEN
            sigmoid_f := 1;
        ELSIF x =- 15781 THEN
            sigmoid_f := 1;
        ELSIF x =- 15780 THEN
            sigmoid_f := 1;
        ELSIF x =- 15779 THEN
            sigmoid_f := 1;
        ELSIF x =- 15778 THEN
            sigmoid_f := 1;
        ELSIF x =- 15777 THEN
            sigmoid_f := 1;
        ELSIF x =- 15776 THEN
            sigmoid_f := 1;
        ELSIF x =- 15775 THEN
            sigmoid_f := 1;
        ELSIF x =- 15774 THEN
            sigmoid_f := 1;
        ELSIF x =- 15773 THEN
            sigmoid_f := 1;
        ELSIF x =- 15772 THEN
            sigmoid_f := 1;
        ELSIF x =- 15771 THEN
            sigmoid_f := 1;
        ELSIF x =- 15770 THEN
            sigmoid_f := 1;
        ELSIF x =- 15769 THEN
            sigmoid_f := 1;
        ELSIF x =- 15768 THEN
            sigmoid_f := 1;
        ELSIF x =- 15767 THEN
            sigmoid_f := 1;
        ELSIF x =- 15766 THEN
            sigmoid_f := 1;
        ELSIF x =- 15765 THEN
            sigmoid_f := 1;
        ELSIF x =- 15764 THEN
            sigmoid_f := 1;
        ELSIF x =- 15763 THEN
            sigmoid_f := 1;
        ELSIF x =- 15762 THEN
            sigmoid_f := 1;
        ELSIF x =- 15761 THEN
            sigmoid_f := 1;
        ELSIF x =- 15760 THEN
            sigmoid_f := 1;
        ELSIF x =- 15759 THEN
            sigmoid_f := 1;
        ELSIF x =- 15758 THEN
            sigmoid_f := 1;
        ELSIF x =- 15757 THEN
            sigmoid_f := 1;
        ELSIF x =- 15756 THEN
            sigmoid_f := 1;
        ELSIF x =- 15755 THEN
            sigmoid_f := 1;
        ELSIF x =- 15754 THEN
            sigmoid_f := 1;
        ELSIF x =- 15753 THEN
            sigmoid_f := 1;
        ELSIF x =- 15752 THEN
            sigmoid_f := 1;
        ELSIF x =- 15751 THEN
            sigmoid_f := 1;
        ELSIF x =- 15750 THEN
            sigmoid_f := 1;
        ELSIF x =- 15749 THEN
            sigmoid_f := 1;
        ELSIF x =- 15748 THEN
            sigmoid_f := 1;
        ELSIF x =- 15747 THEN
            sigmoid_f := 1;
        ELSIF x =- 15746 THEN
            sigmoid_f := 1;
        ELSIF x =- 15745 THEN
            sigmoid_f := 1;
        ELSIF x =- 15744 THEN
            sigmoid_f := 1;
        ELSIF x =- 15743 THEN
            sigmoid_f := 1;
        ELSIF x =- 15742 THEN
            sigmoid_f := 1;
        ELSIF x =- 15741 THEN
            sigmoid_f := 1;
        ELSIF x =- 15740 THEN
            sigmoid_f := 1;
        ELSIF x =- 15739 THEN
            sigmoid_f := 1;
        ELSIF x =- 15738 THEN
            sigmoid_f := 1;
        ELSIF x =- 15737 THEN
            sigmoid_f := 1;
        ELSIF x =- 15736 THEN
            sigmoid_f := 1;
        ELSIF x =- 15735 THEN
            sigmoid_f := 1;
        ELSIF x =- 15734 THEN
            sigmoid_f := 1;
        ELSIF x =- 15733 THEN
            sigmoid_f := 1;
        ELSIF x =- 15732 THEN
            sigmoid_f := 1;
        ELSIF x =- 15731 THEN
            sigmoid_f := 1;
        ELSIF x =- 15730 THEN
            sigmoid_f := 1;
        ELSIF x =- 15729 THEN
            sigmoid_f := 1;
        ELSIF x =- 15728 THEN
            sigmoid_f := 1;
        ELSIF x =- 15727 THEN
            sigmoid_f := 1;
        ELSIF x =- 15726 THEN
            sigmoid_f := 1;
        ELSIF x =- 15725 THEN
            sigmoid_f := 1;
        ELSIF x =- 15724 THEN
            sigmoid_f := 1;
        ELSIF x =- 15723 THEN
            sigmoid_f := 1;
        ELSIF x =- 15722 THEN
            sigmoid_f := 1;
        ELSIF x =- 15721 THEN
            sigmoid_f := 1;
        ELSIF x =- 15720 THEN
            sigmoid_f := 1;
        ELSIF x =- 15719 THEN
            sigmoid_f := 1;
        ELSIF x =- 15718 THEN
            sigmoid_f := 1;
        ELSIF x =- 15717 THEN
            sigmoid_f := 1;
        ELSIF x =- 15716 THEN
            sigmoid_f := 1;
        ELSIF x =- 15715 THEN
            sigmoid_f := 1;
        ELSIF x =- 15714 THEN
            sigmoid_f := 1;
        ELSIF x =- 15713 THEN
            sigmoid_f := 1;
        ELSIF x =- 15712 THEN
            sigmoid_f := 1;
        ELSIF x =- 15711 THEN
            sigmoid_f := 1;
        ELSIF x =- 15710 THEN
            sigmoid_f := 1;
        ELSIF x =- 15709 THEN
            sigmoid_f := 1;
        ELSIF x =- 15708 THEN
            sigmoid_f := 1;
        ELSIF x =- 15707 THEN
            sigmoid_f := 1;
        ELSIF x =- 15706 THEN
            sigmoid_f := 1;
        ELSIF x =- 15705 THEN
            sigmoid_f := 1;
        ELSIF x =- 15704 THEN
            sigmoid_f := 1;
        ELSIF x =- 15703 THEN
            sigmoid_f := 1;
        ELSIF x =- 15702 THEN
            sigmoid_f := 1;
        ELSIF x =- 15701 THEN
            sigmoid_f := 1;
        ELSIF x =- 15700 THEN
            sigmoid_f := 1;
        ELSIF x =- 15699 THEN
            sigmoid_f := 1;
        ELSIF x =- 15698 THEN
            sigmoid_f := 1;
        ELSIF x =- 15697 THEN
            sigmoid_f := 1;
        ELSIF x =- 15696 THEN
            sigmoid_f := 1;
        ELSIF x =- 15695 THEN
            sigmoid_f := 1;
        ELSIF x =- 15694 THEN
            sigmoid_f := 1;
        ELSIF x =- 15693 THEN
            sigmoid_f := 1;
        ELSIF x =- 15692 THEN
            sigmoid_f := 1;
        ELSIF x =- 15691 THEN
            sigmoid_f := 1;
        ELSIF x =- 15690 THEN
            sigmoid_f := 1;
        ELSIF x =- 15689 THEN
            sigmoid_f := 1;
        ELSIF x =- 15688 THEN
            sigmoid_f := 1;
        ELSIF x =- 15687 THEN
            sigmoid_f := 1;
        ELSIF x =- 15686 THEN
            sigmoid_f := 1;
        ELSIF x =- 15685 THEN
            sigmoid_f := 1;
        ELSIF x =- 15684 THEN
            sigmoid_f := 1;
        ELSIF x =- 15683 THEN
            sigmoid_f := 1;
        ELSIF x =- 15682 THEN
            sigmoid_f := 1;
        ELSIF x =- 15681 THEN
            sigmoid_f := 1;
        ELSIF x =- 15680 THEN
            sigmoid_f := 1;
        ELSIF x =- 15679 THEN
            sigmoid_f := 1;
        ELSIF x =- 15678 THEN
            sigmoid_f := 1;
        ELSIF x =- 15677 THEN
            sigmoid_f := 1;
        ELSIF x =- 15676 THEN
            sigmoid_f := 1;
        ELSIF x =- 15675 THEN
            sigmoid_f := 1;
        ELSIF x =- 15674 THEN
            sigmoid_f := 1;
        ELSIF x =- 15673 THEN
            sigmoid_f := 1;
        ELSIF x =- 15672 THEN
            sigmoid_f := 1;
        ELSIF x =- 15671 THEN
            sigmoid_f := 1;
        ELSIF x =- 15670 THEN
            sigmoid_f := 1;
        ELSIF x =- 15669 THEN
            sigmoid_f := 1;
        ELSIF x =- 15668 THEN
            sigmoid_f := 1;
        ELSIF x =- 15667 THEN
            sigmoid_f := 1;
        ELSIF x =- 15666 THEN
            sigmoid_f := 1;
        ELSIF x =- 15665 THEN
            sigmoid_f := 1;
        ELSIF x =- 15664 THEN
            sigmoid_f := 1;
        ELSIF x =- 15663 THEN
            sigmoid_f := 1;
        ELSIF x =- 15662 THEN
            sigmoid_f := 1;
        ELSIF x =- 15661 THEN
            sigmoid_f := 1;
        ELSIF x =- 15660 THEN
            sigmoid_f := 1;
        ELSIF x =- 15659 THEN
            sigmoid_f := 1;
        ELSIF x =- 15658 THEN
            sigmoid_f := 1;
        ELSIF x =- 15657 THEN
            sigmoid_f := 1;
        ELSIF x =- 15656 THEN
            sigmoid_f := 1;
        ELSIF x =- 15655 THEN
            sigmoid_f := 1;
        ELSIF x =- 15654 THEN
            sigmoid_f := 1;
        ELSIF x =- 15653 THEN
            sigmoid_f := 1;
        ELSIF x =- 15652 THEN
            sigmoid_f := 1;
        ELSIF x =- 15651 THEN
            sigmoid_f := 1;
        ELSIF x =- 15650 THEN
            sigmoid_f := 1;
        ELSIF x =- 15649 THEN
            sigmoid_f := 1;
        ELSIF x =- 15648 THEN
            sigmoid_f := 1;
        ELSIF x =- 15647 THEN
            sigmoid_f := 1;
        ELSIF x =- 15646 THEN
            sigmoid_f := 1;
        ELSIF x =- 15645 THEN
            sigmoid_f := 1;
        ELSIF x =- 15644 THEN
            sigmoid_f := 1;
        ELSIF x =- 15643 THEN
            sigmoid_f := 1;
        ELSIF x =- 15642 THEN
            sigmoid_f := 1;
        ELSIF x =- 15641 THEN
            sigmoid_f := 1;
        ELSIF x =- 15640 THEN
            sigmoid_f := 1;
        ELSIF x =- 15639 THEN
            sigmoid_f := 1;
        ELSIF x =- 15638 THEN
            sigmoid_f := 1;
        ELSIF x =- 15637 THEN
            sigmoid_f := 1;
        ELSIF x =- 15636 THEN
            sigmoid_f := 1;
        ELSIF x =- 15635 THEN
            sigmoid_f := 1;
        ELSIF x =- 15634 THEN
            sigmoid_f := 1;
        ELSIF x =- 15633 THEN
            sigmoid_f := 1;
        ELSIF x =- 15632 THEN
            sigmoid_f := 1;
        ELSIF x =- 15631 THEN
            sigmoid_f := 1;
        ELSIF x =- 15630 THEN
            sigmoid_f := 1;
        ELSIF x =- 15629 THEN
            sigmoid_f := 1;
        ELSIF x =- 15628 THEN
            sigmoid_f := 1;
        ELSIF x =- 15627 THEN
            sigmoid_f := 1;
        ELSIF x =- 15626 THEN
            sigmoid_f := 1;
        ELSIF x =- 15625 THEN
            sigmoid_f := 1;
        ELSIF x =- 15624 THEN
            sigmoid_f := 1;
        ELSIF x =- 15623 THEN
            sigmoid_f := 1;
        ELSIF x =- 15622 THEN
            sigmoid_f := 1;
        ELSIF x =- 15621 THEN
            sigmoid_f := 1;
        ELSIF x =- 15620 THEN
            sigmoid_f := 1;
        ELSIF x =- 15619 THEN
            sigmoid_f := 1;
        ELSIF x =- 15618 THEN
            sigmoid_f := 1;
        ELSIF x =- 15617 THEN
            sigmoid_f := 1;
        ELSIF x =- 15616 THEN
            sigmoid_f := 1;
        ELSIF x =- 15615 THEN
            sigmoid_f := 1;
        ELSIF x =- 15614 THEN
            sigmoid_f := 1;
        ELSIF x =- 15613 THEN
            sigmoid_f := 1;
        ELSIF x =- 15612 THEN
            sigmoid_f := 1;
        ELSIF x =- 15611 THEN
            sigmoid_f := 1;
        ELSIF x =- 15610 THEN
            sigmoid_f := 1;
        ELSIF x =- 15609 THEN
            sigmoid_f := 1;
        ELSIF x =- 15608 THEN
            sigmoid_f := 1;
        ELSIF x =- 15607 THEN
            sigmoid_f := 1;
        ELSIF x =- 15606 THEN
            sigmoid_f := 1;
        ELSIF x =- 15605 THEN
            sigmoid_f := 1;
        ELSIF x =- 15604 THEN
            sigmoid_f := 1;
        ELSIF x =- 15603 THEN
            sigmoid_f := 1;
        ELSIF x =- 15602 THEN
            sigmoid_f := 1;
        ELSIF x =- 15601 THEN
            sigmoid_f := 1;
        ELSIF x =- 15600 THEN
            sigmoid_f := 1;
        ELSIF x =- 15599 THEN
            sigmoid_f := 1;
        ELSIF x =- 15598 THEN
            sigmoid_f := 1;
        ELSIF x =- 15597 THEN
            sigmoid_f := 1;
        ELSIF x =- 15596 THEN
            sigmoid_f := 1;
        ELSIF x =- 15595 THEN
            sigmoid_f := 1;
        ELSIF x =- 15594 THEN
            sigmoid_f := 1;
        ELSIF x =- 15593 THEN
            sigmoid_f := 1;
        ELSIF x =- 15592 THEN
            sigmoid_f := 1;
        ELSIF x =- 15591 THEN
            sigmoid_f := 1;
        ELSIF x =- 15590 THEN
            sigmoid_f := 1;
        ELSIF x =- 15589 THEN
            sigmoid_f := 1;
        ELSIF x =- 15588 THEN
            sigmoid_f := 1;
        ELSIF x =- 15587 THEN
            sigmoid_f := 1;
        ELSIF x =- 15586 THEN
            sigmoid_f := 1;
        ELSIF x =- 15585 THEN
            sigmoid_f := 1;
        ELSIF x =- 15584 THEN
            sigmoid_f := 1;
        ELSIF x =- 15583 THEN
            sigmoid_f := 1;
        ELSIF x =- 15582 THEN
            sigmoid_f := 1;
        ELSIF x =- 15581 THEN
            sigmoid_f := 1;
        ELSIF x =- 15580 THEN
            sigmoid_f := 1;
        ELSIF x =- 15579 THEN
            sigmoid_f := 1;
        ELSIF x =- 15578 THEN
            sigmoid_f := 1;
        ELSIF x =- 15577 THEN
            sigmoid_f := 1;
        ELSIF x =- 15576 THEN
            sigmoid_f := 1;
        ELSIF x =- 15575 THEN
            sigmoid_f := 1;
        ELSIF x =- 15574 THEN
            sigmoid_f := 1;
        ELSIF x =- 15573 THEN
            sigmoid_f := 1;
        ELSIF x =- 15572 THEN
            sigmoid_f := 1;
        ELSIF x =- 15571 THEN
            sigmoid_f := 1;
        ELSIF x =- 15570 THEN
            sigmoid_f := 1;
        ELSIF x =- 15569 THEN
            sigmoid_f := 1;
        ELSIF x =- 15568 THEN
            sigmoid_f := 1;
        ELSIF x =- 15567 THEN
            sigmoid_f := 1;
        ELSIF x =- 15566 THEN
            sigmoid_f := 1;
        ELSIF x =- 15565 THEN
            sigmoid_f := 1;
        ELSIF x =- 15564 THEN
            sigmoid_f := 1;
        ELSIF x =- 15563 THEN
            sigmoid_f := 1;
        ELSIF x =- 15562 THEN
            sigmoid_f := 1;
        ELSIF x =- 15561 THEN
            sigmoid_f := 1;
        ELSIF x =- 15560 THEN
            sigmoid_f := 1;
        ELSIF x =- 15559 THEN
            sigmoid_f := 1;
        ELSIF x =- 15558 THEN
            sigmoid_f := 1;
        ELSIF x =- 15557 THEN
            sigmoid_f := 1;
        ELSIF x =- 15556 THEN
            sigmoid_f := 1;
        ELSIF x =- 15555 THEN
            sigmoid_f := 1;
        ELSIF x =- 15554 THEN
            sigmoid_f := 1;
        ELSIF x =- 15553 THEN
            sigmoid_f := 1;
        ELSIF x =- 15552 THEN
            sigmoid_f := 1;
        ELSIF x =- 15551 THEN
            sigmoid_f := 1;
        ELSIF x =- 15550 THEN
            sigmoid_f := 1;
        ELSIF x =- 15549 THEN
            sigmoid_f := 1;
        ELSIF x =- 15548 THEN
            sigmoid_f := 1;
        ELSIF x =- 15547 THEN
            sigmoid_f := 1;
        ELSIF x =- 15546 THEN
            sigmoid_f := 1;
        ELSIF x =- 15545 THEN
            sigmoid_f := 1;
        ELSIF x =- 15544 THEN
            sigmoid_f := 1;
        ELSIF x =- 15543 THEN
            sigmoid_f := 1;
        ELSIF x =- 15542 THEN
            sigmoid_f := 1;
        ELSIF x =- 15541 THEN
            sigmoid_f := 1;
        ELSIF x =- 15540 THEN
            sigmoid_f := 1;
        ELSIF x =- 15539 THEN
            sigmoid_f := 1;
        ELSIF x =- 15538 THEN
            sigmoid_f := 1;
        ELSIF x =- 15537 THEN
            sigmoid_f := 1;
        ELSIF x =- 15536 THEN
            sigmoid_f := 1;
        ELSIF x =- 15535 THEN
            sigmoid_f := 1;
        ELSIF x =- 15534 THEN
            sigmoid_f := 1;
        ELSIF x =- 15533 THEN
            sigmoid_f := 1;
        ELSIF x =- 15532 THEN
            sigmoid_f := 1;
        ELSIF x =- 15531 THEN
            sigmoid_f := 1;
        ELSIF x =- 15530 THEN
            sigmoid_f := 1;
        ELSIF x =- 15529 THEN
            sigmoid_f := 1;
        ELSIF x =- 15528 THEN
            sigmoid_f := 1;
        ELSIF x =- 15527 THEN
            sigmoid_f := 1;
        ELSIF x =- 15526 THEN
            sigmoid_f := 1;
        ELSIF x =- 15525 THEN
            sigmoid_f := 1;
        ELSIF x =- 15524 THEN
            sigmoid_f := 1;
        ELSIF x =- 15523 THEN
            sigmoid_f := 1;
        ELSIF x =- 15522 THEN
            sigmoid_f := 1;
        ELSIF x =- 15521 THEN
            sigmoid_f := 1;
        ELSIF x =- 15520 THEN
            sigmoid_f := 1;
        ELSIF x =- 15519 THEN
            sigmoid_f := 1;
        ELSIF x =- 15518 THEN
            sigmoid_f := 1;
        ELSIF x =- 15517 THEN
            sigmoid_f := 1;
        ELSIF x =- 15516 THEN
            sigmoid_f := 1;
        ELSIF x =- 15515 THEN
            sigmoid_f := 1;
        ELSIF x =- 15514 THEN
            sigmoid_f := 1;
        ELSIF x =- 15513 THEN
            sigmoid_f := 1;
        ELSIF x =- 15512 THEN
            sigmoid_f := 1;
        ELSIF x =- 15511 THEN
            sigmoid_f := 1;
        ELSIF x =- 15510 THEN
            sigmoid_f := 1;
        ELSIF x =- 15509 THEN
            sigmoid_f := 1;
        ELSIF x =- 15508 THEN
            sigmoid_f := 1;
        ELSIF x =- 15507 THEN
            sigmoid_f := 1;
        ELSIF x =- 15506 THEN
            sigmoid_f := 1;
        ELSIF x =- 15505 THEN
            sigmoid_f := 1;
        ELSIF x =- 15504 THEN
            sigmoid_f := 1;
        ELSIF x =- 15503 THEN
            sigmoid_f := 1;
        ELSIF x =- 15502 THEN
            sigmoid_f := 1;
        ELSIF x =- 15501 THEN
            sigmoid_f := 1;
        ELSIF x =- 15500 THEN
            sigmoid_f := 1;
        ELSIF x =- 15499 THEN
            sigmoid_f := 1;
        ELSIF x =- 15498 THEN
            sigmoid_f := 1;
        ELSIF x =- 15497 THEN
            sigmoid_f := 1;
        ELSIF x =- 15496 THEN
            sigmoid_f := 1;
        ELSIF x =- 15495 THEN
            sigmoid_f := 1;
        ELSIF x =- 15494 THEN
            sigmoid_f := 1;
        ELSIF x =- 15493 THEN
            sigmoid_f := 1;
        ELSIF x =- 15492 THEN
            sigmoid_f := 1;
        ELSIF x =- 15491 THEN
            sigmoid_f := 1;
        ELSIF x =- 15490 THEN
            sigmoid_f := 1;
        ELSIF x =- 15489 THEN
            sigmoid_f := 1;
        ELSIF x =- 15488 THEN
            sigmoid_f := 1;
        ELSIF x =- 15487 THEN
            sigmoid_f := 1;
        ELSIF x =- 15486 THEN
            sigmoid_f := 1;
        ELSIF x =- 15485 THEN
            sigmoid_f := 1;
        ELSIF x =- 15484 THEN
            sigmoid_f := 1;
        ELSIF x =- 15483 THEN
            sigmoid_f := 1;
        ELSIF x =- 15482 THEN
            sigmoid_f := 1;
        ELSIF x =- 15481 THEN
            sigmoid_f := 1;
        ELSIF x =- 15480 THEN
            sigmoid_f := 1;
        ELSIF x =- 15479 THEN
            sigmoid_f := 1;
        ELSIF x =- 15478 THEN
            sigmoid_f := 1;
        ELSIF x =- 15477 THEN
            sigmoid_f := 1;
        ELSIF x =- 15476 THEN
            sigmoid_f := 1;
        ELSIF x =- 15475 THEN
            sigmoid_f := 1;
        ELSIF x =- 15474 THEN
            sigmoid_f := 1;
        ELSIF x =- 15473 THEN
            sigmoid_f := 1;
        ELSIF x =- 15472 THEN
            sigmoid_f := 1;
        ELSIF x =- 15471 THEN
            sigmoid_f := 1;
        ELSIF x =- 15470 THEN
            sigmoid_f := 1;
        ELSIF x =- 15469 THEN
            sigmoid_f := 1;
        ELSIF x =- 15468 THEN
            sigmoid_f := 1;
        ELSIF x =- 15467 THEN
            sigmoid_f := 1;
        ELSIF x =- 15466 THEN
            sigmoid_f := 1;
        ELSIF x =- 15465 THEN
            sigmoid_f := 1;
        ELSIF x =- 15464 THEN
            sigmoid_f := 1;
        ELSIF x =- 15463 THEN
            sigmoid_f := 1;
        ELSIF x =- 15462 THEN
            sigmoid_f := 1;
        ELSIF x =- 15461 THEN
            sigmoid_f := 1;
        ELSIF x =- 15460 THEN
            sigmoid_f := 1;
        ELSIF x =- 15459 THEN
            sigmoid_f := 1;
        ELSIF x =- 15458 THEN
            sigmoid_f := 1;
        ELSIF x =- 15457 THEN
            sigmoid_f := 1;
        ELSIF x =- 15456 THEN
            sigmoid_f := 1;
        ELSIF x =- 15455 THEN
            sigmoid_f := 1;
        ELSIF x =- 15454 THEN
            sigmoid_f := 1;
        ELSIF x =- 15453 THEN
            sigmoid_f := 1;
        ELSIF x =- 15452 THEN
            sigmoid_f := 1;
        ELSIF x =- 15451 THEN
            sigmoid_f := 1;
        ELSIF x =- 15450 THEN
            sigmoid_f := 1;
        ELSIF x =- 15449 THEN
            sigmoid_f := 1;
        ELSIF x =- 15448 THEN
            sigmoid_f := 1;
        ELSIF x =- 15447 THEN
            sigmoid_f := 1;
        ELSIF x =- 15446 THEN
            sigmoid_f := 1;
        ELSIF x =- 15445 THEN
            sigmoid_f := 1;
        ELSIF x =- 15444 THEN
            sigmoid_f := 1;
        ELSIF x =- 15443 THEN
            sigmoid_f := 1;
        ELSIF x =- 15442 THEN
            sigmoid_f := 1;
        ELSIF x =- 15441 THEN
            sigmoid_f := 1;
        ELSIF x =- 15440 THEN
            sigmoid_f := 1;
        ELSIF x =- 15439 THEN
            sigmoid_f := 1;
        ELSIF x =- 15438 THEN
            sigmoid_f := 1;
        ELSIF x =- 15437 THEN
            sigmoid_f := 1;
        ELSIF x =- 15436 THEN
            sigmoid_f := 1;
        ELSIF x =- 15435 THEN
            sigmoid_f := 1;
        ELSIF x =- 15434 THEN
            sigmoid_f := 1;
        ELSIF x =- 15433 THEN
            sigmoid_f := 1;
        ELSIF x =- 15432 THEN
            sigmoid_f := 1;
        ELSIF x =- 15431 THEN
            sigmoid_f := 1;
        ELSIF x =- 15430 THEN
            sigmoid_f := 1;
        ELSIF x =- 15429 THEN
            sigmoid_f := 1;
        ELSIF x =- 15428 THEN
            sigmoid_f := 1;
        ELSIF x =- 15427 THEN
            sigmoid_f := 1;
        ELSIF x =- 15426 THEN
            sigmoid_f := 1;
        ELSIF x =- 15425 THEN
            sigmoid_f := 1;
        ELSIF x =- 15424 THEN
            sigmoid_f := 1;
        ELSIF x =- 15423 THEN
            sigmoid_f := 1;
        ELSIF x =- 15422 THEN
            sigmoid_f := 1;
        ELSIF x =- 15421 THEN
            sigmoid_f := 1;
        ELSIF x =- 15420 THEN
            sigmoid_f := 1;
        ELSIF x =- 15419 THEN
            sigmoid_f := 1;
        ELSIF x =- 15418 THEN
            sigmoid_f := 1;
        ELSIF x =- 15417 THEN
            sigmoid_f := 1;
        ELSIF x =- 15416 THEN
            sigmoid_f := 1;
        ELSIF x =- 15415 THEN
            sigmoid_f := 1;
        ELSIF x =- 15414 THEN
            sigmoid_f := 1;
        ELSIF x =- 15413 THEN
            sigmoid_f := 1;
        ELSIF x =- 15412 THEN
            sigmoid_f := 1;
        ELSIF x =- 15411 THEN
            sigmoid_f := 1;
        ELSIF x =- 15410 THEN
            sigmoid_f := 1;
        ELSIF x =- 15409 THEN
            sigmoid_f := 1;
        ELSIF x =- 15408 THEN
            sigmoid_f := 1;
        ELSIF x =- 15407 THEN
            sigmoid_f := 1;
        ELSIF x =- 15406 THEN
            sigmoid_f := 1;
        ELSIF x =- 15405 THEN
            sigmoid_f := 1;
        ELSIF x =- 15404 THEN
            sigmoid_f := 1;
        ELSIF x =- 15403 THEN
            sigmoid_f := 1;
        ELSIF x =- 15402 THEN
            sigmoid_f := 1;
        ELSIF x =- 15401 THEN
            sigmoid_f := 1;
        ELSIF x =- 15400 THEN
            sigmoid_f := 1;
        ELSIF x =- 15399 THEN
            sigmoid_f := 1;
        ELSIF x =- 15398 THEN
            sigmoid_f := 1;
        ELSIF x =- 15397 THEN
            sigmoid_f := 1;
        ELSIF x =- 15396 THEN
            sigmoid_f := 1;
        ELSIF x =- 15395 THEN
            sigmoid_f := 1;
        ELSIF x =- 15394 THEN
            sigmoid_f := 1;
        ELSIF x =- 15393 THEN
            sigmoid_f := 1;
        ELSIF x =- 15392 THEN
            sigmoid_f := 1;
        ELSIF x =- 15391 THEN
            sigmoid_f := 1;
        ELSIF x =- 15390 THEN
            sigmoid_f := 1;
        ELSIF x =- 15389 THEN
            sigmoid_f := 1;
        ELSIF x =- 15388 THEN
            sigmoid_f := 1;
        ELSIF x =- 15387 THEN
            sigmoid_f := 1;
        ELSIF x =- 15386 THEN
            sigmoid_f := 1;
        ELSIF x =- 15385 THEN
            sigmoid_f := 1;
        ELSIF x =- 15384 THEN
            sigmoid_f := 1;
        ELSIF x =- 15383 THEN
            sigmoid_f := 1;
        ELSIF x =- 15382 THEN
            sigmoid_f := 1;
        ELSIF x =- 15381 THEN
            sigmoid_f := 1;
        ELSIF x =- 15380 THEN
            sigmoid_f := 1;
        ELSIF x =- 15379 THEN
            sigmoid_f := 1;
        ELSIF x =- 15378 THEN
            sigmoid_f := 1;
        ELSIF x =- 15377 THEN
            sigmoid_f := 1;
        ELSIF x =- 15376 THEN
            sigmoid_f := 1;
        ELSIF x =- 15375 THEN
            sigmoid_f := 1;
        ELSIF x =- 15374 THEN
            sigmoid_f := 1;
        ELSIF x =- 15373 THEN
            sigmoid_f := 1;
        ELSIF x =- 15372 THEN
            sigmoid_f := 1;
        ELSIF x =- 15371 THEN
            sigmoid_f := 1;
        ELSIF x =- 15370 THEN
            sigmoid_f := 1;
        ELSIF x =- 15369 THEN
            sigmoid_f := 1;
        ELSIF x =- 15368 THEN
            sigmoid_f := 1;
        ELSIF x =- 15367 THEN
            sigmoid_f := 1;
        ELSIF x =- 15366 THEN
            sigmoid_f := 1;
        ELSIF x =- 15365 THEN
            sigmoid_f := 1;
        ELSIF x =- 15364 THEN
            sigmoid_f := 1;
        ELSIF x =- 15363 THEN
            sigmoid_f := 1;
        ELSIF x =- 15362 THEN
            sigmoid_f := 1;
        ELSIF x =- 15361 THEN
            sigmoid_f := 1;
        ELSIF x =- 15360 THEN
            sigmoid_f := 1;
        ELSIF x =- 15359 THEN
            sigmoid_f := 1;
        ELSIF x =- 15358 THEN
            sigmoid_f := 1;
        ELSIF x =- 15357 THEN
            sigmoid_f := 1;
        ELSIF x =- 15356 THEN
            sigmoid_f := 1;
        ELSIF x =- 15355 THEN
            sigmoid_f := 1;
        ELSIF x =- 15354 THEN
            sigmoid_f := 1;
        ELSIF x =- 15353 THEN
            sigmoid_f := 1;
        ELSIF x =- 15352 THEN
            sigmoid_f := 1;
        ELSIF x =- 15351 THEN
            sigmoid_f := 1;
        ELSIF x =- 15350 THEN
            sigmoid_f := 1;
        ELSIF x =- 15349 THEN
            sigmoid_f := 1;
        ELSIF x =- 15348 THEN
            sigmoid_f := 1;
        ELSIF x =- 15347 THEN
            sigmoid_f := 1;
        ELSIF x =- 15346 THEN
            sigmoid_f := 1;
        ELSIF x =- 15345 THEN
            sigmoid_f := 1;
        ELSIF x =- 15344 THEN
            sigmoid_f := 1;
        ELSIF x =- 15343 THEN
            sigmoid_f := 1;
        ELSIF x =- 15342 THEN
            sigmoid_f := 1;
        ELSIF x =- 15341 THEN
            sigmoid_f := 1;
        ELSIF x =- 15340 THEN
            sigmoid_f := 1;
        ELSIF x =- 15339 THEN
            sigmoid_f := 1;
        ELSIF x =- 15338 THEN
            sigmoid_f := 1;
        ELSIF x =- 15337 THEN
            sigmoid_f := 1;
        ELSIF x =- 15336 THEN
            sigmoid_f := 1;
        ELSIF x =- 15335 THEN
            sigmoid_f := 1;
        ELSIF x =- 15334 THEN
            sigmoid_f := 1;
        ELSIF x =- 15333 THEN
            sigmoid_f := 1;
        ELSIF x =- 15332 THEN
            sigmoid_f := 1;
        ELSIF x =- 15331 THEN
            sigmoid_f := 1;
        ELSIF x =- 15330 THEN
            sigmoid_f := 1;
        ELSIF x =- 15329 THEN
            sigmoid_f := 1;
        ELSIF x =- 15328 THEN
            sigmoid_f := 1;
        ELSIF x =- 15327 THEN
            sigmoid_f := 1;
        ELSIF x =- 15326 THEN
            sigmoid_f := 1;
        ELSIF x =- 15325 THEN
            sigmoid_f := 1;
        ELSIF x =- 15324 THEN
            sigmoid_f := 1;
        ELSIF x =- 15323 THEN
            sigmoid_f := 1;
        ELSIF x =- 15322 THEN
            sigmoid_f := 1;
        ELSIF x =- 15321 THEN
            sigmoid_f := 1;
        ELSIF x =- 15320 THEN
            sigmoid_f := 1;
        ELSIF x =- 15319 THEN
            sigmoid_f := 1;
        ELSIF x =- 15318 THEN
            sigmoid_f := 1;
        ELSIF x =- 15317 THEN
            sigmoid_f := 1;
        ELSIF x =- 15316 THEN
            sigmoid_f := 1;
        ELSIF x =- 15315 THEN
            sigmoid_f := 1;
        ELSIF x =- 15314 THEN
            sigmoid_f := 1;
        ELSIF x =- 15313 THEN
            sigmoid_f := 1;
        ELSIF x =- 15312 THEN
            sigmoid_f := 1;
        ELSIF x =- 15311 THEN
            sigmoid_f := 1;
        ELSIF x =- 15310 THEN
            sigmoid_f := 1;
        ELSIF x =- 15309 THEN
            sigmoid_f := 1;
        ELSIF x =- 15308 THEN
            sigmoid_f := 1;
        ELSIF x =- 15307 THEN
            sigmoid_f := 1;
        ELSIF x =- 15306 THEN
            sigmoid_f := 1;
        ELSIF x =- 15305 THEN
            sigmoid_f := 1;
        ELSIF x =- 15304 THEN
            sigmoid_f := 1;
        ELSIF x =- 15303 THEN
            sigmoid_f := 1;
        ELSIF x =- 15302 THEN
            sigmoid_f := 1;
        ELSIF x =- 15301 THEN
            sigmoid_f := 1;
        ELSIF x =- 15300 THEN
            sigmoid_f := 1;
        ELSIF x =- 15299 THEN
            sigmoid_f := 1;
        ELSIF x =- 15298 THEN
            sigmoid_f := 1;
        ELSIF x =- 15297 THEN
            sigmoid_f := 1;
        ELSIF x =- 15296 THEN
            sigmoid_f := 1;
        ELSIF x =- 15295 THEN
            sigmoid_f := 1;
        ELSIF x =- 15294 THEN
            sigmoid_f := 1;
        ELSIF x =- 15293 THEN
            sigmoid_f := 1;
        ELSIF x =- 15292 THEN
            sigmoid_f := 1;
        ELSIF x =- 15291 THEN
            sigmoid_f := 1;
        ELSIF x =- 15290 THEN
            sigmoid_f := 1;
        ELSIF x =- 15289 THEN
            sigmoid_f := 1;
        ELSIF x =- 15288 THEN
            sigmoid_f := 1;
        ELSIF x =- 15287 THEN
            sigmoid_f := 1;
        ELSIF x =- 15286 THEN
            sigmoid_f := 1;
        ELSIF x =- 15285 THEN
            sigmoid_f := 1;
        ELSIF x =- 15284 THEN
            sigmoid_f := 1;
        ELSIF x =- 15283 THEN
            sigmoid_f := 1;
        ELSIF x =- 15282 THEN
            sigmoid_f := 1;
        ELSIF x =- 15281 THEN
            sigmoid_f := 1;
        ELSIF x =- 15280 THEN
            sigmoid_f := 1;
        ELSIF x =- 15279 THEN
            sigmoid_f := 1;
        ELSIF x =- 15278 THEN
            sigmoid_f := 1;
        ELSIF x =- 15277 THEN
            sigmoid_f := 1;
        ELSIF x =- 15276 THEN
            sigmoid_f := 1;
        ELSIF x =- 15275 THEN
            sigmoid_f := 1;
        ELSIF x =- 15274 THEN
            sigmoid_f := 1;
        ELSIF x =- 15273 THEN
            sigmoid_f := 1;
        ELSIF x =- 15272 THEN
            sigmoid_f := 1;
        ELSIF x =- 15271 THEN
            sigmoid_f := 1;
        ELSIF x =- 15270 THEN
            sigmoid_f := 1;
        ELSIF x =- 15269 THEN
            sigmoid_f := 1;
        ELSIF x =- 15268 THEN
            sigmoid_f := 1;
        ELSIF x =- 15267 THEN
            sigmoid_f := 1;
        ELSIF x =- 15266 THEN
            sigmoid_f := 1;
        ELSIF x =- 15265 THEN
            sigmoid_f := 1;
        ELSIF x =- 15264 THEN
            sigmoid_f := 1;
        ELSIF x =- 15263 THEN
            sigmoid_f := 1;
        ELSIF x =- 15262 THEN
            sigmoid_f := 1;
        ELSIF x =- 15261 THEN
            sigmoid_f := 1;
        ELSIF x =- 15260 THEN
            sigmoid_f := 1;
        ELSIF x =- 15259 THEN
            sigmoid_f := 1;
        ELSIF x =- 15258 THEN
            sigmoid_f := 1;
        ELSIF x =- 15257 THEN
            sigmoid_f := 1;
        ELSIF x =- 15256 THEN
            sigmoid_f := 1;
        ELSIF x =- 15255 THEN
            sigmoid_f := 1;
        ELSIF x =- 15254 THEN
            sigmoid_f := 1;
        ELSIF x =- 15253 THEN
            sigmoid_f := 1;
        ELSIF x =- 15252 THEN
            sigmoid_f := 1;
        ELSIF x =- 15251 THEN
            sigmoid_f := 1;
        ELSIF x =- 15250 THEN
            sigmoid_f := 1;
        ELSIF x =- 15249 THEN
            sigmoid_f := 1;
        ELSIF x =- 15248 THEN
            sigmoid_f := 1;
        ELSIF x =- 15247 THEN
            sigmoid_f := 1;
        ELSIF x =- 15246 THEN
            sigmoid_f := 1;
        ELSIF x =- 15245 THEN
            sigmoid_f := 1;
        ELSIF x =- 15244 THEN
            sigmoid_f := 1;
        ELSIF x =- 15243 THEN
            sigmoid_f := 1;
        ELSIF x =- 15242 THEN
            sigmoid_f := 1;
        ELSIF x =- 15241 THEN
            sigmoid_f := 1;
        ELSIF x =- 15240 THEN
            sigmoid_f := 1;
        ELSIF x =- 15239 THEN
            sigmoid_f := 1;
        ELSIF x =- 15238 THEN
            sigmoid_f := 1;
        ELSIF x =- 15237 THEN
            sigmoid_f := 1;
        ELSIF x =- 15236 THEN
            sigmoid_f := 1;
        ELSIF x =- 15235 THEN
            sigmoid_f := 1;
        ELSIF x =- 15234 THEN
            sigmoid_f := 1;
        ELSIF x =- 15233 THEN
            sigmoid_f := 1;
        ELSIF x =- 15232 THEN
            sigmoid_f := 1;
        ELSIF x =- 15231 THEN
            sigmoid_f := 1;
        ELSIF x =- 15230 THEN
            sigmoid_f := 1;
        ELSIF x =- 15229 THEN
            sigmoid_f := 1;
        ELSIF x =- 15228 THEN
            sigmoid_f := 1;
        ELSIF x =- 15227 THEN
            sigmoid_f := 1;
        ELSIF x =- 15226 THEN
            sigmoid_f := 1;
        ELSIF x =- 15225 THEN
            sigmoid_f := 1;
        ELSIF x =- 15224 THEN
            sigmoid_f := 1;
        ELSIF x =- 15223 THEN
            sigmoid_f := 1;
        ELSIF x =- 15222 THEN
            sigmoid_f := 1;
        ELSIF x =- 15221 THEN
            sigmoid_f := 1;
        ELSIF x =- 15220 THEN
            sigmoid_f := 1;
        ELSIF x =- 15219 THEN
            sigmoid_f := 1;
        ELSIF x =- 15218 THEN
            sigmoid_f := 1;
        ELSIF x =- 15217 THEN
            sigmoid_f := 1;
        ELSIF x =- 15216 THEN
            sigmoid_f := 1;
        ELSIF x =- 15215 THEN
            sigmoid_f := 1;
        ELSIF x =- 15214 THEN
            sigmoid_f := 1;
        ELSIF x =- 15213 THEN
            sigmoid_f := 1;
        ELSIF x =- 15212 THEN
            sigmoid_f := 1;
        ELSIF x =- 15211 THEN
            sigmoid_f := 1;
        ELSIF x =- 15210 THEN
            sigmoid_f := 1;
        ELSIF x =- 15209 THEN
            sigmoid_f := 1;
        ELSIF x =- 15208 THEN
            sigmoid_f := 1;
        ELSIF x =- 15207 THEN
            sigmoid_f := 1;
        ELSIF x =- 15206 THEN
            sigmoid_f := 1;
        ELSIF x =- 15205 THEN
            sigmoid_f := 1;
        ELSIF x =- 15204 THEN
            sigmoid_f := 1;
        ELSIF x =- 15203 THEN
            sigmoid_f := 1;
        ELSIF x =- 15202 THEN
            sigmoid_f := 1;
        ELSIF x =- 15201 THEN
            sigmoid_f := 1;
        ELSIF x =- 15200 THEN
            sigmoid_f := 1;
        ELSIF x =- 15199 THEN
            sigmoid_f := 1;
        ELSIF x =- 15198 THEN
            sigmoid_f := 1;
        ELSIF x =- 15197 THEN
            sigmoid_f := 1;
        ELSIF x =- 15196 THEN
            sigmoid_f := 1;
        ELSIF x =- 15195 THEN
            sigmoid_f := 1;
        ELSIF x =- 15194 THEN
            sigmoid_f := 1;
        ELSIF x =- 15193 THEN
            sigmoid_f := 1;
        ELSIF x =- 15192 THEN
            sigmoid_f := 1;
        ELSIF x =- 15191 THEN
            sigmoid_f := 1;
        ELSIF x =- 15190 THEN
            sigmoid_f := 1;
        ELSIF x =- 15189 THEN
            sigmoid_f := 1;
        ELSIF x =- 15188 THEN
            sigmoid_f := 1;
        ELSIF x =- 15187 THEN
            sigmoid_f := 1;
        ELSIF x =- 15186 THEN
            sigmoid_f := 1;
        ELSIF x =- 15185 THEN
            sigmoid_f := 1;
        ELSIF x =- 15184 THEN
            sigmoid_f := 1;
        ELSIF x =- 15183 THEN
            sigmoid_f := 1;
        ELSIF x =- 15182 THEN
            sigmoid_f := 1;
        ELSIF x =- 15181 THEN
            sigmoid_f := 1;
        ELSIF x =- 15180 THEN
            sigmoid_f := 1;
        ELSIF x =- 15179 THEN
            sigmoid_f := 1;
        ELSIF x =- 15178 THEN
            sigmoid_f := 1;
        ELSIF x =- 15177 THEN
            sigmoid_f := 1;
        ELSIF x =- 15176 THEN
            sigmoid_f := 1;
        ELSIF x =- 15175 THEN
            sigmoid_f := 1;
        ELSIF x =- 15174 THEN
            sigmoid_f := 1;
        ELSIF x =- 15173 THEN
            sigmoid_f := 1;
        ELSIF x =- 15172 THEN
            sigmoid_f := 1;
        ELSIF x =- 15171 THEN
            sigmoid_f := 1;
        ELSIF x =- 15170 THEN
            sigmoid_f := 1;
        ELSIF x =- 15169 THEN
            sigmoid_f := 1;
        ELSIF x =- 15168 THEN
            sigmoid_f := 1;
        ELSIF x =- 15167 THEN
            sigmoid_f := 1;
        ELSIF x =- 15166 THEN
            sigmoid_f := 1;
        ELSIF x =- 15165 THEN
            sigmoid_f := 1;
        ELSIF x =- 15164 THEN
            sigmoid_f := 1;
        ELSIF x =- 15163 THEN
            sigmoid_f := 1;
        ELSIF x =- 15162 THEN
            sigmoid_f := 1;
        ELSIF x =- 15161 THEN
            sigmoid_f := 1;
        ELSIF x =- 15160 THEN
            sigmoid_f := 1;
        ELSIF x =- 15159 THEN
            sigmoid_f := 1;
        ELSIF x =- 15158 THEN
            sigmoid_f := 1;
        ELSIF x =- 15157 THEN
            sigmoid_f := 1;
        ELSIF x =- 15156 THEN
            sigmoid_f := 1;
        ELSIF x =- 15155 THEN
            sigmoid_f := 1;
        ELSIF x =- 15154 THEN
            sigmoid_f := 1;
        ELSIF x =- 15153 THEN
            sigmoid_f := 1;
        ELSIF x =- 15152 THEN
            sigmoid_f := 1;
        ELSIF x =- 15151 THEN
            sigmoid_f := 1;
        ELSIF x =- 15150 THEN
            sigmoid_f := 1;
        ELSIF x =- 15149 THEN
            sigmoid_f := 1;
        ELSIF x =- 15148 THEN
            sigmoid_f := 1;
        ELSIF x =- 15147 THEN
            sigmoid_f := 1;
        ELSIF x =- 15146 THEN
            sigmoid_f := 1;
        ELSIF x =- 15145 THEN
            sigmoid_f := 1;
        ELSIF x =- 15144 THEN
            sigmoid_f := 1;
        ELSIF x =- 15143 THEN
            sigmoid_f := 1;
        ELSIF x =- 15142 THEN
            sigmoid_f := 1;
        ELSIF x =- 15141 THEN
            sigmoid_f := 1;
        ELSIF x =- 15140 THEN
            sigmoid_f := 1;
        ELSIF x =- 15139 THEN
            sigmoid_f := 1;
        ELSIF x =- 15138 THEN
            sigmoid_f := 1;
        ELSIF x =- 15137 THEN
            sigmoid_f := 1;
        ELSIF x =- 15136 THEN
            sigmoid_f := 1;
        ELSIF x =- 15135 THEN
            sigmoid_f := 1;
        ELSIF x =- 15134 THEN
            sigmoid_f := 1;
        ELSIF x =- 15133 THEN
            sigmoid_f := 1;
        ELSIF x =- 15132 THEN
            sigmoid_f := 1;
        ELSIF x =- 15131 THEN
            sigmoid_f := 1;
        ELSIF x =- 15130 THEN
            sigmoid_f := 1;
        ELSIF x =- 15129 THEN
            sigmoid_f := 1;
        ELSIF x =- 15128 THEN
            sigmoid_f := 1;
        ELSIF x =- 15127 THEN
            sigmoid_f := 1;
        ELSIF x =- 15126 THEN
            sigmoid_f := 1;
        ELSIF x =- 15125 THEN
            sigmoid_f := 1;
        ELSIF x =- 15124 THEN
            sigmoid_f := 1;
        ELSIF x =- 15123 THEN
            sigmoid_f := 1;
        ELSIF x =- 15122 THEN
            sigmoid_f := 1;
        ELSIF x =- 15121 THEN
            sigmoid_f := 1;
        ELSIF x =- 15120 THEN
            sigmoid_f := 1;
        ELSIF x =- 15119 THEN
            sigmoid_f := 1;
        ELSIF x =- 15118 THEN
            sigmoid_f := 1;
        ELSIF x =- 15117 THEN
            sigmoid_f := 1;
        ELSIF x =- 15116 THEN
            sigmoid_f := 1;
        ELSIF x =- 15115 THEN
            sigmoid_f := 1;
        ELSIF x =- 15114 THEN
            sigmoid_f := 1;
        ELSIF x =- 15113 THEN
            sigmoid_f := 1;
        ELSIF x =- 15112 THEN
            sigmoid_f := 1;
        ELSIF x =- 15111 THEN
            sigmoid_f := 1;
        ELSIF x =- 15110 THEN
            sigmoid_f := 1;
        ELSIF x =- 15109 THEN
            sigmoid_f := 1;
        ELSIF x =- 15108 THEN
            sigmoid_f := 1;
        ELSIF x =- 15107 THEN
            sigmoid_f := 1;
        ELSIF x =- 15106 THEN
            sigmoid_f := 1;
        ELSIF x =- 15105 THEN
            sigmoid_f := 1;
        ELSIF x =- 15104 THEN
            sigmoid_f := 1;
        ELSIF x =- 15103 THEN
            sigmoid_f := 1;
        ELSIF x =- 15102 THEN
            sigmoid_f := 1;
        ELSIF x =- 15101 THEN
            sigmoid_f := 1;
        ELSIF x =- 15100 THEN
            sigmoid_f := 1;
        ELSIF x =- 15099 THEN
            sigmoid_f := 1;
        ELSIF x =- 15098 THEN
            sigmoid_f := 1;
        ELSIF x =- 15097 THEN
            sigmoid_f := 1;
        ELSIF x =- 15096 THEN
            sigmoid_f := 1;
        ELSIF x =- 15095 THEN
            sigmoid_f := 1;
        ELSIF x =- 15094 THEN
            sigmoid_f := 1;
        ELSIF x =- 15093 THEN
            sigmoid_f := 1;
        ELSIF x =- 15092 THEN
            sigmoid_f := 1;
        ELSIF x =- 15091 THEN
            sigmoid_f := 1;
        ELSIF x =- 15090 THEN
            sigmoid_f := 1;
        ELSIF x =- 15089 THEN
            sigmoid_f := 1;
        ELSIF x =- 15088 THEN
            sigmoid_f := 1;
        ELSIF x =- 15087 THEN
            sigmoid_f := 1;
        ELSIF x =- 15086 THEN
            sigmoid_f := 1;
        ELSIF x =- 15085 THEN
            sigmoid_f := 1;
        ELSIF x =- 15084 THEN
            sigmoid_f := 1;
        ELSIF x =- 15083 THEN
            sigmoid_f := 1;
        ELSIF x =- 15082 THEN
            sigmoid_f := 1;
        ELSIF x =- 15081 THEN
            sigmoid_f := 1;
        ELSIF x =- 15080 THEN
            sigmoid_f := 1;
        ELSIF x =- 15079 THEN
            sigmoid_f := 1;
        ELSIF x =- 15078 THEN
            sigmoid_f := 1;
        ELSIF x =- 15077 THEN
            sigmoid_f := 1;
        ELSIF x =- 15076 THEN
            sigmoid_f := 1;
        ELSIF x =- 15075 THEN
            sigmoid_f := 1;
        ELSIF x =- 15074 THEN
            sigmoid_f := 1;
        ELSIF x =- 15073 THEN
            sigmoid_f := 1;
        ELSIF x =- 15072 THEN
            sigmoid_f := 1;
        ELSIF x =- 15071 THEN
            sigmoid_f := 1;
        ELSIF x =- 15070 THEN
            sigmoid_f := 1;
        ELSIF x =- 15069 THEN
            sigmoid_f := 1;
        ELSIF x =- 15068 THEN
            sigmoid_f := 1;
        ELSIF x =- 15067 THEN
            sigmoid_f := 1;
        ELSIF x =- 15066 THEN
            sigmoid_f := 1;
        ELSIF x =- 15065 THEN
            sigmoid_f := 1;
        ELSIF x =- 15064 THEN
            sigmoid_f := 1;
        ELSIF x =- 15063 THEN
            sigmoid_f := 1;
        ELSIF x =- 15062 THEN
            sigmoid_f := 1;
        ELSIF x =- 15061 THEN
            sigmoid_f := 1;
        ELSIF x =- 15060 THEN
            sigmoid_f := 1;
        ELSIF x =- 15059 THEN
            sigmoid_f := 1;
        ELSIF x =- 15058 THEN
            sigmoid_f := 1;
        ELSIF x =- 15057 THEN
            sigmoid_f := 1;
        ELSIF x =- 15056 THEN
            sigmoid_f := 1;
        ELSIF x =- 15055 THEN
            sigmoid_f := 1;
        ELSIF x =- 15054 THEN
            sigmoid_f := 1;
        ELSIF x =- 15053 THEN
            sigmoid_f := 1;
        ELSIF x =- 15052 THEN
            sigmoid_f := 1;
        ELSIF x =- 15051 THEN
            sigmoid_f := 1;
        ELSIF x =- 15050 THEN
            sigmoid_f := 1;
        ELSIF x =- 15049 THEN
            sigmoid_f := 1;
        ELSIF x =- 15048 THEN
            sigmoid_f := 1;
        ELSIF x =- 15047 THEN
            sigmoid_f := 1;
        ELSIF x =- 15046 THEN
            sigmoid_f := 1;
        ELSIF x =- 15045 THEN
            sigmoid_f := 1;
        ELSIF x =- 15044 THEN
            sigmoid_f := 1;
        ELSIF x =- 15043 THEN
            sigmoid_f := 1;
        ELSIF x =- 15042 THEN
            sigmoid_f := 1;
        ELSIF x =- 15041 THEN
            sigmoid_f := 1;
        ELSIF x =- 15040 THEN
            sigmoid_f := 1;
        ELSIF x =- 15039 THEN
            sigmoid_f := 1;
        ELSIF x =- 15038 THEN
            sigmoid_f := 1;
        ELSIF x =- 15037 THEN
            sigmoid_f := 1;
        ELSIF x =- 15036 THEN
            sigmoid_f := 1;
        ELSIF x =- 15035 THEN
            sigmoid_f := 1;
        ELSIF x =- 15034 THEN
            sigmoid_f := 1;
        ELSIF x =- 15033 THEN
            sigmoid_f := 1;
        ELSIF x =- 15032 THEN
            sigmoid_f := 1;
        ELSIF x =- 15031 THEN
            sigmoid_f := 1;
        ELSIF x =- 15030 THEN
            sigmoid_f := 1;
        ELSIF x =- 15029 THEN
            sigmoid_f := 1;
        ELSIF x =- 15028 THEN
            sigmoid_f := 1;
        ELSIF x =- 15027 THEN
            sigmoid_f := 1;
        ELSIF x =- 15026 THEN
            sigmoid_f := 1;
        ELSIF x =- 15025 THEN
            sigmoid_f := 1;
        ELSIF x =- 15024 THEN
            sigmoid_f := 1;
        ELSIF x =- 15023 THEN
            sigmoid_f := 1;
        ELSIF x =- 15022 THEN
            sigmoid_f := 1;
        ELSIF x =- 15021 THEN
            sigmoid_f := 1;
        ELSIF x =- 15020 THEN
            sigmoid_f := 1;
        ELSIF x =- 15019 THEN
            sigmoid_f := 1;
        ELSIF x =- 15018 THEN
            sigmoid_f := 1;
        ELSIF x =- 15017 THEN
            sigmoid_f := 1;
        ELSIF x =- 15016 THEN
            sigmoid_f := 1;
        ELSIF x =- 15015 THEN
            sigmoid_f := 1;
        ELSIF x =- 15014 THEN
            sigmoid_f := 1;
        ELSIF x =- 15013 THEN
            sigmoid_f := 1;
        ELSIF x =- 15012 THEN
            sigmoid_f := 1;
        ELSIF x =- 15011 THEN
            sigmoid_f := 1;
        ELSIF x =- 15010 THEN
            sigmoid_f := 1;
        ELSIF x =- 15009 THEN
            sigmoid_f := 1;
        ELSIF x =- 15008 THEN
            sigmoid_f := 1;
        ELSIF x =- 15007 THEN
            sigmoid_f := 1;
        ELSIF x =- 15006 THEN
            sigmoid_f := 1;
        ELSIF x =- 15005 THEN
            sigmoid_f := 1;
        ELSIF x =- 15004 THEN
            sigmoid_f := 1;
        ELSIF x =- 15003 THEN
            sigmoid_f := 1;
        ELSIF x =- 15002 THEN
            sigmoid_f := 1;
        ELSIF x =- 15001 THEN
            sigmoid_f := 1;
        ELSIF x =- 15000 THEN
            sigmoid_f := 1;
        ELSIF x =- 14999 THEN
            sigmoid_f := 1;
        ELSIF x =- 14998 THEN
            sigmoid_f := 1;
        ELSIF x =- 14997 THEN
            sigmoid_f := 1;
        ELSIF x =- 14996 THEN
            sigmoid_f := 1;
        ELSIF x =- 14995 THEN
            sigmoid_f := 1;
        ELSIF x =- 14994 THEN
            sigmoid_f := 1;
        ELSIF x =- 14993 THEN
            sigmoid_f := 1;
        ELSIF x =- 14992 THEN
            sigmoid_f := 1;
        ELSIF x =- 14991 THEN
            sigmoid_f := 1;
        ELSIF x =- 14990 THEN
            sigmoid_f := 1;
        ELSIF x =- 14989 THEN
            sigmoid_f := 1;
        ELSIF x =- 14988 THEN
            sigmoid_f := 1;
        ELSIF x =- 14987 THEN
            sigmoid_f := 1;
        ELSIF x =- 14986 THEN
            sigmoid_f := 1;
        ELSIF x =- 14985 THEN
            sigmoid_f := 1;
        ELSIF x =- 14984 THEN
            sigmoid_f := 1;
        ELSIF x =- 14983 THEN
            sigmoid_f := 1;
        ELSIF x =- 14982 THEN
            sigmoid_f := 1;
        ELSIF x =- 14981 THEN
            sigmoid_f := 1;
        ELSIF x =- 14980 THEN
            sigmoid_f := 1;
        ELSIF x =- 14979 THEN
            sigmoid_f := 1;
        ELSIF x =- 14978 THEN
            sigmoid_f := 1;
        ELSIF x =- 14977 THEN
            sigmoid_f := 1;
        ELSIF x =- 14976 THEN
            sigmoid_f := 1;
        ELSIF x =- 14975 THEN
            sigmoid_f := 1;
        ELSIF x =- 14974 THEN
            sigmoid_f := 1;
        ELSIF x =- 14973 THEN
            sigmoid_f := 1;
        ELSIF x =- 14972 THEN
            sigmoid_f := 1;
        ELSIF x =- 14971 THEN
            sigmoid_f := 1;
        ELSIF x =- 14970 THEN
            sigmoid_f := 1;
        ELSIF x =- 14969 THEN
            sigmoid_f := 1;
        ELSIF x =- 14968 THEN
            sigmoid_f := 1;
        ELSIF x =- 14967 THEN
            sigmoid_f := 1;
        ELSIF x =- 14966 THEN
            sigmoid_f := 1;
        ELSIF x =- 14965 THEN
            sigmoid_f := 1;
        ELSIF x =- 14964 THEN
            sigmoid_f := 1;
        ELSIF x =- 14963 THEN
            sigmoid_f := 1;
        ELSIF x =- 14962 THEN
            sigmoid_f := 1;
        ELSIF x =- 14961 THEN
            sigmoid_f := 1;
        ELSIF x =- 14960 THEN
            sigmoid_f := 1;
        ELSIF x =- 14959 THEN
            sigmoid_f := 1;
        ELSIF x =- 14958 THEN
            sigmoid_f := 1;
        ELSIF x =- 14957 THEN
            sigmoid_f := 1;
        ELSIF x =- 14956 THEN
            sigmoid_f := 1;
        ELSIF x =- 14955 THEN
            sigmoid_f := 1;
        ELSIF x =- 14954 THEN
            sigmoid_f := 1;
        ELSIF x =- 14953 THEN
            sigmoid_f := 1;
        ELSIF x =- 14952 THEN
            sigmoid_f := 1;
        ELSIF x =- 14951 THEN
            sigmoid_f := 1;
        ELSIF x =- 14950 THEN
            sigmoid_f := 1;
        ELSIF x =- 14949 THEN
            sigmoid_f := 1;
        ELSIF x =- 14948 THEN
            sigmoid_f := 1;
        ELSIF x =- 14947 THEN
            sigmoid_f := 1;
        ELSIF x =- 14946 THEN
            sigmoid_f := 1;
        ELSIF x =- 14945 THEN
            sigmoid_f := 1;
        ELSIF x =- 14944 THEN
            sigmoid_f := 1;
        ELSIF x =- 14943 THEN
            sigmoid_f := 1;
        ELSIF x =- 14942 THEN
            sigmoid_f := 1;
        ELSIF x =- 14941 THEN
            sigmoid_f := 1;
        ELSIF x =- 14940 THEN
            sigmoid_f := 1;
        ELSIF x =- 14939 THEN
            sigmoid_f := 1;
        ELSIF x =- 14938 THEN
            sigmoid_f := 1;
        ELSIF x =- 14937 THEN
            sigmoid_f := 1;
        ELSIF x =- 14936 THEN
            sigmoid_f := 1;
        ELSIF x =- 14935 THEN
            sigmoid_f := 1;
        ELSIF x =- 14934 THEN
            sigmoid_f := 1;
        ELSIF x =- 14933 THEN
            sigmoid_f := 1;
        ELSIF x =- 14932 THEN
            sigmoid_f := 1;
        ELSIF x =- 14931 THEN
            sigmoid_f := 1;
        ELSIF x =- 14930 THEN
            sigmoid_f := 1;
        ELSIF x =- 14929 THEN
            sigmoid_f := 1;
        ELSIF x =- 14928 THEN
            sigmoid_f := 1;
        ELSIF x =- 14927 THEN
            sigmoid_f := 1;
        ELSIF x =- 14926 THEN
            sigmoid_f := 1;
        ELSIF x =- 14925 THEN
            sigmoid_f := 1;
        ELSIF x =- 14924 THEN
            sigmoid_f := 1;
        ELSIF x =- 14923 THEN
            sigmoid_f := 1;
        ELSIF x =- 14922 THEN
            sigmoid_f := 1;
        ELSIF x =- 14921 THEN
            sigmoid_f := 1;
        ELSIF x =- 14920 THEN
            sigmoid_f := 1;
        ELSIF x =- 14919 THEN
            sigmoid_f := 1;
        ELSIF x =- 14918 THEN
            sigmoid_f := 1;
        ELSIF x =- 14917 THEN
            sigmoid_f := 1;
        ELSIF x =- 14916 THEN
            sigmoid_f := 1;
        ELSIF x =- 14915 THEN
            sigmoid_f := 1;
        ELSIF x =- 14914 THEN
            sigmoid_f := 1;
        ELSIF x =- 14913 THEN
            sigmoid_f := 1;
        ELSIF x =- 14912 THEN
            sigmoid_f := 1;
        ELSIF x =- 14911 THEN
            sigmoid_f := 1;
        ELSIF x =- 14910 THEN
            sigmoid_f := 1;
        ELSIF x =- 14909 THEN
            sigmoid_f := 1;
        ELSIF x =- 14908 THEN
            sigmoid_f := 1;
        ELSIF x =- 14907 THEN
            sigmoid_f := 1;
        ELSIF x =- 14906 THEN
            sigmoid_f := 1;
        ELSIF x =- 14905 THEN
            sigmoid_f := 1;
        ELSIF x =- 14904 THEN
            sigmoid_f := 1;
        ELSIF x =- 14903 THEN
            sigmoid_f := 1;
        ELSIF x =- 14902 THEN
            sigmoid_f := 1;
        ELSIF x =- 14901 THEN
            sigmoid_f := 1;
        ELSIF x =- 14900 THEN
            sigmoid_f := 1;
        ELSIF x =- 14899 THEN
            sigmoid_f := 1;
        ELSIF x =- 14898 THEN
            sigmoid_f := 1;
        ELSIF x =- 14897 THEN
            sigmoid_f := 1;
        ELSIF x =- 14896 THEN
            sigmoid_f := 1;
        ELSIF x =- 14895 THEN
            sigmoid_f := 1;
        ELSIF x =- 14894 THEN
            sigmoid_f := 1;
        ELSIF x =- 14893 THEN
            sigmoid_f := 1;
        ELSIF x =- 14892 THEN
            sigmoid_f := 1;
        ELSIF x =- 14891 THEN
            sigmoid_f := 1;
        ELSIF x =- 14890 THEN
            sigmoid_f := 1;
        ELSIF x =- 14889 THEN
            sigmoid_f := 1;
        ELSIF x =- 14888 THEN
            sigmoid_f := 1;
        ELSIF x =- 14887 THEN
            sigmoid_f := 1;
        ELSIF x =- 14886 THEN
            sigmoid_f := 1;
        ELSIF x =- 14885 THEN
            sigmoid_f := 1;
        ELSIF x =- 14884 THEN
            sigmoid_f := 1;
        ELSIF x =- 14883 THEN
            sigmoid_f := 1;
        ELSIF x =- 14882 THEN
            sigmoid_f := 1;
        ELSIF x =- 14881 THEN
            sigmoid_f := 1;
        ELSIF x =- 14880 THEN
            sigmoid_f := 1;
        ELSIF x =- 14879 THEN
            sigmoid_f := 1;
        ELSIF x =- 14878 THEN
            sigmoid_f := 1;
        ELSIF x =- 14877 THEN
            sigmoid_f := 1;
        ELSIF x =- 14876 THEN
            sigmoid_f := 1;
        ELSIF x =- 14875 THEN
            sigmoid_f := 1;
        ELSIF x =- 14874 THEN
            sigmoid_f := 1;
        ELSIF x =- 14873 THEN
            sigmoid_f := 1;
        ELSIF x =- 14872 THEN
            sigmoid_f := 1;
        ELSIF x =- 14871 THEN
            sigmoid_f := 1;
        ELSIF x =- 14870 THEN
            sigmoid_f := 1;
        ELSIF x =- 14869 THEN
            sigmoid_f := 1;
        ELSIF x =- 14868 THEN
            sigmoid_f := 1;
        ELSIF x =- 14867 THEN
            sigmoid_f := 1;
        ELSIF x =- 14866 THEN
            sigmoid_f := 1;
        ELSIF x =- 14865 THEN
            sigmoid_f := 1;
        ELSIF x =- 14864 THEN
            sigmoid_f := 1;
        ELSIF x =- 14863 THEN
            sigmoid_f := 1;
        ELSIF x =- 14862 THEN
            sigmoid_f := 1;
        ELSIF x =- 14861 THEN
            sigmoid_f := 1;
        ELSIF x =- 14860 THEN
            sigmoid_f := 1;
        ELSIF x =- 14859 THEN
            sigmoid_f := 1;
        ELSIF x =- 14858 THEN
            sigmoid_f := 1;
        ELSIF x =- 14857 THEN
            sigmoid_f := 1;
        ELSIF x =- 14856 THEN
            sigmoid_f := 1;
        ELSIF x =- 14855 THEN
            sigmoid_f := 1;
        ELSIF x =- 14854 THEN
            sigmoid_f := 1;
        ELSIF x =- 14853 THEN
            sigmoid_f := 1;
        ELSIF x =- 14852 THEN
            sigmoid_f := 1;
        ELSIF x =- 14851 THEN
            sigmoid_f := 1;
        ELSIF x =- 14850 THEN
            sigmoid_f := 1;
        ELSIF x =- 14849 THEN
            sigmoid_f := 1;
        ELSIF x =- 14848 THEN
            sigmoid_f := 1;
        ELSIF x =- 14847 THEN
            sigmoid_f := 2;
        ELSIF x =- 14846 THEN
            sigmoid_f := 2;
        ELSIF x =- 14845 THEN
            sigmoid_f := 2;
        ELSIF x =- 14844 THEN
            sigmoid_f := 2;
        ELSIF x =- 14843 THEN
            sigmoid_f := 2;
        ELSIF x =- 14842 THEN
            sigmoid_f := 2;
        ELSIF x =- 14841 THEN
            sigmoid_f := 2;
        ELSIF x =- 14840 THEN
            sigmoid_f := 2;
        ELSIF x =- 14839 THEN
            sigmoid_f := 2;
        ELSIF x =- 14838 THEN
            sigmoid_f := 2;
        ELSIF x =- 14837 THEN
            sigmoid_f := 2;
        ELSIF x =- 14836 THEN
            sigmoid_f := 2;
        ELSIF x =- 14835 THEN
            sigmoid_f := 2;
        ELSIF x =- 14834 THEN
            sigmoid_f := 2;
        ELSIF x =- 14833 THEN
            sigmoid_f := 2;
        ELSIF x =- 14832 THEN
            sigmoid_f := 2;
        ELSIF x =- 14831 THEN
            sigmoid_f := 2;
        ELSIF x =- 14830 THEN
            sigmoid_f := 2;
        ELSIF x =- 14829 THEN
            sigmoid_f := 2;
        ELSIF x =- 14828 THEN
            sigmoid_f := 2;
        ELSIF x =- 14827 THEN
            sigmoid_f := 2;
        ELSIF x =- 14826 THEN
            sigmoid_f := 2;
        ELSIF x =- 14825 THEN
            sigmoid_f := 2;
        ELSIF x =- 14824 THEN
            sigmoid_f := 2;
        ELSIF x =- 14823 THEN
            sigmoid_f := 2;
        ELSIF x =- 14822 THEN
            sigmoid_f := 2;
        ELSIF x =- 14821 THEN
            sigmoid_f := 2;
        ELSIF x =- 14820 THEN
            sigmoid_f := 2;
        ELSIF x =- 14819 THEN
            sigmoid_f := 2;
        ELSIF x =- 14818 THEN
            sigmoid_f := 2;
        ELSIF x =- 14817 THEN
            sigmoid_f := 2;
        ELSIF x =- 14816 THEN
            sigmoid_f := 2;
        ELSIF x =- 14815 THEN
            sigmoid_f := 2;
        ELSIF x =- 14814 THEN
            sigmoid_f := 2;
        ELSIF x =- 14813 THEN
            sigmoid_f := 2;
        ELSIF x =- 14812 THEN
            sigmoid_f := 2;
        ELSIF x =- 14811 THEN
            sigmoid_f := 2;
        ELSIF x =- 14810 THEN
            sigmoid_f := 2;
        ELSIF x =- 14809 THEN
            sigmoid_f := 2;
        ELSIF x =- 14808 THEN
            sigmoid_f := 2;
        ELSIF x =- 14807 THEN
            sigmoid_f := 2;
        ELSIF x =- 14806 THEN
            sigmoid_f := 2;
        ELSIF x =- 14805 THEN
            sigmoid_f := 2;
        ELSIF x =- 14804 THEN
            sigmoid_f := 2;
        ELSIF x =- 14803 THEN
            sigmoid_f := 2;
        ELSIF x =- 14802 THEN
            sigmoid_f := 2;
        ELSIF x =- 14801 THEN
            sigmoid_f := 2;
        ELSIF x =- 14800 THEN
            sigmoid_f := 2;
        ELSIF x =- 14799 THEN
            sigmoid_f := 2;
        ELSIF x =- 14798 THEN
            sigmoid_f := 2;
        ELSIF x =- 14797 THEN
            sigmoid_f := 2;
        ELSIF x =- 14796 THEN
            sigmoid_f := 2;
        ELSIF x =- 14795 THEN
            sigmoid_f := 2;
        ELSIF x =- 14794 THEN
            sigmoid_f := 2;
        ELSIF x =- 14793 THEN
            sigmoid_f := 2;
        ELSIF x =- 14792 THEN
            sigmoid_f := 2;
        ELSIF x =- 14791 THEN
            sigmoid_f := 2;
        ELSIF x =- 14790 THEN
            sigmoid_f := 2;
        ELSIF x =- 14789 THEN
            sigmoid_f := 2;
        ELSIF x =- 14788 THEN
            sigmoid_f := 2;
        ELSIF x =- 14787 THEN
            sigmoid_f := 2;
        ELSIF x =- 14786 THEN
            sigmoid_f := 2;
        ELSIF x =- 14785 THEN
            sigmoid_f := 2;
        ELSIF x =- 14784 THEN
            sigmoid_f := 2;
        ELSIF x =- 14783 THEN
            sigmoid_f := 2;
        ELSIF x =- 14782 THEN
            sigmoid_f := 2;
        ELSIF x =- 14781 THEN
            sigmoid_f := 2;
        ELSIF x =- 14780 THEN
            sigmoid_f := 2;
        ELSIF x =- 14779 THEN
            sigmoid_f := 2;
        ELSIF x =- 14778 THEN
            sigmoid_f := 2;
        ELSIF x =- 14777 THEN
            sigmoid_f := 2;
        ELSIF x =- 14776 THEN
            sigmoid_f := 2;
        ELSIF x =- 14775 THEN
            sigmoid_f := 2;
        ELSIF x =- 14774 THEN
            sigmoid_f := 2;
        ELSIF x =- 14773 THEN
            sigmoid_f := 2;
        ELSIF x =- 14772 THEN
            sigmoid_f := 2;
        ELSIF x =- 14771 THEN
            sigmoid_f := 2;
        ELSIF x =- 14770 THEN
            sigmoid_f := 2;
        ELSIF x =- 14769 THEN
            sigmoid_f := 2;
        ELSIF x =- 14768 THEN
            sigmoid_f := 2;
        ELSIF x =- 14767 THEN
            sigmoid_f := 2;
        ELSIF x =- 14766 THEN
            sigmoid_f := 2;
        ELSIF x =- 14765 THEN
            sigmoid_f := 2;
        ELSIF x =- 14764 THEN
            sigmoid_f := 2;
        ELSIF x =- 14763 THEN
            sigmoid_f := 2;
        ELSIF x =- 14762 THEN
            sigmoid_f := 2;
        ELSIF x =- 14761 THEN
            sigmoid_f := 2;
        ELSIF x =- 14760 THEN
            sigmoid_f := 2;
        ELSIF x =- 14759 THEN
            sigmoid_f := 2;
        ELSIF x =- 14758 THEN
            sigmoid_f := 2;
        ELSIF x =- 14757 THEN
            sigmoid_f := 2;
        ELSIF x =- 14756 THEN
            sigmoid_f := 2;
        ELSIF x =- 14755 THEN
            sigmoid_f := 2;
        ELSIF x =- 14754 THEN
            sigmoid_f := 2;
        ELSIF x =- 14753 THEN
            sigmoid_f := 2;
        ELSIF x =- 14752 THEN
            sigmoid_f := 2;
        ELSIF x =- 14751 THEN
            sigmoid_f := 2;
        ELSIF x =- 14750 THEN
            sigmoid_f := 2;
        ELSIF x =- 14749 THEN
            sigmoid_f := 2;
        ELSIF x =- 14748 THEN
            sigmoid_f := 2;
        ELSIF x =- 14747 THEN
            sigmoid_f := 2;
        ELSIF x =- 14746 THEN
            sigmoid_f := 2;
        ELSIF x =- 14745 THEN
            sigmoid_f := 2;
        ELSIF x =- 14744 THEN
            sigmoid_f := 2;
        ELSIF x =- 14743 THEN
            sigmoid_f := 2;
        ELSIF x =- 14742 THEN
            sigmoid_f := 2;
        ELSIF x =- 14741 THEN
            sigmoid_f := 2;
        ELSIF x =- 14740 THEN
            sigmoid_f := 2;
        ELSIF x =- 14739 THEN
            sigmoid_f := 2;
        ELSIF x =- 14738 THEN
            sigmoid_f := 2;
        ELSIF x =- 14737 THEN
            sigmoid_f := 2;
        ELSIF x =- 14736 THEN
            sigmoid_f := 2;
        ELSIF x =- 14735 THEN
            sigmoid_f := 2;
        ELSIF x =- 14734 THEN
            sigmoid_f := 2;
        ELSIF x =- 14733 THEN
            sigmoid_f := 2;
        ELSIF x =- 14732 THEN
            sigmoid_f := 2;
        ELSIF x =- 14731 THEN
            sigmoid_f := 2;
        ELSIF x =- 14730 THEN
            sigmoid_f := 2;
        ELSIF x =- 14729 THEN
            sigmoid_f := 2;
        ELSIF x =- 14728 THEN
            sigmoid_f := 2;
        ELSIF x =- 14727 THEN
            sigmoid_f := 2;
        ELSIF x =- 14726 THEN
            sigmoid_f := 2;
        ELSIF x =- 14725 THEN
            sigmoid_f := 2;
        ELSIF x =- 14724 THEN
            sigmoid_f := 2;
        ELSIF x =- 14723 THEN
            sigmoid_f := 2;
        ELSIF x =- 14722 THEN
            sigmoid_f := 2;
        ELSIF x =- 14721 THEN
            sigmoid_f := 2;
        ELSIF x =- 14720 THEN
            sigmoid_f := 2;
        ELSIF x =- 14719 THEN
            sigmoid_f := 2;
        ELSIF x =- 14718 THEN
            sigmoid_f := 2;
        ELSIF x =- 14717 THEN
            sigmoid_f := 2;
        ELSIF x =- 14716 THEN
            sigmoid_f := 2;
        ELSIF x =- 14715 THEN
            sigmoid_f := 2;
        ELSIF x =- 14714 THEN
            sigmoid_f := 2;
        ELSIF x =- 14713 THEN
            sigmoid_f := 2;
        ELSIF x =- 14712 THEN
            sigmoid_f := 2;
        ELSIF x =- 14711 THEN
            sigmoid_f := 2;
        ELSIF x =- 14710 THEN
            sigmoid_f := 2;
        ELSIF x =- 14709 THEN
            sigmoid_f := 2;
        ELSIF x =- 14708 THEN
            sigmoid_f := 2;
        ELSIF x =- 14707 THEN
            sigmoid_f := 2;
        ELSIF x =- 14706 THEN
            sigmoid_f := 2;
        ELSIF x =- 14705 THEN
            sigmoid_f := 2;
        ELSIF x =- 14704 THEN
            sigmoid_f := 2;
        ELSIF x =- 14703 THEN
            sigmoid_f := 2;
        ELSIF x =- 14702 THEN
            sigmoid_f := 2;
        ELSIF x =- 14701 THEN
            sigmoid_f := 2;
        ELSIF x =- 14700 THEN
            sigmoid_f := 2;
        ELSIF x =- 14699 THEN
            sigmoid_f := 2;
        ELSIF x =- 14698 THEN
            sigmoid_f := 2;
        ELSIF x =- 14697 THEN
            sigmoid_f := 2;
        ELSIF x =- 14696 THEN
            sigmoid_f := 2;
        ELSIF x =- 14695 THEN
            sigmoid_f := 2;
        ELSIF x =- 14694 THEN
            sigmoid_f := 2;
        ELSIF x =- 14693 THEN
            sigmoid_f := 2;
        ELSIF x =- 14692 THEN
            sigmoid_f := 2;
        ELSIF x =- 14691 THEN
            sigmoid_f := 2;
        ELSIF x =- 14690 THEN
            sigmoid_f := 2;
        ELSIF x =- 14689 THEN
            sigmoid_f := 2;
        ELSIF x =- 14688 THEN
            sigmoid_f := 2;
        ELSIF x =- 14687 THEN
            sigmoid_f := 2;
        ELSIF x =- 14686 THEN
            sigmoid_f := 2;
        ELSIF x =- 14685 THEN
            sigmoid_f := 2;
        ELSIF x =- 14684 THEN
            sigmoid_f := 2;
        ELSIF x =- 14683 THEN
            sigmoid_f := 2;
        ELSIF x =- 14682 THEN
            sigmoid_f := 2;
        ELSIF x =- 14681 THEN
            sigmoid_f := 2;
        ELSIF x =- 14680 THEN
            sigmoid_f := 2;
        ELSIF x =- 14679 THEN
            sigmoid_f := 2;
        ELSIF x =- 14678 THEN
            sigmoid_f := 2;
        ELSIF x =- 14677 THEN
            sigmoid_f := 2;
        ELSIF x =- 14676 THEN
            sigmoid_f := 2;
        ELSIF x =- 14675 THEN
            sigmoid_f := 2;
        ELSIF x =- 14674 THEN
            sigmoid_f := 2;
        ELSIF x =- 14673 THEN
            sigmoid_f := 2;
        ELSIF x =- 14672 THEN
            sigmoid_f := 2;
        ELSIF x =- 14671 THEN
            sigmoid_f := 2;
        ELSIF x =- 14670 THEN
            sigmoid_f := 2;
        ELSIF x =- 14669 THEN
            sigmoid_f := 2;
        ELSIF x =- 14668 THEN
            sigmoid_f := 2;
        ELSIF x =- 14667 THEN
            sigmoid_f := 2;
        ELSIF x =- 14666 THEN
            sigmoid_f := 2;
        ELSIF x =- 14665 THEN
            sigmoid_f := 2;
        ELSIF x =- 14664 THEN
            sigmoid_f := 2;
        ELSIF x =- 14663 THEN
            sigmoid_f := 2;
        ELSIF x =- 14662 THEN
            sigmoid_f := 2;
        ELSIF x =- 14661 THEN
            sigmoid_f := 2;
        ELSIF x =- 14660 THEN
            sigmoid_f := 2;
        ELSIF x =- 14659 THEN
            sigmoid_f := 2;
        ELSIF x =- 14658 THEN
            sigmoid_f := 2;
        ELSIF x =- 14657 THEN
            sigmoid_f := 2;
        ELSIF x =- 14656 THEN
            sigmoid_f := 2;
        ELSIF x =- 14655 THEN
            sigmoid_f := 2;
        ELSIF x =- 14654 THEN
            sigmoid_f := 2;
        ELSIF x =- 14653 THEN
            sigmoid_f := 2;
        ELSIF x =- 14652 THEN
            sigmoid_f := 2;
        ELSIF x =- 14651 THEN
            sigmoid_f := 2;
        ELSIF x =- 14650 THEN
            sigmoid_f := 2;
        ELSIF x =- 14649 THEN
            sigmoid_f := 2;
        ELSIF x =- 14648 THEN
            sigmoid_f := 2;
        ELSIF x =- 14647 THEN
            sigmoid_f := 2;
        ELSIF x =- 14646 THEN
            sigmoid_f := 2;
        ELSIF x =- 14645 THEN
            sigmoid_f := 2;
        ELSIF x =- 14644 THEN
            sigmoid_f := 2;
        ELSIF x =- 14643 THEN
            sigmoid_f := 2;
        ELSIF x =- 14642 THEN
            sigmoid_f := 2;
        ELSIF x =- 14641 THEN
            sigmoid_f := 2;
        ELSIF x =- 14640 THEN
            sigmoid_f := 2;
        ELSIF x =- 14639 THEN
            sigmoid_f := 2;
        ELSIF x =- 14638 THEN
            sigmoid_f := 2;
        ELSIF x =- 14637 THEN
            sigmoid_f := 2;
        ELSIF x =- 14636 THEN
            sigmoid_f := 2;
        ELSIF x =- 14635 THEN
            sigmoid_f := 2;
        ELSIF x =- 14634 THEN
            sigmoid_f := 2;
        ELSIF x =- 14633 THEN
            sigmoid_f := 2;
        ELSIF x =- 14632 THEN
            sigmoid_f := 2;
        ELSIF x =- 14631 THEN
            sigmoid_f := 2;
        ELSIF x =- 14630 THEN
            sigmoid_f := 2;
        ELSIF x =- 14629 THEN
            sigmoid_f := 2;
        ELSIF x =- 14628 THEN
            sigmoid_f := 2;
        ELSIF x =- 14627 THEN
            sigmoid_f := 2;
        ELSIF x =- 14626 THEN
            sigmoid_f := 2;
        ELSIF x =- 14625 THEN
            sigmoid_f := 2;
        ELSIF x =- 14624 THEN
            sigmoid_f := 2;
        ELSIF x =- 14623 THEN
            sigmoid_f := 2;
        ELSIF x =- 14622 THEN
            sigmoid_f := 2;
        ELSIF x =- 14621 THEN
            sigmoid_f := 2;
        ELSIF x =- 14620 THEN
            sigmoid_f := 2;
        ELSIF x =- 14619 THEN
            sigmoid_f := 2;
        ELSIF x =- 14618 THEN
            sigmoid_f := 2;
        ELSIF x =- 14617 THEN
            sigmoid_f := 2;
        ELSIF x =- 14616 THEN
            sigmoid_f := 2;
        ELSIF x =- 14615 THEN
            sigmoid_f := 2;
        ELSIF x =- 14614 THEN
            sigmoid_f := 2;
        ELSIF x =- 14613 THEN
            sigmoid_f := 2;
        ELSIF x =- 14612 THEN
            sigmoid_f := 2;
        ELSIF x =- 14611 THEN
            sigmoid_f := 2;
        ELSIF x =- 14610 THEN
            sigmoid_f := 2;
        ELSIF x =- 14609 THEN
            sigmoid_f := 2;
        ELSIF x =- 14608 THEN
            sigmoid_f := 2;
        ELSIF x =- 14607 THEN
            sigmoid_f := 2;
        ELSIF x =- 14606 THEN
            sigmoid_f := 2;
        ELSIF x =- 14605 THEN
            sigmoid_f := 2;
        ELSIF x =- 14604 THEN
            sigmoid_f := 2;
        ELSIF x =- 14603 THEN
            sigmoid_f := 2;
        ELSIF x =- 14602 THEN
            sigmoid_f := 2;
        ELSIF x =- 14601 THEN
            sigmoid_f := 2;
        ELSIF x =- 14600 THEN
            sigmoid_f := 2;
        ELSIF x =- 14599 THEN
            sigmoid_f := 2;
        ELSIF x =- 14598 THEN
            sigmoid_f := 2;
        ELSIF x =- 14597 THEN
            sigmoid_f := 2;
        ELSIF x =- 14596 THEN
            sigmoid_f := 2;
        ELSIF x =- 14595 THEN
            sigmoid_f := 2;
        ELSIF x =- 14594 THEN
            sigmoid_f := 2;
        ELSIF x =- 14593 THEN
            sigmoid_f := 2;
        ELSIF x =- 14592 THEN
            sigmoid_f := 2;
        ELSIF x =- 14591 THEN
            sigmoid_f := 2;
        ELSIF x =- 14590 THEN
            sigmoid_f := 2;
        ELSIF x =- 14589 THEN
            sigmoid_f := 2;
        ELSIF x =- 14588 THEN
            sigmoid_f := 2;
        ELSIF x =- 14587 THEN
            sigmoid_f := 2;
        ELSIF x =- 14586 THEN
            sigmoid_f := 2;
        ELSIF x =- 14585 THEN
            sigmoid_f := 2;
        ELSIF x =- 14584 THEN
            sigmoid_f := 2;
        ELSIF x =- 14583 THEN
            sigmoid_f := 2;
        ELSIF x =- 14582 THEN
            sigmoid_f := 2;
        ELSIF x =- 14581 THEN
            sigmoid_f := 2;
        ELSIF x =- 14580 THEN
            sigmoid_f := 2;
        ELSIF x =- 14579 THEN
            sigmoid_f := 2;
        ELSIF x =- 14578 THEN
            sigmoid_f := 2;
        ELSIF x =- 14577 THEN
            sigmoid_f := 2;
        ELSIF x =- 14576 THEN
            sigmoid_f := 2;
        ELSIF x =- 14575 THEN
            sigmoid_f := 2;
        ELSIF x =- 14574 THEN
            sigmoid_f := 2;
        ELSIF x =- 14573 THEN
            sigmoid_f := 2;
        ELSIF x =- 14572 THEN
            sigmoid_f := 2;
        ELSIF x =- 14571 THEN
            sigmoid_f := 2;
        ELSIF x =- 14570 THEN
            sigmoid_f := 2;
        ELSIF x =- 14569 THEN
            sigmoid_f := 2;
        ELSIF x =- 14568 THEN
            sigmoid_f := 2;
        ELSIF x =- 14567 THEN
            sigmoid_f := 2;
        ELSIF x =- 14566 THEN
            sigmoid_f := 2;
        ELSIF x =- 14565 THEN
            sigmoid_f := 2;
        ELSIF x =- 14564 THEN
            sigmoid_f := 2;
        ELSIF x =- 14563 THEN
            sigmoid_f := 2;
        ELSIF x =- 14562 THEN
            sigmoid_f := 2;
        ELSIF x =- 14561 THEN
            sigmoid_f := 2;
        ELSIF x =- 14560 THEN
            sigmoid_f := 2;
        ELSIF x =- 14559 THEN
            sigmoid_f := 2;
        ELSIF x =- 14558 THEN
            sigmoid_f := 2;
        ELSIF x =- 14557 THEN
            sigmoid_f := 2;
        ELSIF x =- 14556 THEN
            sigmoid_f := 2;
        ELSIF x =- 14555 THEN
            sigmoid_f := 2;
        ELSIF x =- 14554 THEN
            sigmoid_f := 2;
        ELSIF x =- 14553 THEN
            sigmoid_f := 2;
        ELSIF x =- 14552 THEN
            sigmoid_f := 2;
        ELSIF x =- 14551 THEN
            sigmoid_f := 2;
        ELSIF x =- 14550 THEN
            sigmoid_f := 2;
        ELSIF x =- 14549 THEN
            sigmoid_f := 2;
        ELSIF x =- 14548 THEN
            sigmoid_f := 2;
        ELSIF x =- 14547 THEN
            sigmoid_f := 2;
        ELSIF x =- 14546 THEN
            sigmoid_f := 2;
        ELSIF x =- 14545 THEN
            sigmoid_f := 2;
        ELSIF x =- 14544 THEN
            sigmoid_f := 2;
        ELSIF x =- 14543 THEN
            sigmoid_f := 2;
        ELSIF x =- 14542 THEN
            sigmoid_f := 2;
        ELSIF x =- 14541 THEN
            sigmoid_f := 2;
        ELSIF x =- 14540 THEN
            sigmoid_f := 2;
        ELSIF x =- 14539 THEN
            sigmoid_f := 2;
        ELSIF x =- 14538 THEN
            sigmoid_f := 2;
        ELSIF x =- 14537 THEN
            sigmoid_f := 2;
        ELSIF x =- 14536 THEN
            sigmoid_f := 2;
        ELSIF x =- 14535 THEN
            sigmoid_f := 2;
        ELSIF x =- 14534 THEN
            sigmoid_f := 2;
        ELSIF x =- 14533 THEN
            sigmoid_f := 2;
        ELSIF x =- 14532 THEN
            sigmoid_f := 2;
        ELSIF x =- 14531 THEN
            sigmoid_f := 2;
        ELSIF x =- 14530 THEN
            sigmoid_f := 2;
        ELSIF x =- 14529 THEN
            sigmoid_f := 2;
        ELSIF x =- 14528 THEN
            sigmoid_f := 2;
        ELSIF x =- 14527 THEN
            sigmoid_f := 2;
        ELSIF x =- 14526 THEN
            sigmoid_f := 2;
        ELSIF x =- 14525 THEN
            sigmoid_f := 2;
        ELSIF x =- 14524 THEN
            sigmoid_f := 2;
        ELSIF x =- 14523 THEN
            sigmoid_f := 2;
        ELSIF x =- 14522 THEN
            sigmoid_f := 2;
        ELSIF x =- 14521 THEN
            sigmoid_f := 2;
        ELSIF x =- 14520 THEN
            sigmoid_f := 2;
        ELSIF x =- 14519 THEN
            sigmoid_f := 2;
        ELSIF x =- 14518 THEN
            sigmoid_f := 2;
        ELSIF x =- 14517 THEN
            sigmoid_f := 2;
        ELSIF x =- 14516 THEN
            sigmoid_f := 2;
        ELSIF x =- 14515 THEN
            sigmoid_f := 2;
        ELSIF x =- 14514 THEN
            sigmoid_f := 2;
        ELSIF x =- 14513 THEN
            sigmoid_f := 2;
        ELSIF x =- 14512 THEN
            sigmoid_f := 2;
        ELSIF x =- 14511 THEN
            sigmoid_f := 2;
        ELSIF x =- 14510 THEN
            sigmoid_f := 2;
        ELSIF x =- 14509 THEN
            sigmoid_f := 2;
        ELSIF x =- 14508 THEN
            sigmoid_f := 2;
        ELSIF x =- 14507 THEN
            sigmoid_f := 2;
        ELSIF x =- 14506 THEN
            sigmoid_f := 2;
        ELSIF x =- 14505 THEN
            sigmoid_f := 2;
        ELSIF x =- 14504 THEN
            sigmoid_f := 2;
        ELSIF x =- 14503 THEN
            sigmoid_f := 2;
        ELSIF x =- 14502 THEN
            sigmoid_f := 2;
        ELSIF x =- 14501 THEN
            sigmoid_f := 2;
        ELSIF x =- 14500 THEN
            sigmoid_f := 2;
        ELSIF x =- 14499 THEN
            sigmoid_f := 2;
        ELSIF x =- 14498 THEN
            sigmoid_f := 2;
        ELSIF x =- 14497 THEN
            sigmoid_f := 2;
        ELSIF x =- 14496 THEN
            sigmoid_f := 2;
        ELSIF x =- 14495 THEN
            sigmoid_f := 2;
        ELSIF x =- 14494 THEN
            sigmoid_f := 2;
        ELSIF x =- 14493 THEN
            sigmoid_f := 2;
        ELSIF x =- 14492 THEN
            sigmoid_f := 2;
        ELSIF x =- 14491 THEN
            sigmoid_f := 2;
        ELSIF x =- 14490 THEN
            sigmoid_f := 2;
        ELSIF x =- 14489 THEN
            sigmoid_f := 2;
        ELSIF x =- 14488 THEN
            sigmoid_f := 2;
        ELSIF x =- 14487 THEN
            sigmoid_f := 2;
        ELSIF x =- 14486 THEN
            sigmoid_f := 2;
        ELSIF x =- 14485 THEN
            sigmoid_f := 2;
        ELSIF x =- 14484 THEN
            sigmoid_f := 2;
        ELSIF x =- 14483 THEN
            sigmoid_f := 2;
        ELSIF x =- 14482 THEN
            sigmoid_f := 2;
        ELSIF x =- 14481 THEN
            sigmoid_f := 2;
        ELSIF x =- 14480 THEN
            sigmoid_f := 2;
        ELSIF x =- 14479 THEN
            sigmoid_f := 2;
        ELSIF x =- 14478 THEN
            sigmoid_f := 2;
        ELSIF x =- 14477 THEN
            sigmoid_f := 2;
        ELSIF x =- 14476 THEN
            sigmoid_f := 2;
        ELSIF x =- 14475 THEN
            sigmoid_f := 2;
        ELSIF x =- 14474 THEN
            sigmoid_f := 2;
        ELSIF x =- 14473 THEN
            sigmoid_f := 2;
        ELSIF x =- 14472 THEN
            sigmoid_f := 2;
        ELSIF x =- 14471 THEN
            sigmoid_f := 2;
        ELSIF x =- 14470 THEN
            sigmoid_f := 2;
        ELSIF x =- 14469 THEN
            sigmoid_f := 2;
        ELSIF x =- 14468 THEN
            sigmoid_f := 2;
        ELSIF x =- 14467 THEN
            sigmoid_f := 2;
        ELSIF x =- 14466 THEN
            sigmoid_f := 2;
        ELSIF x =- 14465 THEN
            sigmoid_f := 2;
        ELSIF x =- 14464 THEN
            sigmoid_f := 2;
        ELSIF x =- 14463 THEN
            sigmoid_f := 2;
        ELSIF x =- 14462 THEN
            sigmoid_f := 2;
        ELSIF x =- 14461 THEN
            sigmoid_f := 2;
        ELSIF x =- 14460 THEN
            sigmoid_f := 2;
        ELSIF x =- 14459 THEN
            sigmoid_f := 2;
        ELSIF x =- 14458 THEN
            sigmoid_f := 2;
        ELSIF x =- 14457 THEN
            sigmoid_f := 2;
        ELSIF x =- 14456 THEN
            sigmoid_f := 2;
        ELSIF x =- 14455 THEN
            sigmoid_f := 2;
        ELSIF x =- 14454 THEN
            sigmoid_f := 2;
        ELSIF x =- 14453 THEN
            sigmoid_f := 2;
        ELSIF x =- 14452 THEN
            sigmoid_f := 2;
        ELSIF x =- 14451 THEN
            sigmoid_f := 2;
        ELSIF x =- 14450 THEN
            sigmoid_f := 2;
        ELSIF x =- 14449 THEN
            sigmoid_f := 2;
        ELSIF x =- 14448 THEN
            sigmoid_f := 2;
        ELSIF x =- 14447 THEN
            sigmoid_f := 2;
        ELSIF x =- 14446 THEN
            sigmoid_f := 2;
        ELSIF x =- 14445 THEN
            sigmoid_f := 2;
        ELSIF x =- 14444 THEN
            sigmoid_f := 2;
        ELSIF x =- 14443 THEN
            sigmoid_f := 2;
        ELSIF x =- 14442 THEN
            sigmoid_f := 2;
        ELSIF x =- 14441 THEN
            sigmoid_f := 2;
        ELSIF x =- 14440 THEN
            sigmoid_f := 2;
        ELSIF x =- 14439 THEN
            sigmoid_f := 2;
        ELSIF x =- 14438 THEN
            sigmoid_f := 2;
        ELSIF x =- 14437 THEN
            sigmoid_f := 2;
        ELSIF x =- 14436 THEN
            sigmoid_f := 2;
        ELSIF x =- 14435 THEN
            sigmoid_f := 2;
        ELSIF x =- 14434 THEN
            sigmoid_f := 2;
        ELSIF x =- 14433 THEN
            sigmoid_f := 2;
        ELSIF x =- 14432 THEN
            sigmoid_f := 2;
        ELSIF x =- 14431 THEN
            sigmoid_f := 2;
        ELSIF x =- 14430 THEN
            sigmoid_f := 2;
        ELSIF x =- 14429 THEN
            sigmoid_f := 2;
        ELSIF x =- 14428 THEN
            sigmoid_f := 2;
        ELSIF x =- 14427 THEN
            sigmoid_f := 2;
        ELSIF x =- 14426 THEN
            sigmoid_f := 2;
        ELSIF x =- 14425 THEN
            sigmoid_f := 2;
        ELSIF x =- 14424 THEN
            sigmoid_f := 2;
        ELSIF x =- 14423 THEN
            sigmoid_f := 2;
        ELSIF x =- 14422 THEN
            sigmoid_f := 2;
        ELSIF x =- 14421 THEN
            sigmoid_f := 2;
        ELSIF x =- 14420 THEN
            sigmoid_f := 2;
        ELSIF x =- 14419 THEN
            sigmoid_f := 2;
        ELSIF x =- 14418 THEN
            sigmoid_f := 2;
        ELSIF x =- 14417 THEN
            sigmoid_f := 2;
        ELSIF x =- 14416 THEN
            sigmoid_f := 2;
        ELSIF x =- 14415 THEN
            sigmoid_f := 2;
        ELSIF x =- 14414 THEN
            sigmoid_f := 2;
        ELSIF x =- 14413 THEN
            sigmoid_f := 2;
        ELSIF x =- 14412 THEN
            sigmoid_f := 2;
        ELSIF x =- 14411 THEN
            sigmoid_f := 2;
        ELSIF x =- 14410 THEN
            sigmoid_f := 2;
        ELSIF x =- 14409 THEN
            sigmoid_f := 2;
        ELSIF x =- 14408 THEN
            sigmoid_f := 2;
        ELSIF x =- 14407 THEN
            sigmoid_f := 2;
        ELSIF x =- 14406 THEN
            sigmoid_f := 2;
        ELSIF x =- 14405 THEN
            sigmoid_f := 2;
        ELSIF x =- 14404 THEN
            sigmoid_f := 2;
        ELSIF x =- 14403 THEN
            sigmoid_f := 2;
        ELSIF x =- 14402 THEN
            sigmoid_f := 2;
        ELSIF x =- 14401 THEN
            sigmoid_f := 2;
        ELSIF x =- 14400 THEN
            sigmoid_f := 2;
        ELSIF x =- 14399 THEN
            sigmoid_f := 2;
        ELSIF x =- 14398 THEN
            sigmoid_f := 2;
        ELSIF x =- 14397 THEN
            sigmoid_f := 2;
        ELSIF x =- 14396 THEN
            sigmoid_f := 2;
        ELSIF x =- 14395 THEN
            sigmoid_f := 2;
        ELSIF x =- 14394 THEN
            sigmoid_f := 2;
        ELSIF x =- 14393 THEN
            sigmoid_f := 2;
        ELSIF x =- 14392 THEN
            sigmoid_f := 2;
        ELSIF x =- 14391 THEN
            sigmoid_f := 2;
        ELSIF x =- 14390 THEN
            sigmoid_f := 2;
        ELSIF x =- 14389 THEN
            sigmoid_f := 2;
        ELSIF x =- 14388 THEN
            sigmoid_f := 2;
        ELSIF x =- 14387 THEN
            sigmoid_f := 2;
        ELSIF x =- 14386 THEN
            sigmoid_f := 2;
        ELSIF x =- 14385 THEN
            sigmoid_f := 2;
        ELSIF x =- 14384 THEN
            sigmoid_f := 2;
        ELSIF x =- 14383 THEN
            sigmoid_f := 2;
        ELSIF x =- 14382 THEN
            sigmoid_f := 2;
        ELSIF x =- 14381 THEN
            sigmoid_f := 2;
        ELSIF x =- 14380 THEN
            sigmoid_f := 2;
        ELSIF x =- 14379 THEN
            sigmoid_f := 2;
        ELSIF x =- 14378 THEN
            sigmoid_f := 2;
        ELSIF x =- 14377 THEN
            sigmoid_f := 2;
        ELSIF x =- 14376 THEN
            sigmoid_f := 2;
        ELSIF x =- 14375 THEN
            sigmoid_f := 2;
        ELSIF x =- 14374 THEN
            sigmoid_f := 2;
        ELSIF x =- 14373 THEN
            sigmoid_f := 2;
        ELSIF x =- 14372 THEN
            sigmoid_f := 2;
        ELSIF x =- 14371 THEN
            sigmoid_f := 2;
        ELSIF x =- 14370 THEN
            sigmoid_f := 2;
        ELSIF x =- 14369 THEN
            sigmoid_f := 2;
        ELSIF x =- 14368 THEN
            sigmoid_f := 2;
        ELSIF x =- 14367 THEN
            sigmoid_f := 2;
        ELSIF x =- 14366 THEN
            sigmoid_f := 2;
        ELSIF x =- 14365 THEN
            sigmoid_f := 2;
        ELSIF x =- 14364 THEN
            sigmoid_f := 2;
        ELSIF x =- 14363 THEN
            sigmoid_f := 2;
        ELSIF x =- 14362 THEN
            sigmoid_f := 2;
        ELSIF x =- 14361 THEN
            sigmoid_f := 2;
        ELSIF x =- 14360 THEN
            sigmoid_f := 2;
        ELSIF x =- 14359 THEN
            sigmoid_f := 2;
        ELSIF x =- 14358 THEN
            sigmoid_f := 2;
        ELSIF x =- 14357 THEN
            sigmoid_f := 2;
        ELSIF x =- 14356 THEN
            sigmoid_f := 2;
        ELSIF x =- 14355 THEN
            sigmoid_f := 2;
        ELSIF x =- 14354 THEN
            sigmoid_f := 2;
        ELSIF x =- 14353 THEN
            sigmoid_f := 2;
        ELSIF x =- 14352 THEN
            sigmoid_f := 2;
        ELSIF x =- 14351 THEN
            sigmoid_f := 2;
        ELSIF x =- 14350 THEN
            sigmoid_f := 2;
        ELSIF x =- 14349 THEN
            sigmoid_f := 2;
        ELSIF x =- 14348 THEN
            sigmoid_f := 2;
        ELSIF x =- 14347 THEN
            sigmoid_f := 2;
        ELSIF x =- 14346 THEN
            sigmoid_f := 2;
        ELSIF x =- 14345 THEN
            sigmoid_f := 2;
        ELSIF x =- 14344 THEN
            sigmoid_f := 2;
        ELSIF x =- 14343 THEN
            sigmoid_f := 2;
        ELSIF x =- 14342 THEN
            sigmoid_f := 2;
        ELSIF x =- 14341 THEN
            sigmoid_f := 2;
        ELSIF x =- 14340 THEN
            sigmoid_f := 2;
        ELSIF x =- 14339 THEN
            sigmoid_f := 2;
        ELSIF x =- 14338 THEN
            sigmoid_f := 2;
        ELSIF x =- 14337 THEN
            sigmoid_f := 2;
        ELSIF x =- 14336 THEN
            sigmoid_f := 2;
        ELSIF x =- 14335 THEN
            sigmoid_f := 2;
        ELSIF x =- 14334 THEN
            sigmoid_f := 2;
        ELSIF x =- 14333 THEN
            sigmoid_f := 2;
        ELSIF x =- 14332 THEN
            sigmoid_f := 2;
        ELSIF x =- 14331 THEN
            sigmoid_f := 2;
        ELSIF x =- 14330 THEN
            sigmoid_f := 2;
        ELSIF x =- 14329 THEN
            sigmoid_f := 2;
        ELSIF x =- 14328 THEN
            sigmoid_f := 2;
        ELSIF x =- 14327 THEN
            sigmoid_f := 2;
        ELSIF x =- 14326 THEN
            sigmoid_f := 2;
        ELSIF x =- 14325 THEN
            sigmoid_f := 2;
        ELSIF x =- 14324 THEN
            sigmoid_f := 2;
        ELSIF x =- 14323 THEN
            sigmoid_f := 2;
        ELSIF x =- 14322 THEN
            sigmoid_f := 2;
        ELSIF x =- 14321 THEN
            sigmoid_f := 2;
        ELSIF x =- 14320 THEN
            sigmoid_f := 2;
        ELSIF x =- 14319 THEN
            sigmoid_f := 2;
        ELSIF x =- 14318 THEN
            sigmoid_f := 2;
        ELSIF x =- 14317 THEN
            sigmoid_f := 2;
        ELSIF x =- 14316 THEN
            sigmoid_f := 2;
        ELSIF x =- 14315 THEN
            sigmoid_f := 2;
        ELSIF x =- 14314 THEN
            sigmoid_f := 2;
        ELSIF x =- 14313 THEN
            sigmoid_f := 2;
        ELSIF x =- 14312 THEN
            sigmoid_f := 2;
        ELSIF x =- 14311 THEN
            sigmoid_f := 2;
        ELSIF x =- 14310 THEN
            sigmoid_f := 2;
        ELSIF x =- 14309 THEN
            sigmoid_f := 2;
        ELSIF x =- 14308 THEN
            sigmoid_f := 2;
        ELSIF x =- 14307 THEN
            sigmoid_f := 2;
        ELSIF x =- 14306 THEN
            sigmoid_f := 2;
        ELSIF x =- 14305 THEN
            sigmoid_f := 2;
        ELSIF x =- 14304 THEN
            sigmoid_f := 2;
        ELSIF x =- 14303 THEN
            sigmoid_f := 2;
        ELSIF x =- 14302 THEN
            sigmoid_f := 2;
        ELSIF x =- 14301 THEN
            sigmoid_f := 2;
        ELSIF x =- 14300 THEN
            sigmoid_f := 2;
        ELSIF x =- 14299 THEN
            sigmoid_f := 2;
        ELSIF x =- 14298 THEN
            sigmoid_f := 2;
        ELSIF x =- 14297 THEN
            sigmoid_f := 2;
        ELSIF x =- 14296 THEN
            sigmoid_f := 2;
        ELSIF x =- 14295 THEN
            sigmoid_f := 2;
        ELSIF x =- 14294 THEN
            sigmoid_f := 2;
        ELSIF x =- 14293 THEN
            sigmoid_f := 2;
        ELSIF x =- 14292 THEN
            sigmoid_f := 2;
        ELSIF x =- 14291 THEN
            sigmoid_f := 2;
        ELSIF x =- 14290 THEN
            sigmoid_f := 2;
        ELSIF x =- 14289 THEN
            sigmoid_f := 2;
        ELSIF x =- 14288 THEN
            sigmoid_f := 2;
        ELSIF x =- 14287 THEN
            sigmoid_f := 2;
        ELSIF x =- 14286 THEN
            sigmoid_f := 2;
        ELSIF x =- 14285 THEN
            sigmoid_f := 2;
        ELSIF x =- 14284 THEN
            sigmoid_f := 2;
        ELSIF x =- 14283 THEN
            sigmoid_f := 2;
        ELSIF x =- 14282 THEN
            sigmoid_f := 2;
        ELSIF x =- 14281 THEN
            sigmoid_f := 2;
        ELSIF x =- 14280 THEN
            sigmoid_f := 2;
        ELSIF x =- 14279 THEN
            sigmoid_f := 2;
        ELSIF x =- 14278 THEN
            sigmoid_f := 2;
        ELSIF x =- 14277 THEN
            sigmoid_f := 2;
        ELSIF x =- 14276 THEN
            sigmoid_f := 2;
        ELSIF x =- 14275 THEN
            sigmoid_f := 2;
        ELSIF x =- 14274 THEN
            sigmoid_f := 2;
        ELSIF x =- 14273 THEN
            sigmoid_f := 2;
        ELSIF x =- 14272 THEN
            sigmoid_f := 2;
        ELSIF x =- 14271 THEN
            sigmoid_f := 2;
        ELSIF x =- 14270 THEN
            sigmoid_f := 2;
        ELSIF x =- 14269 THEN
            sigmoid_f := 2;
        ELSIF x =- 14268 THEN
            sigmoid_f := 2;
        ELSIF x =- 14267 THEN
            sigmoid_f := 2;
        ELSIF x =- 14266 THEN
            sigmoid_f := 2;
        ELSIF x =- 14265 THEN
            sigmoid_f := 2;
        ELSIF x =- 14264 THEN
            sigmoid_f := 2;
        ELSIF x =- 14263 THEN
            sigmoid_f := 2;
        ELSIF x =- 14262 THEN
            sigmoid_f := 2;
        ELSIF x =- 14261 THEN
            sigmoid_f := 2;
        ELSIF x =- 14260 THEN
            sigmoid_f := 2;
        ELSIF x =- 14259 THEN
            sigmoid_f := 2;
        ELSIF x =- 14258 THEN
            sigmoid_f := 2;
        ELSIF x =- 14257 THEN
            sigmoid_f := 2;
        ELSIF x =- 14256 THEN
            sigmoid_f := 2;
        ELSIF x =- 14255 THEN
            sigmoid_f := 2;
        ELSIF x =- 14254 THEN
            sigmoid_f := 2;
        ELSIF x =- 14253 THEN
            sigmoid_f := 2;
        ELSIF x =- 14252 THEN
            sigmoid_f := 2;
        ELSIF x =- 14251 THEN
            sigmoid_f := 2;
        ELSIF x =- 14250 THEN
            sigmoid_f := 2;
        ELSIF x =- 14249 THEN
            sigmoid_f := 2;
        ELSIF x =- 14248 THEN
            sigmoid_f := 2;
        ELSIF x =- 14247 THEN
            sigmoid_f := 2;
        ELSIF x =- 14246 THEN
            sigmoid_f := 2;
        ELSIF x =- 14245 THEN
            sigmoid_f := 2;
        ELSIF x =- 14244 THEN
            sigmoid_f := 2;
        ELSIF x =- 14243 THEN
            sigmoid_f := 2;
        ELSIF x =- 14242 THEN
            sigmoid_f := 2;
        ELSIF x =- 14241 THEN
            sigmoid_f := 2;
        ELSIF x =- 14240 THEN
            sigmoid_f := 2;
        ELSIF x =- 14239 THEN
            sigmoid_f := 2;
        ELSIF x =- 14238 THEN
            sigmoid_f := 2;
        ELSIF x =- 14237 THEN
            sigmoid_f := 2;
        ELSIF x =- 14236 THEN
            sigmoid_f := 2;
        ELSIF x =- 14235 THEN
            sigmoid_f := 2;
        ELSIF x =- 14234 THEN
            sigmoid_f := 2;
        ELSIF x =- 14233 THEN
            sigmoid_f := 2;
        ELSIF x =- 14232 THEN
            sigmoid_f := 2;
        ELSIF x =- 14231 THEN
            sigmoid_f := 2;
        ELSIF x =- 14230 THEN
            sigmoid_f := 2;
        ELSIF x =- 14229 THEN
            sigmoid_f := 2;
        ELSIF x =- 14228 THEN
            sigmoid_f := 2;
        ELSIF x =- 14227 THEN
            sigmoid_f := 2;
        ELSIF x =- 14226 THEN
            sigmoid_f := 2;
        ELSIF x =- 14225 THEN
            sigmoid_f := 2;
        ELSIF x =- 14224 THEN
            sigmoid_f := 2;
        ELSIF x =- 14223 THEN
            sigmoid_f := 2;
        ELSIF x =- 14222 THEN
            sigmoid_f := 2;
        ELSIF x =- 14221 THEN
            sigmoid_f := 2;
        ELSIF x =- 14220 THEN
            sigmoid_f := 2;
        ELSIF x =- 14219 THEN
            sigmoid_f := 2;
        ELSIF x =- 14218 THEN
            sigmoid_f := 2;
        ELSIF x =- 14217 THEN
            sigmoid_f := 2;
        ELSIF x =- 14216 THEN
            sigmoid_f := 2;
        ELSIF x =- 14215 THEN
            sigmoid_f := 2;
        ELSIF x =- 14214 THEN
            sigmoid_f := 2;
        ELSIF x =- 14213 THEN
            sigmoid_f := 2;
        ELSIF x =- 14212 THEN
            sigmoid_f := 2;
        ELSIF x =- 14211 THEN
            sigmoid_f := 2;
        ELSIF x =- 14210 THEN
            sigmoid_f := 2;
        ELSIF x =- 14209 THEN
            sigmoid_f := 2;
        ELSIF x =- 14208 THEN
            sigmoid_f := 2;
        ELSIF x =- 14207 THEN
            sigmoid_f := 2;
        ELSIF x =- 14206 THEN
            sigmoid_f := 2;
        ELSIF x =- 14205 THEN
            sigmoid_f := 2;
        ELSIF x =- 14204 THEN
            sigmoid_f := 2;
        ELSIF x =- 14203 THEN
            sigmoid_f := 2;
        ELSIF x =- 14202 THEN
            sigmoid_f := 2;
        ELSIF x =- 14201 THEN
            sigmoid_f := 2;
        ELSIF x =- 14200 THEN
            sigmoid_f := 2;
        ELSIF x =- 14199 THEN
            sigmoid_f := 2;
        ELSIF x =- 14198 THEN
            sigmoid_f := 2;
        ELSIF x =- 14197 THEN
            sigmoid_f := 2;
        ELSIF x =- 14196 THEN
            sigmoid_f := 2;
        ELSIF x =- 14195 THEN
            sigmoid_f := 2;
        ELSIF x =- 14194 THEN
            sigmoid_f := 2;
        ELSIF x =- 14193 THEN
            sigmoid_f := 2;
        ELSIF x =- 14192 THEN
            sigmoid_f := 2;
        ELSIF x =- 14191 THEN
            sigmoid_f := 2;
        ELSIF x =- 14190 THEN
            sigmoid_f := 2;
        ELSIF x =- 14189 THEN
            sigmoid_f := 2;
        ELSIF x =- 14188 THEN
            sigmoid_f := 2;
        ELSIF x =- 14187 THEN
            sigmoid_f := 2;
        ELSIF x =- 14186 THEN
            sigmoid_f := 2;
        ELSIF x =- 14185 THEN
            sigmoid_f := 2;
        ELSIF x =- 14184 THEN
            sigmoid_f := 2;
        ELSIF x =- 14183 THEN
            sigmoid_f := 2;
        ELSIF x =- 14182 THEN
            sigmoid_f := 2;
        ELSIF x =- 14181 THEN
            sigmoid_f := 2;
        ELSIF x =- 14180 THEN
            sigmoid_f := 2;
        ELSIF x =- 14179 THEN
            sigmoid_f := 2;
        ELSIF x =- 14178 THEN
            sigmoid_f := 2;
        ELSIF x =- 14177 THEN
            sigmoid_f := 2;
        ELSIF x =- 14176 THEN
            sigmoid_f := 2;
        ELSIF x =- 14175 THEN
            sigmoid_f := 2;
        ELSIF x =- 14174 THEN
            sigmoid_f := 2;
        ELSIF x =- 14173 THEN
            sigmoid_f := 2;
        ELSIF x =- 14172 THEN
            sigmoid_f := 2;
        ELSIF x =- 14171 THEN
            sigmoid_f := 2;
        ELSIF x =- 14170 THEN
            sigmoid_f := 2;
        ELSIF x =- 14169 THEN
            sigmoid_f := 2;
        ELSIF x =- 14168 THEN
            sigmoid_f := 2;
        ELSIF x =- 14167 THEN
            sigmoid_f := 2;
        ELSIF x =- 14166 THEN
            sigmoid_f := 2;
        ELSIF x =- 14165 THEN
            sigmoid_f := 2;
        ELSIF x =- 14164 THEN
            sigmoid_f := 2;
        ELSIF x =- 14163 THEN
            sigmoid_f := 2;
        ELSIF x =- 14162 THEN
            sigmoid_f := 2;
        ELSIF x =- 14161 THEN
            sigmoid_f := 2;
        ELSIF x =- 14160 THEN
            sigmoid_f := 2;
        ELSIF x =- 14159 THEN
            sigmoid_f := 2;
        ELSIF x =- 14158 THEN
            sigmoid_f := 2;
        ELSIF x =- 14157 THEN
            sigmoid_f := 2;
        ELSIF x =- 14156 THEN
            sigmoid_f := 2;
        ELSIF x =- 14155 THEN
            sigmoid_f := 2;
        ELSIF x =- 14154 THEN
            sigmoid_f := 2;
        ELSIF x =- 14153 THEN
            sigmoid_f := 2;
        ELSIF x =- 14152 THEN
            sigmoid_f := 2;
        ELSIF x =- 14151 THEN
            sigmoid_f := 2;
        ELSIF x =- 14150 THEN
            sigmoid_f := 2;
        ELSIF x =- 14149 THEN
            sigmoid_f := 2;
        ELSIF x =- 14148 THEN
            sigmoid_f := 2;
        ELSIF x =- 14147 THEN
            sigmoid_f := 2;
        ELSIF x =- 14146 THEN
            sigmoid_f := 2;
        ELSIF x =- 14145 THEN
            sigmoid_f := 2;
        ELSIF x =- 14144 THEN
            sigmoid_f := 2;
        ELSIF x =- 14143 THEN
            sigmoid_f := 2;
        ELSIF x =- 14142 THEN
            sigmoid_f := 2;
        ELSIF x =- 14141 THEN
            sigmoid_f := 2;
        ELSIF x =- 14140 THEN
            sigmoid_f := 2;
        ELSIF x =- 14139 THEN
            sigmoid_f := 2;
        ELSIF x =- 14138 THEN
            sigmoid_f := 2;
        ELSIF x =- 14137 THEN
            sigmoid_f := 2;
        ELSIF x =- 14136 THEN
            sigmoid_f := 2;
        ELSIF x =- 14135 THEN
            sigmoid_f := 2;
        ELSIF x =- 14134 THEN
            sigmoid_f := 2;
        ELSIF x =- 14133 THEN
            sigmoid_f := 2;
        ELSIF x =- 14132 THEN
            sigmoid_f := 2;
        ELSIF x =- 14131 THEN
            sigmoid_f := 2;
        ELSIF x =- 14130 THEN
            sigmoid_f := 2;
        ELSIF x =- 14129 THEN
            sigmoid_f := 2;
        ELSIF x =- 14128 THEN
            sigmoid_f := 2;
        ELSIF x =- 14127 THEN
            sigmoid_f := 2;
        ELSIF x =- 14126 THEN
            sigmoid_f := 2;
        ELSIF x =- 14125 THEN
            sigmoid_f := 2;
        ELSIF x =- 14124 THEN
            sigmoid_f := 2;
        ELSIF x =- 14123 THEN
            sigmoid_f := 2;
        ELSIF x =- 14122 THEN
            sigmoid_f := 2;
        ELSIF x =- 14121 THEN
            sigmoid_f := 2;
        ELSIF x =- 14120 THEN
            sigmoid_f := 2;
        ELSIF x =- 14119 THEN
            sigmoid_f := 2;
        ELSIF x =- 14118 THEN
            sigmoid_f := 2;
        ELSIF x =- 14117 THEN
            sigmoid_f := 2;
        ELSIF x =- 14116 THEN
            sigmoid_f := 2;
        ELSIF x =- 14115 THEN
            sigmoid_f := 2;
        ELSIF x =- 14114 THEN
            sigmoid_f := 2;
        ELSIF x =- 14113 THEN
            sigmoid_f := 2;
        ELSIF x =- 14112 THEN
            sigmoid_f := 2;
        ELSIF x =- 14111 THEN
            sigmoid_f := 2;
        ELSIF x =- 14110 THEN
            sigmoid_f := 2;
        ELSIF x =- 14109 THEN
            sigmoid_f := 2;
        ELSIF x =- 14108 THEN
            sigmoid_f := 2;
        ELSIF x =- 14107 THEN
            sigmoid_f := 2;
        ELSIF x =- 14106 THEN
            sigmoid_f := 2;
        ELSIF x =- 14105 THEN
            sigmoid_f := 2;
        ELSIF x =- 14104 THEN
            sigmoid_f := 2;
        ELSIF x =- 14103 THEN
            sigmoid_f := 2;
        ELSIF x =- 14102 THEN
            sigmoid_f := 2;
        ELSIF x =- 14101 THEN
            sigmoid_f := 2;
        ELSIF x =- 14100 THEN
            sigmoid_f := 2;
        ELSIF x =- 14099 THEN
            sigmoid_f := 2;
        ELSIF x =- 14098 THEN
            sigmoid_f := 2;
        ELSIF x =- 14097 THEN
            sigmoid_f := 2;
        ELSIF x =- 14096 THEN
            sigmoid_f := 2;
        ELSIF x =- 14095 THEN
            sigmoid_f := 2;
        ELSIF x =- 14094 THEN
            sigmoid_f := 2;
        ELSIF x =- 14093 THEN
            sigmoid_f := 2;
        ELSIF x =- 14092 THEN
            sigmoid_f := 2;
        ELSIF x =- 14091 THEN
            sigmoid_f := 2;
        ELSIF x =- 14090 THEN
            sigmoid_f := 2;
        ELSIF x =- 14089 THEN
            sigmoid_f := 2;
        ELSIF x =- 14088 THEN
            sigmoid_f := 2;
        ELSIF x =- 14087 THEN
            sigmoid_f := 2;
        ELSIF x =- 14086 THEN
            sigmoid_f := 2;
        ELSIF x =- 14085 THEN
            sigmoid_f := 2;
        ELSIF x =- 14084 THEN
            sigmoid_f := 2;
        ELSIF x =- 14083 THEN
            sigmoid_f := 2;
        ELSIF x =- 14082 THEN
            sigmoid_f := 2;
        ELSIF x =- 14081 THEN
            sigmoid_f := 2;
        ELSIF x =- 14080 THEN
            sigmoid_f := 2;
        ELSIF x =- 14079 THEN
            sigmoid_f := 2;
        ELSIF x =- 14078 THEN
            sigmoid_f := 2;
        ELSIF x =- 14077 THEN
            sigmoid_f := 2;
        ELSIF x =- 14076 THEN
            sigmoid_f := 2;
        ELSIF x =- 14075 THEN
            sigmoid_f := 2;
        ELSIF x =- 14074 THEN
            sigmoid_f := 2;
        ELSIF x =- 14073 THEN
            sigmoid_f := 2;
        ELSIF x =- 14072 THEN
            sigmoid_f := 2;
        ELSIF x =- 14071 THEN
            sigmoid_f := 2;
        ELSIF x =- 14070 THEN
            sigmoid_f := 2;
        ELSIF x =- 14069 THEN
            sigmoid_f := 2;
        ELSIF x =- 14068 THEN
            sigmoid_f := 2;
        ELSIF x =- 14067 THEN
            sigmoid_f := 2;
        ELSIF x =- 14066 THEN
            sigmoid_f := 2;
        ELSIF x =- 14065 THEN
            sigmoid_f := 2;
        ELSIF x =- 14064 THEN
            sigmoid_f := 2;
        ELSIF x =- 14063 THEN
            sigmoid_f := 2;
        ELSIF x =- 14062 THEN
            sigmoid_f := 2;
        ELSIF x =- 14061 THEN
            sigmoid_f := 2;
        ELSIF x =- 14060 THEN
            sigmoid_f := 2;
        ELSIF x =- 14059 THEN
            sigmoid_f := 2;
        ELSIF x =- 14058 THEN
            sigmoid_f := 2;
        ELSIF x =- 14057 THEN
            sigmoid_f := 2;
        ELSIF x =- 14056 THEN
            sigmoid_f := 2;
        ELSIF x =- 14055 THEN
            sigmoid_f := 2;
        ELSIF x =- 14054 THEN
            sigmoid_f := 2;
        ELSIF x =- 14053 THEN
            sigmoid_f := 2;
        ELSIF x =- 14052 THEN
            sigmoid_f := 2;
        ELSIF x =- 14051 THEN
            sigmoid_f := 2;
        ELSIF x =- 14050 THEN
            sigmoid_f := 2;
        ELSIF x =- 14049 THEN
            sigmoid_f := 2;
        ELSIF x =- 14048 THEN
            sigmoid_f := 2;
        ELSIF x =- 14047 THEN
            sigmoid_f := 2;
        ELSIF x =- 14046 THEN
            sigmoid_f := 2;
        ELSIF x =- 14045 THEN
            sigmoid_f := 2;
        ELSIF x =- 14044 THEN
            sigmoid_f := 2;
        ELSIF x =- 14043 THEN
            sigmoid_f := 2;
        ELSIF x =- 14042 THEN
            sigmoid_f := 2;
        ELSIF x =- 14041 THEN
            sigmoid_f := 2;
        ELSIF x =- 14040 THEN
            sigmoid_f := 2;
        ELSIF x =- 14039 THEN
            sigmoid_f := 2;
        ELSIF x =- 14038 THEN
            sigmoid_f := 2;
        ELSIF x =- 14037 THEN
            sigmoid_f := 2;
        ELSIF x =- 14036 THEN
            sigmoid_f := 2;
        ELSIF x =- 14035 THEN
            sigmoid_f := 2;
        ELSIF x =- 14034 THEN
            sigmoid_f := 2;
        ELSIF x =- 14033 THEN
            sigmoid_f := 2;
        ELSIF x =- 14032 THEN
            sigmoid_f := 2;
        ELSIF x =- 14031 THEN
            sigmoid_f := 2;
        ELSIF x =- 14030 THEN
            sigmoid_f := 2;
        ELSIF x =- 14029 THEN
            sigmoid_f := 2;
        ELSIF x =- 14028 THEN
            sigmoid_f := 2;
        ELSIF x =- 14027 THEN
            sigmoid_f := 2;
        ELSIF x =- 14026 THEN
            sigmoid_f := 2;
        ELSIF x =- 14025 THEN
            sigmoid_f := 2;
        ELSIF x =- 14024 THEN
            sigmoid_f := 2;
        ELSIF x =- 14023 THEN
            sigmoid_f := 2;
        ELSIF x =- 14022 THEN
            sigmoid_f := 2;
        ELSIF x =- 14021 THEN
            sigmoid_f := 2;
        ELSIF x =- 14020 THEN
            sigmoid_f := 2;
        ELSIF x =- 14019 THEN
            sigmoid_f := 2;
        ELSIF x =- 14018 THEN
            sigmoid_f := 2;
        ELSIF x =- 14017 THEN
            sigmoid_f := 2;
        ELSIF x =- 14016 THEN
            sigmoid_f := 2;
        ELSIF x =- 14015 THEN
            sigmoid_f := 2;
        ELSIF x =- 14014 THEN
            sigmoid_f := 2;
        ELSIF x =- 14013 THEN
            sigmoid_f := 2;
        ELSIF x =- 14012 THEN
            sigmoid_f := 2;
        ELSIF x =- 14011 THEN
            sigmoid_f := 2;
        ELSIF x =- 14010 THEN
            sigmoid_f := 2;
        ELSIF x =- 14009 THEN
            sigmoid_f := 2;
        ELSIF x =- 14008 THEN
            sigmoid_f := 2;
        ELSIF x =- 14007 THEN
            sigmoid_f := 2;
        ELSIF x =- 14006 THEN
            sigmoid_f := 2;
        ELSIF x =- 14005 THEN
            sigmoid_f := 2;
        ELSIF x =- 14004 THEN
            sigmoid_f := 2;
        ELSIF x =- 14003 THEN
            sigmoid_f := 2;
        ELSIF x =- 14002 THEN
            sigmoid_f := 2;
        ELSIF x =- 14001 THEN
            sigmoid_f := 2;
        ELSIF x =- 14000 THEN
            sigmoid_f := 2;
        ELSIF x =- 13999 THEN
            sigmoid_f := 2;
        ELSIF x =- 13998 THEN
            sigmoid_f := 2;
        ELSIF x =- 13997 THEN
            sigmoid_f := 2;
        ELSIF x =- 13996 THEN
            sigmoid_f := 2;
        ELSIF x =- 13995 THEN
            sigmoid_f := 2;
        ELSIF x =- 13994 THEN
            sigmoid_f := 2;
        ELSIF x =- 13993 THEN
            sigmoid_f := 2;
        ELSIF x =- 13992 THEN
            sigmoid_f := 2;
        ELSIF x =- 13991 THEN
            sigmoid_f := 2;
        ELSIF x =- 13990 THEN
            sigmoid_f := 2;
        ELSIF x =- 13989 THEN
            sigmoid_f := 2;
        ELSIF x =- 13988 THEN
            sigmoid_f := 2;
        ELSIF x =- 13987 THEN
            sigmoid_f := 2;
        ELSIF x =- 13986 THEN
            sigmoid_f := 2;
        ELSIF x =- 13985 THEN
            sigmoid_f := 2;
        ELSIF x =- 13984 THEN
            sigmoid_f := 2;
        ELSIF x =- 13983 THEN
            sigmoid_f := 2;
        ELSIF x =- 13982 THEN
            sigmoid_f := 2;
        ELSIF x =- 13981 THEN
            sigmoid_f := 2;
        ELSIF x =- 13980 THEN
            sigmoid_f := 2;
        ELSIF x =- 13979 THEN
            sigmoid_f := 2;
        ELSIF x =- 13978 THEN
            sigmoid_f := 2;
        ELSIF x =- 13977 THEN
            sigmoid_f := 2;
        ELSIF x =- 13976 THEN
            sigmoid_f := 2;
        ELSIF x =- 13975 THEN
            sigmoid_f := 2;
        ELSIF x =- 13974 THEN
            sigmoid_f := 2;
        ELSIF x =- 13973 THEN
            sigmoid_f := 2;
        ELSIF x =- 13972 THEN
            sigmoid_f := 2;
        ELSIF x =- 13971 THEN
            sigmoid_f := 2;
        ELSIF x =- 13970 THEN
            sigmoid_f := 2;
        ELSIF x =- 13969 THEN
            sigmoid_f := 2;
        ELSIF x =- 13968 THEN
            sigmoid_f := 2;
        ELSIF x =- 13967 THEN
            sigmoid_f := 2;
        ELSIF x =- 13966 THEN
            sigmoid_f := 2;
        ELSIF x =- 13965 THEN
            sigmoid_f := 2;
        ELSIF x =- 13964 THEN
            sigmoid_f := 2;
        ELSIF x =- 13963 THEN
            sigmoid_f := 2;
        ELSIF x =- 13962 THEN
            sigmoid_f := 2;
        ELSIF x =- 13961 THEN
            sigmoid_f := 2;
        ELSIF x =- 13960 THEN
            sigmoid_f := 2;
        ELSIF x =- 13959 THEN
            sigmoid_f := 2;
        ELSIF x =- 13958 THEN
            sigmoid_f := 2;
        ELSIF x =- 13957 THEN
            sigmoid_f := 2;
        ELSIF x =- 13956 THEN
            sigmoid_f := 2;
        ELSIF x =- 13955 THEN
            sigmoid_f := 2;
        ELSIF x =- 13954 THEN
            sigmoid_f := 2;
        ELSIF x =- 13953 THEN
            sigmoid_f := 2;
        ELSIF x =- 13952 THEN
            sigmoid_f := 2;
        ELSIF x =- 13951 THEN
            sigmoid_f := 2;
        ELSIF x =- 13950 THEN
            sigmoid_f := 2;
        ELSIF x =- 13949 THEN
            sigmoid_f := 2;
        ELSIF x =- 13948 THEN
            sigmoid_f := 2;
        ELSIF x =- 13947 THEN
            sigmoid_f := 2;
        ELSIF x =- 13946 THEN
            sigmoid_f := 2;
        ELSIF x =- 13945 THEN
            sigmoid_f := 2;
        ELSIF x =- 13944 THEN
            sigmoid_f := 2;
        ELSIF x =- 13943 THEN
            sigmoid_f := 2;
        ELSIF x =- 13942 THEN
            sigmoid_f := 2;
        ELSIF x =- 13941 THEN
            sigmoid_f := 2;
        ELSIF x =- 13940 THEN
            sigmoid_f := 2;
        ELSIF x =- 13939 THEN
            sigmoid_f := 2;
        ELSIF x =- 13938 THEN
            sigmoid_f := 2;
        ELSIF x =- 13937 THEN
            sigmoid_f := 2;
        ELSIF x =- 13936 THEN
            sigmoid_f := 2;
        ELSIF x =- 13935 THEN
            sigmoid_f := 2;
        ELSIF x =- 13934 THEN
            sigmoid_f := 2;
        ELSIF x =- 13933 THEN
            sigmoid_f := 2;
        ELSIF x =- 13932 THEN
            sigmoid_f := 2;
        ELSIF x =- 13931 THEN
            sigmoid_f := 2;
        ELSIF x =- 13930 THEN
            sigmoid_f := 2;
        ELSIF x =- 13929 THEN
            sigmoid_f := 2;
        ELSIF x =- 13928 THEN
            sigmoid_f := 2;
        ELSIF x =- 13927 THEN
            sigmoid_f := 2;
        ELSIF x =- 13926 THEN
            sigmoid_f := 2;
        ELSIF x =- 13925 THEN
            sigmoid_f := 2;
        ELSIF x =- 13924 THEN
            sigmoid_f := 2;
        ELSIF x =- 13923 THEN
            sigmoid_f := 2;
        ELSIF x =- 13922 THEN
            sigmoid_f := 2;
        ELSIF x =- 13921 THEN
            sigmoid_f := 2;
        ELSIF x =- 13920 THEN
            sigmoid_f := 2;
        ELSIF x =- 13919 THEN
            sigmoid_f := 2;
        ELSIF x =- 13918 THEN
            sigmoid_f := 2;
        ELSIF x =- 13917 THEN
            sigmoid_f := 2;
        ELSIF x =- 13916 THEN
            sigmoid_f := 2;
        ELSIF x =- 13915 THEN
            sigmoid_f := 2;
        ELSIF x =- 13914 THEN
            sigmoid_f := 2;
        ELSIF x =- 13913 THEN
            sigmoid_f := 2;
        ELSIF x =- 13912 THEN
            sigmoid_f := 2;
        ELSIF x =- 13911 THEN
            sigmoid_f := 2;
        ELSIF x =- 13910 THEN
            sigmoid_f := 2;
        ELSIF x =- 13909 THEN
            sigmoid_f := 2;
        ELSIF x =- 13908 THEN
            sigmoid_f := 2;
        ELSIF x =- 13907 THEN
            sigmoid_f := 2;
        ELSIF x =- 13906 THEN
            sigmoid_f := 2;
        ELSIF x =- 13905 THEN
            sigmoid_f := 2;
        ELSIF x =- 13904 THEN
            sigmoid_f := 2;
        ELSIF x =- 13903 THEN
            sigmoid_f := 2;
        ELSIF x =- 13902 THEN
            sigmoid_f := 2;
        ELSIF x =- 13901 THEN
            sigmoid_f := 2;
        ELSIF x =- 13900 THEN
            sigmoid_f := 2;
        ELSIF x =- 13899 THEN
            sigmoid_f := 2;
        ELSIF x =- 13898 THEN
            sigmoid_f := 2;
        ELSIF x =- 13897 THEN
            sigmoid_f := 2;
        ELSIF x =- 13896 THEN
            sigmoid_f := 2;
        ELSIF x =- 13895 THEN
            sigmoid_f := 2;
        ELSIF x =- 13894 THEN
            sigmoid_f := 2;
        ELSIF x =- 13893 THEN
            sigmoid_f := 2;
        ELSIF x =- 13892 THEN
            sigmoid_f := 2;
        ELSIF x =- 13891 THEN
            sigmoid_f := 2;
        ELSIF x =- 13890 THEN
            sigmoid_f := 2;
        ELSIF x =- 13889 THEN
            sigmoid_f := 2;
        ELSIF x =- 13888 THEN
            sigmoid_f := 2;
        ELSIF x =- 13887 THEN
            sigmoid_f := 2;
        ELSIF x =- 13886 THEN
            sigmoid_f := 2;
        ELSIF x =- 13885 THEN
            sigmoid_f := 2;
        ELSIF x =- 13884 THEN
            sigmoid_f := 2;
        ELSIF x =- 13883 THEN
            sigmoid_f := 2;
        ELSIF x =- 13882 THEN
            sigmoid_f := 2;
        ELSIF x =- 13881 THEN
            sigmoid_f := 2;
        ELSIF x =- 13880 THEN
            sigmoid_f := 2;
        ELSIF x =- 13879 THEN
            sigmoid_f := 2;
        ELSIF x =- 13878 THEN
            sigmoid_f := 2;
        ELSIF x =- 13877 THEN
            sigmoid_f := 2;
        ELSIF x =- 13876 THEN
            sigmoid_f := 2;
        ELSIF x =- 13875 THEN
            sigmoid_f := 2;
        ELSIF x =- 13874 THEN
            sigmoid_f := 2;
        ELSIF x =- 13873 THEN
            sigmoid_f := 2;
        ELSIF x =- 13872 THEN
            sigmoid_f := 2;
        ELSIF x =- 13871 THEN
            sigmoid_f := 2;
        ELSIF x =- 13870 THEN
            sigmoid_f := 2;
        ELSIF x =- 13869 THEN
            sigmoid_f := 2;
        ELSIF x =- 13868 THEN
            sigmoid_f := 2;
        ELSIF x =- 13867 THEN
            sigmoid_f := 2;
        ELSIF x =- 13866 THEN
            sigmoid_f := 2;
        ELSIF x =- 13865 THEN
            sigmoid_f := 2;
        ELSIF x =- 13864 THEN
            sigmoid_f := 2;
        ELSIF x =- 13863 THEN
            sigmoid_f := 2;
        ELSIF x =- 13862 THEN
            sigmoid_f := 2;
        ELSIF x =- 13861 THEN
            sigmoid_f := 2;
        ELSIF x =- 13860 THEN
            sigmoid_f := 2;
        ELSIF x =- 13859 THEN
            sigmoid_f := 2;
        ELSIF x =- 13858 THEN
            sigmoid_f := 2;
        ELSIF x =- 13857 THEN
            sigmoid_f := 2;
        ELSIF x =- 13856 THEN
            sigmoid_f := 2;
        ELSIF x =- 13855 THEN
            sigmoid_f := 2;
        ELSIF x =- 13854 THEN
            sigmoid_f := 2;
        ELSIF x =- 13853 THEN
            sigmoid_f := 2;
        ELSIF x =- 13852 THEN
            sigmoid_f := 2;
        ELSIF x =- 13851 THEN
            sigmoid_f := 2;
        ELSIF x =- 13850 THEN
            sigmoid_f := 2;
        ELSIF x =- 13849 THEN
            sigmoid_f := 2;
        ELSIF x =- 13848 THEN
            sigmoid_f := 2;
        ELSIF x =- 13847 THEN
            sigmoid_f := 2;
        ELSIF x =- 13846 THEN
            sigmoid_f := 2;
        ELSIF x =- 13845 THEN
            sigmoid_f := 2;
        ELSIF x =- 13844 THEN
            sigmoid_f := 2;
        ELSIF x =- 13843 THEN
            sigmoid_f := 2;
        ELSIF x =- 13842 THEN
            sigmoid_f := 2;
        ELSIF x =- 13841 THEN
            sigmoid_f := 2;
        ELSIF x =- 13840 THEN
            sigmoid_f := 2;
        ELSIF x =- 13839 THEN
            sigmoid_f := 2;
        ELSIF x =- 13838 THEN
            sigmoid_f := 2;
        ELSIF x =- 13837 THEN
            sigmoid_f := 2;
        ELSIF x =- 13836 THEN
            sigmoid_f := 2;
        ELSIF x =- 13835 THEN
            sigmoid_f := 2;
        ELSIF x =- 13834 THEN
            sigmoid_f := 2;
        ELSIF x =- 13833 THEN
            sigmoid_f := 2;
        ELSIF x =- 13832 THEN
            sigmoid_f := 2;
        ELSIF x =- 13831 THEN
            sigmoid_f := 2;
        ELSIF x =- 13830 THEN
            sigmoid_f := 2;
        ELSIF x =- 13829 THEN
            sigmoid_f := 2;
        ELSIF x =- 13828 THEN
            sigmoid_f := 2;
        ELSIF x =- 13827 THEN
            sigmoid_f := 2;
        ELSIF x =- 13826 THEN
            sigmoid_f := 2;
        ELSIF x =- 13825 THEN
            sigmoid_f := 2;
        ELSIF x =- 13824 THEN
            sigmoid_f := 2;
        ELSIF x =- 13823 THEN
            sigmoid_f := 3;
        ELSIF x =- 13822 THEN
            sigmoid_f := 3;
        ELSIF x =- 13821 THEN
            sigmoid_f := 3;
        ELSIF x =- 13820 THEN
            sigmoid_f := 3;
        ELSIF x =- 13819 THEN
            sigmoid_f := 3;
        ELSIF x =- 13818 THEN
            sigmoid_f := 3;
        ELSIF x =- 13817 THEN
            sigmoid_f := 3;
        ELSIF x =- 13816 THEN
            sigmoid_f := 3;
        ELSIF x =- 13815 THEN
            sigmoid_f := 3;
        ELSIF x =- 13814 THEN
            sigmoid_f := 3;
        ELSIF x =- 13813 THEN
            sigmoid_f := 3;
        ELSIF x =- 13812 THEN
            sigmoid_f := 3;
        ELSIF x =- 13811 THEN
            sigmoid_f := 3;
        ELSIF x =- 13810 THEN
            sigmoid_f := 3;
        ELSIF x =- 13809 THEN
            sigmoid_f := 3;
        ELSIF x =- 13808 THEN
            sigmoid_f := 3;
        ELSIF x =- 13807 THEN
            sigmoid_f := 3;
        ELSIF x =- 13806 THEN
            sigmoid_f := 3;
        ELSIF x =- 13805 THEN
            sigmoid_f := 3;
        ELSIF x =- 13804 THEN
            sigmoid_f := 3;
        ELSIF x =- 13803 THEN
            sigmoid_f := 3;
        ELSIF x =- 13802 THEN
            sigmoid_f := 3;
        ELSIF x =- 13801 THEN
            sigmoid_f := 3;
        ELSIF x =- 13800 THEN
            sigmoid_f := 3;
        ELSIF x =- 13799 THEN
            sigmoid_f := 3;
        ELSIF x =- 13798 THEN
            sigmoid_f := 3;
        ELSIF x =- 13797 THEN
            sigmoid_f := 3;
        ELSIF x =- 13796 THEN
            sigmoid_f := 3;
        ELSIF x =- 13795 THEN
            sigmoid_f := 3;
        ELSIF x =- 13794 THEN
            sigmoid_f := 3;
        ELSIF x =- 13793 THEN
            sigmoid_f := 3;
        ELSIF x =- 13792 THEN
            sigmoid_f := 3;
        ELSIF x =- 13791 THEN
            sigmoid_f := 3;
        ELSIF x =- 13790 THEN
            sigmoid_f := 3;
        ELSIF x =- 13789 THEN
            sigmoid_f := 3;
        ELSIF x =- 13788 THEN
            sigmoid_f := 3;
        ELSIF x =- 13787 THEN
            sigmoid_f := 3;
        ELSIF x =- 13786 THEN
            sigmoid_f := 3;
        ELSIF x =- 13785 THEN
            sigmoid_f := 3;
        ELSIF x =- 13784 THEN
            sigmoid_f := 3;
        ELSIF x =- 13783 THEN
            sigmoid_f := 3;
        ELSIF x =- 13782 THEN
            sigmoid_f := 3;
        ELSIF x =- 13781 THEN
            sigmoid_f := 3;
        ELSIF x =- 13780 THEN
            sigmoid_f := 3;
        ELSIF x =- 13779 THEN
            sigmoid_f := 3;
        ELSIF x =- 13778 THEN
            sigmoid_f := 3;
        ELSIF x =- 13777 THEN
            sigmoid_f := 3;
        ELSIF x =- 13776 THEN
            sigmoid_f := 3;
        ELSIF x =- 13775 THEN
            sigmoid_f := 3;
        ELSIF x =- 13774 THEN
            sigmoid_f := 3;
        ELSIF x =- 13773 THEN
            sigmoid_f := 3;
        ELSIF x =- 13772 THEN
            sigmoid_f := 3;
        ELSIF x =- 13771 THEN
            sigmoid_f := 3;
        ELSIF x =- 13770 THEN
            sigmoid_f := 3;
        ELSIF x =- 13769 THEN
            sigmoid_f := 3;
        ELSIF x =- 13768 THEN
            sigmoid_f := 3;
        ELSIF x =- 13767 THEN
            sigmoid_f := 3;
        ELSIF x =- 13766 THEN
            sigmoid_f := 3;
        ELSIF x =- 13765 THEN
            sigmoid_f := 3;
        ELSIF x =- 13764 THEN
            sigmoid_f := 3;
        ELSIF x =- 13763 THEN
            sigmoid_f := 3;
        ELSIF x =- 13762 THEN
            sigmoid_f := 3;
        ELSIF x =- 13761 THEN
            sigmoid_f := 3;
        ELSIF x =- 13760 THEN
            sigmoid_f := 3;
        ELSIF x =- 13759 THEN
            sigmoid_f := 3;
        ELSIF x =- 13758 THEN
            sigmoid_f := 3;
        ELSIF x =- 13757 THEN
            sigmoid_f := 3;
        ELSIF x =- 13756 THEN
            sigmoid_f := 3;
        ELSIF x =- 13755 THEN
            sigmoid_f := 3;
        ELSIF x =- 13754 THEN
            sigmoid_f := 3;
        ELSIF x =- 13753 THEN
            sigmoid_f := 3;
        ELSIF x =- 13752 THEN
            sigmoid_f := 3;
        ELSIF x =- 13751 THEN
            sigmoid_f := 3;
        ELSIF x =- 13750 THEN
            sigmoid_f := 3;
        ELSIF x =- 13749 THEN
            sigmoid_f := 3;
        ELSIF x =- 13748 THEN
            sigmoid_f := 3;
        ELSIF x =- 13747 THEN
            sigmoid_f := 3;
        ELSIF x =- 13746 THEN
            sigmoid_f := 3;
        ELSIF x =- 13745 THEN
            sigmoid_f := 3;
        ELSIF x =- 13744 THEN
            sigmoid_f := 3;
        ELSIF x =- 13743 THEN
            sigmoid_f := 3;
        ELSIF x =- 13742 THEN
            sigmoid_f := 3;
        ELSIF x =- 13741 THEN
            sigmoid_f := 3;
        ELSIF x =- 13740 THEN
            sigmoid_f := 3;
        ELSIF x =- 13739 THEN
            sigmoid_f := 3;
        ELSIF x =- 13738 THEN
            sigmoid_f := 3;
        ELSIF x =- 13737 THEN
            sigmoid_f := 3;
        ELSIF x =- 13736 THEN
            sigmoid_f := 3;
        ELSIF x =- 13735 THEN
            sigmoid_f := 3;
        ELSIF x =- 13734 THEN
            sigmoid_f := 3;
        ELSIF x =- 13733 THEN
            sigmoid_f := 3;
        ELSIF x =- 13732 THEN
            sigmoid_f := 3;
        ELSIF x =- 13731 THEN
            sigmoid_f := 3;
        ELSIF x =- 13730 THEN
            sigmoid_f := 3;
        ELSIF x =- 13729 THEN
            sigmoid_f := 3;
        ELSIF x =- 13728 THEN
            sigmoid_f := 3;
        ELSIF x =- 13727 THEN
            sigmoid_f := 3;
        ELSIF x =- 13726 THEN
            sigmoid_f := 3;
        ELSIF x =- 13725 THEN
            sigmoid_f := 3;
        ELSIF x =- 13724 THEN
            sigmoid_f := 3;
        ELSIF x =- 13723 THEN
            sigmoid_f := 3;
        ELSIF x =- 13722 THEN
            sigmoid_f := 3;
        ELSIF x =- 13721 THEN
            sigmoid_f := 3;
        ELSIF x =- 13720 THEN
            sigmoid_f := 3;
        ELSIF x =- 13719 THEN
            sigmoid_f := 3;
        ELSIF x =- 13718 THEN
            sigmoid_f := 3;
        ELSIF x =- 13717 THEN
            sigmoid_f := 3;
        ELSIF x =- 13716 THEN
            sigmoid_f := 3;
        ELSIF x =- 13715 THEN
            sigmoid_f := 3;
        ELSIF x =- 13714 THEN
            sigmoid_f := 3;
        ELSIF x =- 13713 THEN
            sigmoid_f := 3;
        ELSIF x =- 13712 THEN
            sigmoid_f := 3;
        ELSIF x =- 13711 THEN
            sigmoid_f := 3;
        ELSIF x =- 13710 THEN
            sigmoid_f := 3;
        ELSIF x =- 13709 THEN
            sigmoid_f := 3;
        ELSIF x =- 13708 THEN
            sigmoid_f := 3;
        ELSIF x =- 13707 THEN
            sigmoid_f := 3;
        ELSIF x =- 13706 THEN
            sigmoid_f := 3;
        ELSIF x =- 13705 THEN
            sigmoid_f := 3;
        ELSIF x =- 13704 THEN
            sigmoid_f := 3;
        ELSIF x =- 13703 THEN
            sigmoid_f := 3;
        ELSIF x =- 13702 THEN
            sigmoid_f := 3;
        ELSIF x =- 13701 THEN
            sigmoid_f := 3;
        ELSIF x =- 13700 THEN
            sigmoid_f := 3;
        ELSIF x =- 13699 THEN
            sigmoid_f := 3;
        ELSIF x =- 13698 THEN
            sigmoid_f := 3;
        ELSIF x =- 13697 THEN
            sigmoid_f := 3;
        ELSIF x =- 13696 THEN
            sigmoid_f := 3;
        ELSIF x =- 13695 THEN
            sigmoid_f := 3;
        ELSIF x =- 13694 THEN
            sigmoid_f := 3;
        ELSIF x =- 13693 THEN
            sigmoid_f := 3;
        ELSIF x =- 13692 THEN
            sigmoid_f := 3;
        ELSIF x =- 13691 THEN
            sigmoid_f := 3;
        ELSIF x =- 13690 THEN
            sigmoid_f := 3;
        ELSIF x =- 13689 THEN
            sigmoid_f := 3;
        ELSIF x =- 13688 THEN
            sigmoid_f := 3;
        ELSIF x =- 13687 THEN
            sigmoid_f := 3;
        ELSIF x =- 13686 THEN
            sigmoid_f := 3;
        ELSIF x =- 13685 THEN
            sigmoid_f := 3;
        ELSIF x =- 13684 THEN
            sigmoid_f := 3;
        ELSIF x =- 13683 THEN
            sigmoid_f := 3;
        ELSIF x =- 13682 THEN
            sigmoid_f := 3;
        ELSIF x =- 13681 THEN
            sigmoid_f := 3;
        ELSIF x =- 13680 THEN
            sigmoid_f := 3;
        ELSIF x =- 13679 THEN
            sigmoid_f := 3;
        ELSIF x =- 13678 THEN
            sigmoid_f := 3;
        ELSIF x =- 13677 THEN
            sigmoid_f := 3;
        ELSIF x =- 13676 THEN
            sigmoid_f := 3;
        ELSIF x =- 13675 THEN
            sigmoid_f := 3;
        ELSIF x =- 13674 THEN
            sigmoid_f := 3;
        ELSIF x =- 13673 THEN
            sigmoid_f := 3;
        ELSIF x =- 13672 THEN
            sigmoid_f := 3;
        ELSIF x =- 13671 THEN
            sigmoid_f := 3;
        ELSIF x =- 13670 THEN
            sigmoid_f := 3;
        ELSIF x =- 13669 THEN
            sigmoid_f := 3;
        ELSIF x =- 13668 THEN
            sigmoid_f := 3;
        ELSIF x =- 13667 THEN
            sigmoid_f := 3;
        ELSIF x =- 13666 THEN
            sigmoid_f := 3;
        ELSIF x =- 13665 THEN
            sigmoid_f := 3;
        ELSIF x =- 13664 THEN
            sigmoid_f := 3;
        ELSIF x =- 13663 THEN
            sigmoid_f := 3;
        ELSIF x =- 13662 THEN
            sigmoid_f := 3;
        ELSIF x =- 13661 THEN
            sigmoid_f := 3;
        ELSIF x =- 13660 THEN
            sigmoid_f := 3;
        ELSIF x =- 13659 THEN
            sigmoid_f := 3;
        ELSIF x =- 13658 THEN
            sigmoid_f := 3;
        ELSIF x =- 13657 THEN
            sigmoid_f := 3;
        ELSIF x =- 13656 THEN
            sigmoid_f := 3;
        ELSIF x =- 13655 THEN
            sigmoid_f := 3;
        ELSIF x =- 13654 THEN
            sigmoid_f := 3;
        ELSIF x =- 13653 THEN
            sigmoid_f := 3;
        ELSIF x =- 13652 THEN
            sigmoid_f := 3;
        ELSIF x =- 13651 THEN
            sigmoid_f := 3;
        ELSIF x =- 13650 THEN
            sigmoid_f := 3;
        ELSIF x =- 13649 THEN
            sigmoid_f := 3;
        ELSIF x =- 13648 THEN
            sigmoid_f := 3;
        ELSIF x =- 13647 THEN
            sigmoid_f := 3;
        ELSIF x =- 13646 THEN
            sigmoid_f := 3;
        ELSIF x =- 13645 THEN
            sigmoid_f := 3;
        ELSIF x =- 13644 THEN
            sigmoid_f := 3;
        ELSIF x =- 13643 THEN
            sigmoid_f := 3;
        ELSIF x =- 13642 THEN
            sigmoid_f := 3;
        ELSIF x =- 13641 THEN
            sigmoid_f := 3;
        ELSIF x =- 13640 THEN
            sigmoid_f := 3;
        ELSIF x =- 13639 THEN
            sigmoid_f := 3;
        ELSIF x =- 13638 THEN
            sigmoid_f := 3;
        ELSIF x =- 13637 THEN
            sigmoid_f := 3;
        ELSIF x =- 13636 THEN
            sigmoid_f := 3;
        ELSIF x =- 13635 THEN
            sigmoid_f := 3;
        ELSIF x =- 13634 THEN
            sigmoid_f := 3;
        ELSIF x =- 13633 THEN
            sigmoid_f := 3;
        ELSIF x =- 13632 THEN
            sigmoid_f := 3;
        ELSIF x =- 13631 THEN
            sigmoid_f := 3;
        ELSIF x =- 13630 THEN
            sigmoid_f := 3;
        ELSIF x =- 13629 THEN
            sigmoid_f := 3;
        ELSIF x =- 13628 THEN
            sigmoid_f := 3;
        ELSIF x =- 13627 THEN
            sigmoid_f := 3;
        ELSIF x =- 13626 THEN
            sigmoid_f := 3;
        ELSIF x =- 13625 THEN
            sigmoid_f := 3;
        ELSIF x =- 13624 THEN
            sigmoid_f := 3;
        ELSIF x =- 13623 THEN
            sigmoid_f := 3;
        ELSIF x =- 13622 THEN
            sigmoid_f := 3;
        ELSIF x =- 13621 THEN
            sigmoid_f := 3;
        ELSIF x =- 13620 THEN
            sigmoid_f := 3;
        ELSIF x =- 13619 THEN
            sigmoid_f := 3;
        ELSIF x =- 13618 THEN
            sigmoid_f := 3;
        ELSIF x =- 13617 THEN
            sigmoid_f := 3;
        ELSIF x =- 13616 THEN
            sigmoid_f := 3;
        ELSIF x =- 13615 THEN
            sigmoid_f := 3;
        ELSIF x =- 13614 THEN
            sigmoid_f := 3;
        ELSIF x =- 13613 THEN
            sigmoid_f := 3;
        ELSIF x =- 13612 THEN
            sigmoid_f := 3;
        ELSIF x =- 13611 THEN
            sigmoid_f := 3;
        ELSIF x =- 13610 THEN
            sigmoid_f := 3;
        ELSIF x =- 13609 THEN
            sigmoid_f := 3;
        ELSIF x =- 13608 THEN
            sigmoid_f := 3;
        ELSIF x =- 13607 THEN
            sigmoid_f := 3;
        ELSIF x =- 13606 THEN
            sigmoid_f := 3;
        ELSIF x =- 13605 THEN
            sigmoid_f := 3;
        ELSIF x =- 13604 THEN
            sigmoid_f := 3;
        ELSIF x =- 13603 THEN
            sigmoid_f := 3;
        ELSIF x =- 13602 THEN
            sigmoid_f := 3;
        ELSIF x =- 13601 THEN
            sigmoid_f := 3;
        ELSIF x =- 13600 THEN
            sigmoid_f := 3;
        ELSIF x =- 13599 THEN
            sigmoid_f := 3;
        ELSIF x =- 13598 THEN
            sigmoid_f := 3;
        ELSIF x =- 13597 THEN
            sigmoid_f := 3;
        ELSIF x =- 13596 THEN
            sigmoid_f := 3;
        ELSIF x =- 13595 THEN
            sigmoid_f := 3;
        ELSIF x =- 13594 THEN
            sigmoid_f := 3;
        ELSIF x =- 13593 THEN
            sigmoid_f := 3;
        ELSIF x =- 13592 THEN
            sigmoid_f := 3;
        ELSIF x =- 13591 THEN
            sigmoid_f := 3;
        ELSIF x =- 13590 THEN
            sigmoid_f := 3;
        ELSIF x =- 13589 THEN
            sigmoid_f := 3;
        ELSIF x =- 13588 THEN
            sigmoid_f := 3;
        ELSIF x =- 13587 THEN
            sigmoid_f := 3;
        ELSIF x =- 13586 THEN
            sigmoid_f := 3;
        ELSIF x =- 13585 THEN
            sigmoid_f := 3;
        ELSIF x =- 13584 THEN
            sigmoid_f := 3;
        ELSIF x =- 13583 THEN
            sigmoid_f := 3;
        ELSIF x =- 13582 THEN
            sigmoid_f := 3;
        ELSIF x =- 13581 THEN
            sigmoid_f := 3;
        ELSIF x =- 13580 THEN
            sigmoid_f := 3;
        ELSIF x =- 13579 THEN
            sigmoid_f := 3;
        ELSIF x =- 13578 THEN
            sigmoid_f := 3;
        ELSIF x =- 13577 THEN
            sigmoid_f := 3;
        ELSIF x =- 13576 THEN
            sigmoid_f := 3;
        ELSIF x =- 13575 THEN
            sigmoid_f := 3;
        ELSIF x =- 13574 THEN
            sigmoid_f := 3;
        ELSIF x =- 13573 THEN
            sigmoid_f := 3;
        ELSIF x =- 13572 THEN
            sigmoid_f := 3;
        ELSIF x =- 13571 THEN
            sigmoid_f := 3;
        ELSIF x =- 13570 THEN
            sigmoid_f := 3;
        ELSIF x =- 13569 THEN
            sigmoid_f := 3;
        ELSIF x =- 13568 THEN
            sigmoid_f := 3;
        ELSIF x =- 13567 THEN
            sigmoid_f := 3;
        ELSIF x =- 13566 THEN
            sigmoid_f := 3;
        ELSIF x =- 13565 THEN
            sigmoid_f := 3;
        ELSIF x =- 13564 THEN
            sigmoid_f := 3;
        ELSIF x =- 13563 THEN
            sigmoid_f := 3;
        ELSIF x =- 13562 THEN
            sigmoid_f := 3;
        ELSIF x =- 13561 THEN
            sigmoid_f := 3;
        ELSIF x =- 13560 THEN
            sigmoid_f := 3;
        ELSIF x =- 13559 THEN
            sigmoid_f := 3;
        ELSIF x =- 13558 THEN
            sigmoid_f := 3;
        ELSIF x =- 13557 THEN
            sigmoid_f := 3;
        ELSIF x =- 13556 THEN
            sigmoid_f := 3;
        ELSIF x =- 13555 THEN
            sigmoid_f := 3;
        ELSIF x =- 13554 THEN
            sigmoid_f := 3;
        ELSIF x =- 13553 THEN
            sigmoid_f := 3;
        ELSIF x =- 13552 THEN
            sigmoid_f := 3;
        ELSIF x =- 13551 THEN
            sigmoid_f := 3;
        ELSIF x =- 13550 THEN
            sigmoid_f := 3;
        ELSIF x =- 13549 THEN
            sigmoid_f := 3;
        ELSIF x =- 13548 THEN
            sigmoid_f := 3;
        ELSIF x =- 13547 THEN
            sigmoid_f := 3;
        ELSIF x =- 13546 THEN
            sigmoid_f := 3;
        ELSIF x =- 13545 THEN
            sigmoid_f := 3;
        ELSIF x =- 13544 THEN
            sigmoid_f := 3;
        ELSIF x =- 13543 THEN
            sigmoid_f := 3;
        ELSIF x =- 13542 THEN
            sigmoid_f := 3;
        ELSIF x =- 13541 THEN
            sigmoid_f := 3;
        ELSIF x =- 13540 THEN
            sigmoid_f := 3;
        ELSIF x =- 13539 THEN
            sigmoid_f := 3;
        ELSIF x =- 13538 THEN
            sigmoid_f := 3;
        ELSIF x =- 13537 THEN
            sigmoid_f := 3;
        ELSIF x =- 13536 THEN
            sigmoid_f := 3;
        ELSIF x =- 13535 THEN
            sigmoid_f := 3;
        ELSIF x =- 13534 THEN
            sigmoid_f := 3;
        ELSIF x =- 13533 THEN
            sigmoid_f := 3;
        ELSIF x =- 13532 THEN
            sigmoid_f := 3;
        ELSIF x =- 13531 THEN
            sigmoid_f := 3;
        ELSIF x =- 13530 THEN
            sigmoid_f := 3;
        ELSIF x =- 13529 THEN
            sigmoid_f := 3;
        ELSIF x =- 13528 THEN
            sigmoid_f := 3;
        ELSIF x =- 13527 THEN
            sigmoid_f := 3;
        ELSIF x =- 13526 THEN
            sigmoid_f := 3;
        ELSIF x =- 13525 THEN
            sigmoid_f := 3;
        ELSIF x =- 13524 THEN
            sigmoid_f := 3;
        ELSIF x =- 13523 THEN
            sigmoid_f := 3;
        ELSIF x =- 13522 THEN
            sigmoid_f := 3;
        ELSIF x =- 13521 THEN
            sigmoid_f := 3;
        ELSIF x =- 13520 THEN
            sigmoid_f := 3;
        ELSIF x =- 13519 THEN
            sigmoid_f := 3;
        ELSIF x =- 13518 THEN
            sigmoid_f := 3;
        ELSIF x =- 13517 THEN
            sigmoid_f := 3;
        ELSIF x =- 13516 THEN
            sigmoid_f := 3;
        ELSIF x =- 13515 THEN
            sigmoid_f := 3;
        ELSIF x =- 13514 THEN
            sigmoid_f := 3;
        ELSIF x =- 13513 THEN
            sigmoid_f := 3;
        ELSIF x =- 13512 THEN
            sigmoid_f := 3;
        ELSIF x =- 13511 THEN
            sigmoid_f := 3;
        ELSIF x =- 13510 THEN
            sigmoid_f := 3;
        ELSIF x =- 13509 THEN
            sigmoid_f := 3;
        ELSIF x =- 13508 THEN
            sigmoid_f := 3;
        ELSIF x =- 13507 THEN
            sigmoid_f := 3;
        ELSIF x =- 13506 THEN
            sigmoid_f := 3;
        ELSIF x =- 13505 THEN
            sigmoid_f := 3;
        ELSIF x =- 13504 THEN
            sigmoid_f := 3;
        ELSIF x =- 13503 THEN
            sigmoid_f := 3;
        ELSIF x =- 13502 THEN
            sigmoid_f := 3;
        ELSIF x =- 13501 THEN
            sigmoid_f := 3;
        ELSIF x =- 13500 THEN
            sigmoid_f := 3;
        ELSIF x =- 13499 THEN
            sigmoid_f := 3;
        ELSIF x =- 13498 THEN
            sigmoid_f := 3;
        ELSIF x =- 13497 THEN
            sigmoid_f := 3;
        ELSIF x =- 13496 THEN
            sigmoid_f := 3;
        ELSIF x =- 13495 THEN
            sigmoid_f := 3;
        ELSIF x =- 13494 THEN
            sigmoid_f := 3;
        ELSIF x =- 13493 THEN
            sigmoid_f := 3;
        ELSIF x =- 13492 THEN
            sigmoid_f := 3;
        ELSIF x =- 13491 THEN
            sigmoid_f := 3;
        ELSIF x =- 13490 THEN
            sigmoid_f := 3;
        ELSIF x =- 13489 THEN
            sigmoid_f := 3;
        ELSIF x =- 13488 THEN
            sigmoid_f := 3;
        ELSIF x =- 13487 THEN
            sigmoid_f := 3;
        ELSIF x =- 13486 THEN
            sigmoid_f := 3;
        ELSIF x =- 13485 THEN
            sigmoid_f := 3;
        ELSIF x =- 13484 THEN
            sigmoid_f := 3;
        ELSIF x =- 13483 THEN
            sigmoid_f := 3;
        ELSIF x =- 13482 THEN
            sigmoid_f := 3;
        ELSIF x =- 13481 THEN
            sigmoid_f := 3;
        ELSIF x =- 13480 THEN
            sigmoid_f := 3;
        ELSIF x =- 13479 THEN
            sigmoid_f := 3;
        ELSIF x =- 13478 THEN
            sigmoid_f := 3;
        ELSIF x =- 13477 THEN
            sigmoid_f := 3;
        ELSIF x =- 13476 THEN
            sigmoid_f := 3;
        ELSIF x =- 13475 THEN
            sigmoid_f := 3;
        ELSIF x =- 13474 THEN
            sigmoid_f := 3;
        ELSIF x =- 13473 THEN
            sigmoid_f := 3;
        ELSIF x =- 13472 THEN
            sigmoid_f := 3;
        ELSIF x =- 13471 THEN
            sigmoid_f := 3;
        ELSIF x =- 13470 THEN
            sigmoid_f := 3;
        ELSIF x =- 13469 THEN
            sigmoid_f := 3;
        ELSIF x =- 13468 THEN
            sigmoid_f := 3;
        ELSIF x =- 13467 THEN
            sigmoid_f := 3;
        ELSIF x =- 13466 THEN
            sigmoid_f := 3;
        ELSIF x =- 13465 THEN
            sigmoid_f := 3;
        ELSIF x =- 13464 THEN
            sigmoid_f := 3;
        ELSIF x =- 13463 THEN
            sigmoid_f := 3;
        ELSIF x =- 13462 THEN
            sigmoid_f := 3;
        ELSIF x =- 13461 THEN
            sigmoid_f := 3;
        ELSIF x =- 13460 THEN
            sigmoid_f := 3;
        ELSIF x =- 13459 THEN
            sigmoid_f := 3;
        ELSIF x =- 13458 THEN
            sigmoid_f := 3;
        ELSIF x =- 13457 THEN
            sigmoid_f := 3;
        ELSIF x =- 13456 THEN
            sigmoid_f := 3;
        ELSIF x =- 13455 THEN
            sigmoid_f := 3;
        ELSIF x =- 13454 THEN
            sigmoid_f := 3;
        ELSIF x =- 13453 THEN
            sigmoid_f := 3;
        ELSIF x =- 13452 THEN
            sigmoid_f := 3;
        ELSIF x =- 13451 THEN
            sigmoid_f := 3;
        ELSIF x =- 13450 THEN
            sigmoid_f := 3;
        ELSIF x =- 13449 THEN
            sigmoid_f := 3;
        ELSIF x =- 13448 THEN
            sigmoid_f := 3;
        ELSIF x =- 13447 THEN
            sigmoid_f := 3;
        ELSIF x =- 13446 THEN
            sigmoid_f := 3;
        ELSIF x =- 13445 THEN
            sigmoid_f := 3;
        ELSIF x =- 13444 THEN
            sigmoid_f := 3;
        ELSIF x =- 13443 THEN
            sigmoid_f := 3;
        ELSIF x =- 13442 THEN
            sigmoid_f := 3;
        ELSIF x =- 13441 THEN
            sigmoid_f := 3;
        ELSIF x =- 13440 THEN
            sigmoid_f := 3;
        ELSIF x =- 13439 THEN
            sigmoid_f := 3;
        ELSIF x =- 13438 THEN
            sigmoid_f := 3;
        ELSIF x =- 13437 THEN
            sigmoid_f := 3;
        ELSIF x =- 13436 THEN
            sigmoid_f := 3;
        ELSIF x =- 13435 THEN
            sigmoid_f := 3;
        ELSIF x =- 13434 THEN
            sigmoid_f := 3;
        ELSIF x =- 13433 THEN
            sigmoid_f := 3;
        ELSIF x =- 13432 THEN
            sigmoid_f := 3;
        ELSIF x =- 13431 THEN
            sigmoid_f := 3;
        ELSIF x =- 13430 THEN
            sigmoid_f := 3;
        ELSIF x =- 13429 THEN
            sigmoid_f := 3;
        ELSIF x =- 13428 THEN
            sigmoid_f := 3;
        ELSIF x =- 13427 THEN
            sigmoid_f := 3;
        ELSIF x =- 13426 THEN
            sigmoid_f := 3;
        ELSIF x =- 13425 THEN
            sigmoid_f := 3;
        ELSIF x =- 13424 THEN
            sigmoid_f := 3;
        ELSIF x =- 13423 THEN
            sigmoid_f := 3;
        ELSIF x =- 13422 THEN
            sigmoid_f := 3;
        ELSIF x =- 13421 THEN
            sigmoid_f := 3;
        ELSIF x =- 13420 THEN
            sigmoid_f := 3;
        ELSIF x =- 13419 THEN
            sigmoid_f := 3;
        ELSIF x =- 13418 THEN
            sigmoid_f := 3;
        ELSIF x =- 13417 THEN
            sigmoid_f := 3;
        ELSIF x =- 13416 THEN
            sigmoid_f := 3;
        ELSIF x =- 13415 THEN
            sigmoid_f := 3;
        ELSIF x =- 13414 THEN
            sigmoid_f := 3;
        ELSIF x =- 13413 THEN
            sigmoid_f := 3;
        ELSIF x =- 13412 THEN
            sigmoid_f := 3;
        ELSIF x =- 13411 THEN
            sigmoid_f := 3;
        ELSIF x =- 13410 THEN
            sigmoid_f := 3;
        ELSIF x =- 13409 THEN
            sigmoid_f := 3;
        ELSIF x =- 13408 THEN
            sigmoid_f := 3;
        ELSIF x =- 13407 THEN
            sigmoid_f := 3;
        ELSIF x =- 13406 THEN
            sigmoid_f := 3;
        ELSIF x =- 13405 THEN
            sigmoid_f := 3;
        ELSIF x =- 13404 THEN
            sigmoid_f := 3;
        ELSIF x =- 13403 THEN
            sigmoid_f := 3;
        ELSIF x =- 13402 THEN
            sigmoid_f := 3;
        ELSIF x =- 13401 THEN
            sigmoid_f := 3;
        ELSIF x =- 13400 THEN
            sigmoid_f := 3;
        ELSIF x =- 13399 THEN
            sigmoid_f := 3;
        ELSIF x =- 13398 THEN
            sigmoid_f := 3;
        ELSIF x =- 13397 THEN
            sigmoid_f := 3;
        ELSIF x =- 13396 THEN
            sigmoid_f := 3;
        ELSIF x =- 13395 THEN
            sigmoid_f := 3;
        ELSIF x =- 13394 THEN
            sigmoid_f := 3;
        ELSIF x =- 13393 THEN
            sigmoid_f := 3;
        ELSIF x =- 13392 THEN
            sigmoid_f := 3;
        ELSIF x =- 13391 THEN
            sigmoid_f := 3;
        ELSIF x =- 13390 THEN
            sigmoid_f := 3;
        ELSIF x =- 13389 THEN
            sigmoid_f := 3;
        ELSIF x =- 13388 THEN
            sigmoid_f := 3;
        ELSIF x =- 13387 THEN
            sigmoid_f := 3;
        ELSIF x =- 13386 THEN
            sigmoid_f := 3;
        ELSIF x =- 13385 THEN
            sigmoid_f := 3;
        ELSIF x =- 13384 THEN
            sigmoid_f := 3;
        ELSIF x =- 13383 THEN
            sigmoid_f := 3;
        ELSIF x =- 13382 THEN
            sigmoid_f := 3;
        ELSIF x =- 13381 THEN
            sigmoid_f := 3;
        ELSIF x =- 13380 THEN
            sigmoid_f := 3;
        ELSIF x =- 13379 THEN
            sigmoid_f := 3;
        ELSIF x =- 13378 THEN
            sigmoid_f := 3;
        ELSIF x =- 13377 THEN
            sigmoid_f := 3;
        ELSIF x =- 13376 THEN
            sigmoid_f := 3;
        ELSIF x =- 13375 THEN
            sigmoid_f := 3;
        ELSIF x =- 13374 THEN
            sigmoid_f := 3;
        ELSIF x =- 13373 THEN
            sigmoid_f := 3;
        ELSIF x =- 13372 THEN
            sigmoid_f := 3;
        ELSIF x =- 13371 THEN
            sigmoid_f := 3;
        ELSIF x =- 13370 THEN
            sigmoid_f := 3;
        ELSIF x =- 13369 THEN
            sigmoid_f := 3;
        ELSIF x =- 13368 THEN
            sigmoid_f := 3;
        ELSIF x =- 13367 THEN
            sigmoid_f := 3;
        ELSIF x =- 13366 THEN
            sigmoid_f := 3;
        ELSIF x =- 13365 THEN
            sigmoid_f := 3;
        ELSIF x =- 13364 THEN
            sigmoid_f := 3;
        ELSIF x =- 13363 THEN
            sigmoid_f := 3;
        ELSIF x =- 13362 THEN
            sigmoid_f := 3;
        ELSIF x =- 13361 THEN
            sigmoid_f := 3;
        ELSIF x =- 13360 THEN
            sigmoid_f := 3;
        ELSIF x =- 13359 THEN
            sigmoid_f := 3;
        ELSIF x =- 13358 THEN
            sigmoid_f := 3;
        ELSIF x =- 13357 THEN
            sigmoid_f := 3;
        ELSIF x =- 13356 THEN
            sigmoid_f := 3;
        ELSIF x =- 13355 THEN
            sigmoid_f := 3;
        ELSIF x =- 13354 THEN
            sigmoid_f := 3;
        ELSIF x =- 13353 THEN
            sigmoid_f := 3;
        ELSIF x =- 13352 THEN
            sigmoid_f := 3;
        ELSIF x =- 13351 THEN
            sigmoid_f := 3;
        ELSIF x =- 13350 THEN
            sigmoid_f := 3;
        ELSIF x =- 13349 THEN
            sigmoid_f := 3;
        ELSIF x =- 13348 THEN
            sigmoid_f := 3;
        ELSIF x =- 13347 THEN
            sigmoid_f := 3;
        ELSIF x =- 13346 THEN
            sigmoid_f := 3;
        ELSIF x =- 13345 THEN
            sigmoid_f := 3;
        ELSIF x =- 13344 THEN
            sigmoid_f := 3;
        ELSIF x =- 13343 THEN
            sigmoid_f := 3;
        ELSIF x =- 13342 THEN
            sigmoid_f := 3;
        ELSIF x =- 13341 THEN
            sigmoid_f := 3;
        ELSIF x =- 13340 THEN
            sigmoid_f := 3;
        ELSIF x =- 13339 THEN
            sigmoid_f := 3;
        ELSIF x =- 13338 THEN
            sigmoid_f := 3;
        ELSIF x =- 13337 THEN
            sigmoid_f := 3;
        ELSIF x =- 13336 THEN
            sigmoid_f := 3;
        ELSIF x =- 13335 THEN
            sigmoid_f := 3;
        ELSIF x =- 13334 THEN
            sigmoid_f := 3;
        ELSIF x =- 13333 THEN
            sigmoid_f := 3;
        ELSIF x =- 13332 THEN
            sigmoid_f := 3;
        ELSIF x =- 13331 THEN
            sigmoid_f := 3;
        ELSIF x =- 13330 THEN
            sigmoid_f := 3;
        ELSIF x =- 13329 THEN
            sigmoid_f := 3;
        ELSIF x =- 13328 THEN
            sigmoid_f := 3;
        ELSIF x =- 13327 THEN
            sigmoid_f := 3;
        ELSIF x =- 13326 THEN
            sigmoid_f := 3;
        ELSIF x =- 13325 THEN
            sigmoid_f := 3;
        ELSIF x =- 13324 THEN
            sigmoid_f := 3;
        ELSIF x =- 13323 THEN
            sigmoid_f := 3;
        ELSIF x =- 13322 THEN
            sigmoid_f := 3;
        ELSIF x =- 13321 THEN
            sigmoid_f := 3;
        ELSIF x =- 13320 THEN
            sigmoid_f := 3;
        ELSIF x =- 13319 THEN
            sigmoid_f := 3;
        ELSIF x =- 13318 THEN
            sigmoid_f := 3;
        ELSIF x =- 13317 THEN
            sigmoid_f := 3;
        ELSIF x =- 13316 THEN
            sigmoid_f := 3;
        ELSIF x =- 13315 THEN
            sigmoid_f := 3;
        ELSIF x =- 13314 THEN
            sigmoid_f := 3;
        ELSIF x =- 13313 THEN
            sigmoid_f := 3;
        ELSIF x =- 13312 THEN
            sigmoid_f := 3;
        ELSIF x =- 13311 THEN
            sigmoid_f := 3;
        ELSIF x =- 13310 THEN
            sigmoid_f := 3;
        ELSIF x =- 13309 THEN
            sigmoid_f := 3;
        ELSIF x =- 13308 THEN
            sigmoid_f := 3;
        ELSIF x =- 13307 THEN
            sigmoid_f := 3;
        ELSIF x =- 13306 THEN
            sigmoid_f := 3;
        ELSIF x =- 13305 THEN
            sigmoid_f := 3;
        ELSIF x =- 13304 THEN
            sigmoid_f := 3;
        ELSIF x =- 13303 THEN
            sigmoid_f := 3;
        ELSIF x =- 13302 THEN
            sigmoid_f := 3;
        ELSIF x =- 13301 THEN
            sigmoid_f := 3;
        ELSIF x =- 13300 THEN
            sigmoid_f := 3;
        ELSIF x =- 13299 THEN
            sigmoid_f := 3;
        ELSIF x =- 13298 THEN
            sigmoid_f := 3;
        ELSIF x =- 13297 THEN
            sigmoid_f := 3;
        ELSIF x =- 13296 THEN
            sigmoid_f := 3;
        ELSIF x =- 13295 THEN
            sigmoid_f := 3;
        ELSIF x =- 13294 THEN
            sigmoid_f := 3;
        ELSIF x =- 13293 THEN
            sigmoid_f := 3;
        ELSIF x =- 13292 THEN
            sigmoid_f := 3;
        ELSIF x =- 13291 THEN
            sigmoid_f := 3;
        ELSIF x =- 13290 THEN
            sigmoid_f := 3;
        ELSIF x =- 13289 THEN
            sigmoid_f := 3;
        ELSIF x =- 13288 THEN
            sigmoid_f := 3;
        ELSIF x =- 13287 THEN
            sigmoid_f := 3;
        ELSIF x =- 13286 THEN
            sigmoid_f := 3;
        ELSIF x =- 13285 THEN
            sigmoid_f := 3;
        ELSIF x =- 13284 THEN
            sigmoid_f := 3;
        ELSIF x =- 13283 THEN
            sigmoid_f := 3;
        ELSIF x =- 13282 THEN
            sigmoid_f := 3;
        ELSIF x =- 13281 THEN
            sigmoid_f := 3;
        ELSIF x =- 13280 THEN
            sigmoid_f := 3;
        ELSIF x =- 13279 THEN
            sigmoid_f := 3;
        ELSIF x =- 13278 THEN
            sigmoid_f := 3;
        ELSIF x =- 13277 THEN
            sigmoid_f := 3;
        ELSIF x =- 13276 THEN
            sigmoid_f := 3;
        ELSIF x =- 13275 THEN
            sigmoid_f := 3;
        ELSIF x =- 13274 THEN
            sigmoid_f := 3;
        ELSIF x =- 13273 THEN
            sigmoid_f := 3;
        ELSIF x =- 13272 THEN
            sigmoid_f := 3;
        ELSIF x =- 13271 THEN
            sigmoid_f := 3;
        ELSIF x =- 13270 THEN
            sigmoid_f := 3;
        ELSIF x =- 13269 THEN
            sigmoid_f := 3;
        ELSIF x =- 13268 THEN
            sigmoid_f := 3;
        ELSIF x =- 13267 THEN
            sigmoid_f := 3;
        ELSIF x =- 13266 THEN
            sigmoid_f := 3;
        ELSIF x =- 13265 THEN
            sigmoid_f := 3;
        ELSIF x =- 13264 THEN
            sigmoid_f := 3;
        ELSIF x =- 13263 THEN
            sigmoid_f := 3;
        ELSIF x =- 13262 THEN
            sigmoid_f := 3;
        ELSIF x =- 13261 THEN
            sigmoid_f := 3;
        ELSIF x =- 13260 THEN
            sigmoid_f := 3;
        ELSIF x =- 13259 THEN
            sigmoid_f := 3;
        ELSIF x =- 13258 THEN
            sigmoid_f := 3;
        ELSIF x =- 13257 THEN
            sigmoid_f := 3;
        ELSIF x =- 13256 THEN
            sigmoid_f := 3;
        ELSIF x =- 13255 THEN
            sigmoid_f := 3;
        ELSIF x =- 13254 THEN
            sigmoid_f := 3;
        ELSIF x =- 13253 THEN
            sigmoid_f := 3;
        ELSIF x =- 13252 THEN
            sigmoid_f := 3;
        ELSIF x =- 13251 THEN
            sigmoid_f := 3;
        ELSIF x =- 13250 THEN
            sigmoid_f := 3;
        ELSIF x =- 13249 THEN
            sigmoid_f := 3;
        ELSIF x =- 13248 THEN
            sigmoid_f := 3;
        ELSIF x =- 13247 THEN
            sigmoid_f := 3;
        ELSIF x =- 13246 THEN
            sigmoid_f := 3;
        ELSIF x =- 13245 THEN
            sigmoid_f := 3;
        ELSIF x =- 13244 THEN
            sigmoid_f := 3;
        ELSIF x =- 13243 THEN
            sigmoid_f := 3;
        ELSIF x =- 13242 THEN
            sigmoid_f := 3;
        ELSIF x =- 13241 THEN
            sigmoid_f := 3;
        ELSIF x =- 13240 THEN
            sigmoid_f := 3;
        ELSIF x =- 13239 THEN
            sigmoid_f := 3;
        ELSIF x =- 13238 THEN
            sigmoid_f := 3;
        ELSIF x =- 13237 THEN
            sigmoid_f := 3;
        ELSIF x =- 13236 THEN
            sigmoid_f := 3;
        ELSIF x =- 13235 THEN
            sigmoid_f := 3;
        ELSIF x =- 13234 THEN
            sigmoid_f := 3;
        ELSIF x =- 13233 THEN
            sigmoid_f := 3;
        ELSIF x =- 13232 THEN
            sigmoid_f := 3;
        ELSIF x =- 13231 THEN
            sigmoid_f := 3;
        ELSIF x =- 13230 THEN
            sigmoid_f := 3;
        ELSIF x =- 13229 THEN
            sigmoid_f := 3;
        ELSIF x =- 13228 THEN
            sigmoid_f := 3;
        ELSIF x =- 13227 THEN
            sigmoid_f := 3;
        ELSIF x =- 13226 THEN
            sigmoid_f := 3;
        ELSIF x =- 13225 THEN
            sigmoid_f := 3;
        ELSIF x =- 13224 THEN
            sigmoid_f := 3;
        ELSIF x =- 13223 THEN
            sigmoid_f := 3;
        ELSIF x =- 13222 THEN
            sigmoid_f := 3;
        ELSIF x =- 13221 THEN
            sigmoid_f := 3;
        ELSIF x =- 13220 THEN
            sigmoid_f := 3;
        ELSIF x =- 13219 THEN
            sigmoid_f := 3;
        ELSIF x =- 13218 THEN
            sigmoid_f := 3;
        ELSIF x =- 13217 THEN
            sigmoid_f := 3;
        ELSIF x =- 13216 THEN
            sigmoid_f := 3;
        ELSIF x =- 13215 THEN
            sigmoid_f := 3;
        ELSIF x =- 13214 THEN
            sigmoid_f := 3;
        ELSIF x =- 13213 THEN
            sigmoid_f := 3;
        ELSIF x =- 13212 THEN
            sigmoid_f := 3;
        ELSIF x =- 13211 THEN
            sigmoid_f := 3;
        ELSIF x =- 13210 THEN
            sigmoid_f := 3;
        ELSIF x =- 13209 THEN
            sigmoid_f := 3;
        ELSIF x =- 13208 THEN
            sigmoid_f := 3;
        ELSIF x =- 13207 THEN
            sigmoid_f := 3;
        ELSIF x =- 13206 THEN
            sigmoid_f := 3;
        ELSIF x =- 13205 THEN
            sigmoid_f := 3;
        ELSIF x =- 13204 THEN
            sigmoid_f := 3;
        ELSIF x =- 13203 THEN
            sigmoid_f := 3;
        ELSIF x =- 13202 THEN
            sigmoid_f := 3;
        ELSIF x =- 13201 THEN
            sigmoid_f := 3;
        ELSIF x =- 13200 THEN
            sigmoid_f := 3;
        ELSIF x =- 13199 THEN
            sigmoid_f := 3;
        ELSIF x =- 13198 THEN
            sigmoid_f := 3;
        ELSIF x =- 13197 THEN
            sigmoid_f := 3;
        ELSIF x =- 13196 THEN
            sigmoid_f := 3;
        ELSIF x =- 13195 THEN
            sigmoid_f := 3;
        ELSIF x =- 13194 THEN
            sigmoid_f := 3;
        ELSIF x =- 13193 THEN
            sigmoid_f := 3;
        ELSIF x =- 13192 THEN
            sigmoid_f := 3;
        ELSIF x =- 13191 THEN
            sigmoid_f := 3;
        ELSIF x =- 13190 THEN
            sigmoid_f := 3;
        ELSIF x =- 13189 THEN
            sigmoid_f := 3;
        ELSIF x =- 13188 THEN
            sigmoid_f := 3;
        ELSIF x =- 13187 THEN
            sigmoid_f := 3;
        ELSIF x =- 13186 THEN
            sigmoid_f := 3;
        ELSIF x =- 13185 THEN
            sigmoid_f := 3;
        ELSIF x =- 13184 THEN
            sigmoid_f := 3;
        ELSIF x =- 13183 THEN
            sigmoid_f := 3;
        ELSIF x =- 13182 THEN
            sigmoid_f := 3;
        ELSIF x =- 13181 THEN
            sigmoid_f := 3;
        ELSIF x =- 13180 THEN
            sigmoid_f := 3;
        ELSIF x =- 13179 THEN
            sigmoid_f := 3;
        ELSIF x =- 13178 THEN
            sigmoid_f := 3;
        ELSIF x =- 13177 THEN
            sigmoid_f := 3;
        ELSIF x =- 13176 THEN
            sigmoid_f := 3;
        ELSIF x =- 13175 THEN
            sigmoid_f := 3;
        ELSIF x =- 13174 THEN
            sigmoid_f := 3;
        ELSIF x =- 13173 THEN
            sigmoid_f := 3;
        ELSIF x =- 13172 THEN
            sigmoid_f := 3;
        ELSIF x =- 13171 THEN
            sigmoid_f := 3;
        ELSIF x =- 13170 THEN
            sigmoid_f := 3;
        ELSIF x =- 13169 THEN
            sigmoid_f := 3;
        ELSIF x =- 13168 THEN
            sigmoid_f := 3;
        ELSIF x =- 13167 THEN
            sigmoid_f := 3;
        ELSIF x =- 13166 THEN
            sigmoid_f := 3;
        ELSIF x =- 13165 THEN
            sigmoid_f := 3;
        ELSIF x =- 13164 THEN
            sigmoid_f := 3;
        ELSIF x =- 13163 THEN
            sigmoid_f := 3;
        ELSIF x =- 13162 THEN
            sigmoid_f := 3;
        ELSIF x =- 13161 THEN
            sigmoid_f := 3;
        ELSIF x =- 13160 THEN
            sigmoid_f := 3;
        ELSIF x =- 13159 THEN
            sigmoid_f := 3;
        ELSIF x =- 13158 THEN
            sigmoid_f := 3;
        ELSIF x =- 13157 THEN
            sigmoid_f := 3;
        ELSIF x =- 13156 THEN
            sigmoid_f := 3;
        ELSIF x =- 13155 THEN
            sigmoid_f := 3;
        ELSIF x =- 13154 THEN
            sigmoid_f := 3;
        ELSIF x =- 13153 THEN
            sigmoid_f := 3;
        ELSIF x =- 13152 THEN
            sigmoid_f := 3;
        ELSIF x =- 13151 THEN
            sigmoid_f := 3;
        ELSIF x =- 13150 THEN
            sigmoid_f := 3;
        ELSIF x =- 13149 THEN
            sigmoid_f := 3;
        ELSIF x =- 13148 THEN
            sigmoid_f := 3;
        ELSIF x =- 13147 THEN
            sigmoid_f := 3;
        ELSIF x =- 13146 THEN
            sigmoid_f := 3;
        ELSIF x =- 13145 THEN
            sigmoid_f := 3;
        ELSIF x =- 13144 THEN
            sigmoid_f := 3;
        ELSIF x =- 13143 THEN
            sigmoid_f := 3;
        ELSIF x =- 13142 THEN
            sigmoid_f := 3;
        ELSIF x =- 13141 THEN
            sigmoid_f := 3;
        ELSIF x =- 13140 THEN
            sigmoid_f := 3;
        ELSIF x =- 13139 THEN
            sigmoid_f := 3;
        ELSIF x =- 13138 THEN
            sigmoid_f := 3;
        ELSIF x =- 13137 THEN
            sigmoid_f := 3;
        ELSIF x =- 13136 THEN
            sigmoid_f := 3;
        ELSIF x =- 13135 THEN
            sigmoid_f := 3;
        ELSIF x =- 13134 THEN
            sigmoid_f := 3;
        ELSIF x =- 13133 THEN
            sigmoid_f := 3;
        ELSIF x =- 13132 THEN
            sigmoid_f := 3;
        ELSIF x =- 13131 THEN
            sigmoid_f := 3;
        ELSIF x =- 13130 THEN
            sigmoid_f := 3;
        ELSIF x =- 13129 THEN
            sigmoid_f := 3;
        ELSIF x =- 13128 THEN
            sigmoid_f := 3;
        ELSIF x =- 13127 THEN
            sigmoid_f := 3;
        ELSIF x =- 13126 THEN
            sigmoid_f := 3;
        ELSIF x =- 13125 THEN
            sigmoid_f := 3;
        ELSIF x =- 13124 THEN
            sigmoid_f := 3;
        ELSIF x =- 13123 THEN
            sigmoid_f := 3;
        ELSIF x =- 13122 THEN
            sigmoid_f := 3;
        ELSIF x =- 13121 THEN
            sigmoid_f := 3;
        ELSIF x =- 13120 THEN
            sigmoid_f := 3;
        ELSIF x =- 13119 THEN
            sigmoid_f := 3;
        ELSIF x =- 13118 THEN
            sigmoid_f := 3;
        ELSIF x =- 13117 THEN
            sigmoid_f := 3;
        ELSIF x =- 13116 THEN
            sigmoid_f := 3;
        ELSIF x =- 13115 THEN
            sigmoid_f := 3;
        ELSIF x =- 13114 THEN
            sigmoid_f := 3;
        ELSIF x =- 13113 THEN
            sigmoid_f := 3;
        ELSIF x =- 13112 THEN
            sigmoid_f := 3;
        ELSIF x =- 13111 THEN
            sigmoid_f := 3;
        ELSIF x =- 13110 THEN
            sigmoid_f := 3;
        ELSIF x =- 13109 THEN
            sigmoid_f := 3;
        ELSIF x =- 13108 THEN
            sigmoid_f := 3;
        ELSIF x =- 13107 THEN
            sigmoid_f := 3;
        ELSIF x =- 13106 THEN
            sigmoid_f := 3;
        ELSIF x =- 13105 THEN
            sigmoid_f := 3;
        ELSIF x =- 13104 THEN
            sigmoid_f := 3;
        ELSIF x =- 13103 THEN
            sigmoid_f := 3;
        ELSIF x =- 13102 THEN
            sigmoid_f := 3;
        ELSIF x =- 13101 THEN
            sigmoid_f := 3;
        ELSIF x =- 13100 THEN
            sigmoid_f := 3;
        ELSIF x =- 13099 THEN
            sigmoid_f := 3;
        ELSIF x =- 13098 THEN
            sigmoid_f := 3;
        ELSIF x =- 13097 THEN
            sigmoid_f := 3;
        ELSIF x =- 13096 THEN
            sigmoid_f := 3;
        ELSIF x =- 13095 THEN
            sigmoid_f := 3;
        ELSIF x =- 13094 THEN
            sigmoid_f := 3;
        ELSIF x =- 13093 THEN
            sigmoid_f := 3;
        ELSIF x =- 13092 THEN
            sigmoid_f := 3;
        ELSIF x =- 13091 THEN
            sigmoid_f := 3;
        ELSIF x =- 13090 THEN
            sigmoid_f := 3;
        ELSIF x =- 13089 THEN
            sigmoid_f := 3;
        ELSIF x =- 13088 THEN
            sigmoid_f := 3;
        ELSIF x =- 13087 THEN
            sigmoid_f := 3;
        ELSIF x =- 13086 THEN
            sigmoid_f := 3;
        ELSIF x =- 13085 THEN
            sigmoid_f := 3;
        ELSIF x =- 13084 THEN
            sigmoid_f := 3;
        ELSIF x =- 13083 THEN
            sigmoid_f := 3;
        ELSIF x =- 13082 THEN
            sigmoid_f := 3;
        ELSIF x =- 13081 THEN
            sigmoid_f := 3;
        ELSIF x =- 13080 THEN
            sigmoid_f := 3;
        ELSIF x =- 13079 THEN
            sigmoid_f := 3;
        ELSIF x =- 13078 THEN
            sigmoid_f := 3;
        ELSIF x =- 13077 THEN
            sigmoid_f := 3;
        ELSIF x =- 13076 THEN
            sigmoid_f := 3;
        ELSIF x =- 13075 THEN
            sigmoid_f := 3;
        ELSIF x =- 13074 THEN
            sigmoid_f := 3;
        ELSIF x =- 13073 THEN
            sigmoid_f := 3;
        ELSIF x =- 13072 THEN
            sigmoid_f := 3;
        ELSIF x =- 13071 THEN
            sigmoid_f := 3;
        ELSIF x =- 13070 THEN
            sigmoid_f := 3;
        ELSIF x =- 13069 THEN
            sigmoid_f := 3;
        ELSIF x =- 13068 THEN
            sigmoid_f := 3;
        ELSIF x =- 13067 THEN
            sigmoid_f := 3;
        ELSIF x =- 13066 THEN
            sigmoid_f := 3;
        ELSIF x =- 13065 THEN
            sigmoid_f := 3;
        ELSIF x =- 13064 THEN
            sigmoid_f := 3;
        ELSIF x =- 13063 THEN
            sigmoid_f := 3;
        ELSIF x =- 13062 THEN
            sigmoid_f := 3;
        ELSIF x =- 13061 THEN
            sigmoid_f := 3;
        ELSIF x =- 13060 THEN
            sigmoid_f := 3;
        ELSIF x =- 13059 THEN
            sigmoid_f := 3;
        ELSIF x =- 13058 THEN
            sigmoid_f := 3;
        ELSIF x =- 13057 THEN
            sigmoid_f := 3;
        ELSIF x =- 13056 THEN
            sigmoid_f := 3;
        ELSIF x =- 13055 THEN
            sigmoid_f := 3;
        ELSIF x =- 13054 THEN
            sigmoid_f := 3;
        ELSIF x =- 13053 THEN
            sigmoid_f := 3;
        ELSIF x =- 13052 THEN
            sigmoid_f := 3;
        ELSIF x =- 13051 THEN
            sigmoid_f := 3;
        ELSIF x =- 13050 THEN
            sigmoid_f := 3;
        ELSIF x =- 13049 THEN
            sigmoid_f := 3;
        ELSIF x =- 13048 THEN
            sigmoid_f := 3;
        ELSIF x =- 13047 THEN
            sigmoid_f := 3;
        ELSIF x =- 13046 THEN
            sigmoid_f := 3;
        ELSIF x =- 13045 THEN
            sigmoid_f := 3;
        ELSIF x =- 13044 THEN
            sigmoid_f := 3;
        ELSIF x =- 13043 THEN
            sigmoid_f := 3;
        ELSIF x =- 13042 THEN
            sigmoid_f := 3;
        ELSIF x =- 13041 THEN
            sigmoid_f := 3;
        ELSIF x =- 13040 THEN
            sigmoid_f := 3;
        ELSIF x =- 13039 THEN
            sigmoid_f := 3;
        ELSIF x =- 13038 THEN
            sigmoid_f := 3;
        ELSIF x =- 13037 THEN
            sigmoid_f := 3;
        ELSIF x =- 13036 THEN
            sigmoid_f := 3;
        ELSIF x =- 13035 THEN
            sigmoid_f := 3;
        ELSIF x =- 13034 THEN
            sigmoid_f := 3;
        ELSIF x =- 13033 THEN
            sigmoid_f := 3;
        ELSIF x =- 13032 THEN
            sigmoid_f := 3;
        ELSIF x =- 13031 THEN
            sigmoid_f := 3;
        ELSIF x =- 13030 THEN
            sigmoid_f := 3;
        ELSIF x =- 13029 THEN
            sigmoid_f := 3;
        ELSIF x =- 13028 THEN
            sigmoid_f := 3;
        ELSIF x =- 13027 THEN
            sigmoid_f := 3;
        ELSIF x =- 13026 THEN
            sigmoid_f := 3;
        ELSIF x =- 13025 THEN
            sigmoid_f := 3;
        ELSIF x =- 13024 THEN
            sigmoid_f := 3;
        ELSIF x =- 13023 THEN
            sigmoid_f := 3;
        ELSIF x =- 13022 THEN
            sigmoid_f := 3;
        ELSIF x =- 13021 THEN
            sigmoid_f := 3;
        ELSIF x =- 13020 THEN
            sigmoid_f := 3;
        ELSIF x =- 13019 THEN
            sigmoid_f := 3;
        ELSIF x =- 13018 THEN
            sigmoid_f := 3;
        ELSIF x =- 13017 THEN
            sigmoid_f := 3;
        ELSIF x =- 13016 THEN
            sigmoid_f := 3;
        ELSIF x =- 13015 THEN
            sigmoid_f := 3;
        ELSIF x =- 13014 THEN
            sigmoid_f := 3;
        ELSIF x =- 13013 THEN
            sigmoid_f := 3;
        ELSIF x =- 13012 THEN
            sigmoid_f := 3;
        ELSIF x =- 13011 THEN
            sigmoid_f := 3;
        ELSIF x =- 13010 THEN
            sigmoid_f := 3;
        ELSIF x =- 13009 THEN
            sigmoid_f := 3;
        ELSIF x =- 13008 THEN
            sigmoid_f := 3;
        ELSIF x =- 13007 THEN
            sigmoid_f := 3;
        ELSIF x =- 13006 THEN
            sigmoid_f := 3;
        ELSIF x =- 13005 THEN
            sigmoid_f := 3;
        ELSIF x =- 13004 THEN
            sigmoid_f := 3;
        ELSIF x =- 13003 THEN
            sigmoid_f := 3;
        ELSIF x =- 13002 THEN
            sigmoid_f := 3;
        ELSIF x =- 13001 THEN
            sigmoid_f := 3;
        ELSIF x =- 13000 THEN
            sigmoid_f := 3;
        ELSIF x =- 12999 THEN
            sigmoid_f := 3;
        ELSIF x =- 12998 THEN
            sigmoid_f := 3;
        ELSIF x =- 12997 THEN
            sigmoid_f := 3;
        ELSIF x =- 12996 THEN
            sigmoid_f := 3;
        ELSIF x =- 12995 THEN
            sigmoid_f := 3;
        ELSIF x =- 12994 THEN
            sigmoid_f := 3;
        ELSIF x =- 12993 THEN
            sigmoid_f := 3;
        ELSIF x =- 12992 THEN
            sigmoid_f := 3;
        ELSIF x =- 12991 THEN
            sigmoid_f := 3;
        ELSIF x =- 12990 THEN
            sigmoid_f := 3;
        ELSIF x =- 12989 THEN
            sigmoid_f := 3;
        ELSIF x =- 12988 THEN
            sigmoid_f := 3;
        ELSIF x =- 12987 THEN
            sigmoid_f := 3;
        ELSIF x =- 12986 THEN
            sigmoid_f := 3;
        ELSIF x =- 12985 THEN
            sigmoid_f := 3;
        ELSIF x =- 12984 THEN
            sigmoid_f := 3;
        ELSIF x =- 12983 THEN
            sigmoid_f := 3;
        ELSIF x =- 12982 THEN
            sigmoid_f := 3;
        ELSIF x =- 12981 THEN
            sigmoid_f := 3;
        ELSIF x =- 12980 THEN
            sigmoid_f := 3;
        ELSIF x =- 12979 THEN
            sigmoid_f := 3;
        ELSIF x =- 12978 THEN
            sigmoid_f := 3;
        ELSIF x =- 12977 THEN
            sigmoid_f := 3;
        ELSIF x =- 12976 THEN
            sigmoid_f := 3;
        ELSIF x =- 12975 THEN
            sigmoid_f := 3;
        ELSIF x =- 12974 THEN
            sigmoid_f := 3;
        ELSIF x =- 12973 THEN
            sigmoid_f := 3;
        ELSIF x =- 12972 THEN
            sigmoid_f := 3;
        ELSIF x =- 12971 THEN
            sigmoid_f := 3;
        ELSIF x =- 12970 THEN
            sigmoid_f := 3;
        ELSIF x =- 12969 THEN
            sigmoid_f := 3;
        ELSIF x =- 12968 THEN
            sigmoid_f := 3;
        ELSIF x =- 12967 THEN
            sigmoid_f := 3;
        ELSIF x =- 12966 THEN
            sigmoid_f := 3;
        ELSIF x =- 12965 THEN
            sigmoid_f := 3;
        ELSIF x =- 12964 THEN
            sigmoid_f := 3;
        ELSIF x =- 12963 THEN
            sigmoid_f := 3;
        ELSIF x =- 12962 THEN
            sigmoid_f := 3;
        ELSIF x =- 12961 THEN
            sigmoid_f := 3;
        ELSIF x =- 12960 THEN
            sigmoid_f := 3;
        ELSIF x =- 12959 THEN
            sigmoid_f := 3;
        ELSIF x =- 12958 THEN
            sigmoid_f := 3;
        ELSIF x =- 12957 THEN
            sigmoid_f := 3;
        ELSIF x =- 12956 THEN
            sigmoid_f := 3;
        ELSIF x =- 12955 THEN
            sigmoid_f := 3;
        ELSIF x =- 12954 THEN
            sigmoid_f := 3;
        ELSIF x =- 12953 THEN
            sigmoid_f := 3;
        ELSIF x =- 12952 THEN
            sigmoid_f := 3;
        ELSIF x =- 12951 THEN
            sigmoid_f := 3;
        ELSIF x =- 12950 THEN
            sigmoid_f := 3;
        ELSIF x =- 12949 THEN
            sigmoid_f := 3;
        ELSIF x =- 12948 THEN
            sigmoid_f := 3;
        ELSIF x =- 12947 THEN
            sigmoid_f := 3;
        ELSIF x =- 12946 THEN
            sigmoid_f := 3;
        ELSIF x =- 12945 THEN
            sigmoid_f := 3;
        ELSIF x =- 12944 THEN
            sigmoid_f := 3;
        ELSIF x =- 12943 THEN
            sigmoid_f := 3;
        ELSIF x =- 12942 THEN
            sigmoid_f := 3;
        ELSIF x =- 12941 THEN
            sigmoid_f := 3;
        ELSIF x =- 12940 THEN
            sigmoid_f := 3;
        ELSIF x =- 12939 THEN
            sigmoid_f := 3;
        ELSIF x =- 12938 THEN
            sigmoid_f := 3;
        ELSIF x =- 12937 THEN
            sigmoid_f := 3;
        ELSIF x =- 12936 THEN
            sigmoid_f := 3;
        ELSIF x =- 12935 THEN
            sigmoid_f := 3;
        ELSIF x =- 12934 THEN
            sigmoid_f := 3;
        ELSIF x =- 12933 THEN
            sigmoid_f := 3;
        ELSIF x =- 12932 THEN
            sigmoid_f := 3;
        ELSIF x =- 12931 THEN
            sigmoid_f := 3;
        ELSIF x =- 12930 THEN
            sigmoid_f := 3;
        ELSIF x =- 12929 THEN
            sigmoid_f := 3;
        ELSIF x =- 12928 THEN
            sigmoid_f := 3;
        ELSIF x =- 12927 THEN
            sigmoid_f := 3;
        ELSIF x =- 12926 THEN
            sigmoid_f := 3;
        ELSIF x =- 12925 THEN
            sigmoid_f := 3;
        ELSIF x =- 12924 THEN
            sigmoid_f := 3;
        ELSIF x =- 12923 THEN
            sigmoid_f := 3;
        ELSIF x =- 12922 THEN
            sigmoid_f := 3;
        ELSIF x =- 12921 THEN
            sigmoid_f := 3;
        ELSIF x =- 12920 THEN
            sigmoid_f := 3;
        ELSIF x =- 12919 THEN
            sigmoid_f := 3;
        ELSIF x =- 12918 THEN
            sigmoid_f := 3;
        ELSIF x =- 12917 THEN
            sigmoid_f := 3;
        ELSIF x =- 12916 THEN
            sigmoid_f := 3;
        ELSIF x =- 12915 THEN
            sigmoid_f := 3;
        ELSIF x =- 12914 THEN
            sigmoid_f := 3;
        ELSIF x =- 12913 THEN
            sigmoid_f := 3;
        ELSIF x =- 12912 THEN
            sigmoid_f := 3;
        ELSIF x =- 12911 THEN
            sigmoid_f := 3;
        ELSIF x =- 12910 THEN
            sigmoid_f := 3;
        ELSIF x =- 12909 THEN
            sigmoid_f := 3;
        ELSIF x =- 12908 THEN
            sigmoid_f := 3;
        ELSIF x =- 12907 THEN
            sigmoid_f := 3;
        ELSIF x =- 12906 THEN
            sigmoid_f := 3;
        ELSIF x =- 12905 THEN
            sigmoid_f := 3;
        ELSIF x =- 12904 THEN
            sigmoid_f := 3;
        ELSIF x =- 12903 THEN
            sigmoid_f := 3;
        ELSIF x =- 12902 THEN
            sigmoid_f := 3;
        ELSIF x =- 12901 THEN
            sigmoid_f := 3;
        ELSIF x =- 12900 THEN
            sigmoid_f := 3;
        ELSIF x =- 12899 THEN
            sigmoid_f := 3;
        ELSIF x =- 12898 THEN
            sigmoid_f := 3;
        ELSIF x =- 12897 THEN
            sigmoid_f := 3;
        ELSIF x =- 12896 THEN
            sigmoid_f := 3;
        ELSIF x =- 12895 THEN
            sigmoid_f := 3;
        ELSIF x =- 12894 THEN
            sigmoid_f := 3;
        ELSIF x =- 12893 THEN
            sigmoid_f := 3;
        ELSIF x =- 12892 THEN
            sigmoid_f := 3;
        ELSIF x =- 12891 THEN
            sigmoid_f := 3;
        ELSIF x =- 12890 THEN
            sigmoid_f := 3;
        ELSIF x =- 12889 THEN
            sigmoid_f := 3;
        ELSIF x =- 12888 THEN
            sigmoid_f := 3;
        ELSIF x =- 12887 THEN
            sigmoid_f := 3;
        ELSIF x =- 12886 THEN
            sigmoid_f := 3;
        ELSIF x =- 12885 THEN
            sigmoid_f := 3;
        ELSIF x =- 12884 THEN
            sigmoid_f := 3;
        ELSIF x =- 12883 THEN
            sigmoid_f := 3;
        ELSIF x =- 12882 THEN
            sigmoid_f := 3;
        ELSIF x =- 12881 THEN
            sigmoid_f := 3;
        ELSIF x =- 12880 THEN
            sigmoid_f := 3;
        ELSIF x =- 12879 THEN
            sigmoid_f := 3;
        ELSIF x =- 12878 THEN
            sigmoid_f := 3;
        ELSIF x =- 12877 THEN
            sigmoid_f := 3;
        ELSIF x =- 12876 THEN
            sigmoid_f := 3;
        ELSIF x =- 12875 THEN
            sigmoid_f := 3;
        ELSIF x =- 12874 THEN
            sigmoid_f := 3;
        ELSIF x =- 12873 THEN
            sigmoid_f := 3;
        ELSIF x =- 12872 THEN
            sigmoid_f := 3;
        ELSIF x =- 12871 THEN
            sigmoid_f := 3;
        ELSIF x =- 12870 THEN
            sigmoid_f := 3;
        ELSIF x =- 12869 THEN
            sigmoid_f := 3;
        ELSIF x =- 12868 THEN
            sigmoid_f := 3;
        ELSIF x =- 12867 THEN
            sigmoid_f := 3;
        ELSIF x =- 12866 THEN
            sigmoid_f := 3;
        ELSIF x =- 12865 THEN
            sigmoid_f := 3;
        ELSIF x =- 12864 THEN
            sigmoid_f := 3;
        ELSIF x =- 12863 THEN
            sigmoid_f := 3;
        ELSIF x =- 12862 THEN
            sigmoid_f := 3;
        ELSIF x =- 12861 THEN
            sigmoid_f := 3;
        ELSIF x =- 12860 THEN
            sigmoid_f := 3;
        ELSIF x =- 12859 THEN
            sigmoid_f := 3;
        ELSIF x =- 12858 THEN
            sigmoid_f := 3;
        ELSIF x =- 12857 THEN
            sigmoid_f := 3;
        ELSIF x =- 12856 THEN
            sigmoid_f := 3;
        ELSIF x =- 12855 THEN
            sigmoid_f := 3;
        ELSIF x =- 12854 THEN
            sigmoid_f := 3;
        ELSIF x =- 12853 THEN
            sigmoid_f := 3;
        ELSIF x =- 12852 THEN
            sigmoid_f := 3;
        ELSIF x =- 12851 THEN
            sigmoid_f := 3;
        ELSIF x =- 12850 THEN
            sigmoid_f := 3;
        ELSIF x =- 12849 THEN
            sigmoid_f := 3;
        ELSIF x =- 12848 THEN
            sigmoid_f := 3;
        ELSIF x =- 12847 THEN
            sigmoid_f := 3;
        ELSIF x =- 12846 THEN
            sigmoid_f := 3;
        ELSIF x =- 12845 THEN
            sigmoid_f := 3;
        ELSIF x =- 12844 THEN
            sigmoid_f := 3;
        ELSIF x =- 12843 THEN
            sigmoid_f := 3;
        ELSIF x =- 12842 THEN
            sigmoid_f := 3;
        ELSIF x =- 12841 THEN
            sigmoid_f := 3;
        ELSIF x =- 12840 THEN
            sigmoid_f := 3;
        ELSIF x =- 12839 THEN
            sigmoid_f := 3;
        ELSIF x =- 12838 THEN
            sigmoid_f := 3;
        ELSIF x =- 12837 THEN
            sigmoid_f := 3;
        ELSIF x =- 12836 THEN
            sigmoid_f := 3;
        ELSIF x =- 12835 THEN
            sigmoid_f := 3;
        ELSIF x =- 12834 THEN
            sigmoid_f := 3;
        ELSIF x =- 12833 THEN
            sigmoid_f := 3;
        ELSIF x =- 12832 THEN
            sigmoid_f := 3;
        ELSIF x =- 12831 THEN
            sigmoid_f := 3;
        ELSIF x =- 12830 THEN
            sigmoid_f := 3;
        ELSIF x =- 12829 THEN
            sigmoid_f := 3;
        ELSIF x =- 12828 THEN
            sigmoid_f := 3;
        ELSIF x =- 12827 THEN
            sigmoid_f := 3;
        ELSIF x =- 12826 THEN
            sigmoid_f := 3;
        ELSIF x =- 12825 THEN
            sigmoid_f := 3;
        ELSIF x =- 12824 THEN
            sigmoid_f := 3;
        ELSIF x =- 12823 THEN
            sigmoid_f := 3;
        ELSIF x =- 12822 THEN
            sigmoid_f := 3;
        ELSIF x =- 12821 THEN
            sigmoid_f := 3;
        ELSIF x =- 12820 THEN
            sigmoid_f := 3;
        ELSIF x =- 12819 THEN
            sigmoid_f := 3;
        ELSIF x =- 12818 THEN
            sigmoid_f := 3;
        ELSIF x =- 12817 THEN
            sigmoid_f := 3;
        ELSIF x =- 12816 THEN
            sigmoid_f := 3;
        ELSIF x =- 12815 THEN
            sigmoid_f := 3;
        ELSIF x =- 12814 THEN
            sigmoid_f := 3;
        ELSIF x =- 12813 THEN
            sigmoid_f := 3;
        ELSIF x =- 12812 THEN
            sigmoid_f := 3;
        ELSIF x =- 12811 THEN
            sigmoid_f := 3;
        ELSIF x =- 12810 THEN
            sigmoid_f := 3;
        ELSIF x =- 12809 THEN
            sigmoid_f := 3;
        ELSIF x =- 12808 THEN
            sigmoid_f := 3;
        ELSIF x =- 12807 THEN
            sigmoid_f := 3;
        ELSIF x =- 12806 THEN
            sigmoid_f := 3;
        ELSIF x =- 12805 THEN
            sigmoid_f := 3;
        ELSIF x =- 12804 THEN
            sigmoid_f := 3;
        ELSIF x =- 12803 THEN
            sigmoid_f := 3;
        ELSIF x =- 12802 THEN
            sigmoid_f := 3;
        ELSIF x =- 12801 THEN
            sigmoid_f := 3;
        ELSIF x =- 12800 THEN
            sigmoid_f := 3;
        ELSIF x =- 12799 THEN
            sigmoid_f := 4;
        ELSIF x =- 12798 THEN
            sigmoid_f := 4;
        ELSIF x =- 12797 THEN
            sigmoid_f := 4;
        ELSIF x =- 12796 THEN
            sigmoid_f := 4;
        ELSIF x =- 12795 THEN
            sigmoid_f := 4;
        ELSIF x =- 12794 THEN
            sigmoid_f := 4;
        ELSIF x =- 12793 THEN
            sigmoid_f := 4;
        ELSIF x =- 12792 THEN
            sigmoid_f := 4;
        ELSIF x =- 12791 THEN
            sigmoid_f := 4;
        ELSIF x =- 12790 THEN
            sigmoid_f := 4;
        ELSIF x =- 12789 THEN
            sigmoid_f := 4;
        ELSIF x =- 12788 THEN
            sigmoid_f := 4;
        ELSIF x =- 12787 THEN
            sigmoid_f := 4;
        ELSIF x =- 12786 THEN
            sigmoid_f := 4;
        ELSIF x =- 12785 THEN
            sigmoid_f := 4;
        ELSIF x =- 12784 THEN
            sigmoid_f := 4;
        ELSIF x =- 12783 THEN
            sigmoid_f := 4;
        ELSIF x =- 12782 THEN
            sigmoid_f := 4;
        ELSIF x =- 12781 THEN
            sigmoid_f := 4;
        ELSIF x =- 12780 THEN
            sigmoid_f := 4;
        ELSIF x =- 12779 THEN
            sigmoid_f := 4;
        ELSIF x =- 12778 THEN
            sigmoid_f := 4;
        ELSIF x =- 12777 THEN
            sigmoid_f := 4;
        ELSIF x =- 12776 THEN
            sigmoid_f := 4;
        ELSIF x =- 12775 THEN
            sigmoid_f := 4;
        ELSIF x =- 12774 THEN
            sigmoid_f := 4;
        ELSIF x =- 12773 THEN
            sigmoid_f := 4;
        ELSIF x =- 12772 THEN
            sigmoid_f := 4;
        ELSIF x =- 12771 THEN
            sigmoid_f := 4;
        ELSIF x =- 12770 THEN
            sigmoid_f := 4;
        ELSIF x =- 12769 THEN
            sigmoid_f := 4;
        ELSIF x =- 12768 THEN
            sigmoid_f := 4;
        ELSIF x =- 12767 THEN
            sigmoid_f := 4;
        ELSIF x =- 12766 THEN
            sigmoid_f := 4;
        ELSIF x =- 12765 THEN
            sigmoid_f := 4;
        ELSIF x =- 12764 THEN
            sigmoid_f := 4;
        ELSIF x =- 12763 THEN
            sigmoid_f := 4;
        ELSIF x =- 12762 THEN
            sigmoid_f := 4;
        ELSIF x =- 12761 THEN
            sigmoid_f := 4;
        ELSIF x =- 12760 THEN
            sigmoid_f := 4;
        ELSIF x =- 12759 THEN
            sigmoid_f := 4;
        ELSIF x =- 12758 THEN
            sigmoid_f := 4;
        ELSIF x =- 12757 THEN
            sigmoid_f := 4;
        ELSIF x =- 12756 THEN
            sigmoid_f := 4;
        ELSIF x =- 12755 THEN
            sigmoid_f := 4;
        ELSIF x =- 12754 THEN
            sigmoid_f := 4;
        ELSIF x =- 12753 THEN
            sigmoid_f := 4;
        ELSIF x =- 12752 THEN
            sigmoid_f := 4;
        ELSIF x =- 12751 THEN
            sigmoid_f := 4;
        ELSIF x =- 12750 THEN
            sigmoid_f := 4;
        ELSIF x =- 12749 THEN
            sigmoid_f := 4;
        ELSIF x =- 12748 THEN
            sigmoid_f := 4;
        ELSIF x =- 12747 THEN
            sigmoid_f := 4;
        ELSIF x =- 12746 THEN
            sigmoid_f := 4;
        ELSIF x =- 12745 THEN
            sigmoid_f := 4;
        ELSIF x =- 12744 THEN
            sigmoid_f := 4;
        ELSIF x =- 12743 THEN
            sigmoid_f := 4;
        ELSIF x =- 12742 THEN
            sigmoid_f := 4;
        ELSIF x =- 12741 THEN
            sigmoid_f := 4;
        ELSIF x =- 12740 THEN
            sigmoid_f := 4;
        ELSIF x =- 12739 THEN
            sigmoid_f := 4;
        ELSIF x =- 12738 THEN
            sigmoid_f := 4;
        ELSIF x =- 12737 THEN
            sigmoid_f := 4;
        ELSIF x =- 12736 THEN
            sigmoid_f := 4;
        ELSIF x =- 12735 THEN
            sigmoid_f := 4;
        ELSIF x =- 12734 THEN
            sigmoid_f := 4;
        ELSIF x =- 12733 THEN
            sigmoid_f := 4;
        ELSIF x =- 12732 THEN
            sigmoid_f := 4;
        ELSIF x =- 12731 THEN
            sigmoid_f := 4;
        ELSIF x =- 12730 THEN
            sigmoid_f := 4;
        ELSIF x =- 12729 THEN
            sigmoid_f := 4;
        ELSIF x =- 12728 THEN
            sigmoid_f := 4;
        ELSIF x =- 12727 THEN
            sigmoid_f := 4;
        ELSIF x =- 12726 THEN
            sigmoid_f := 4;
        ELSIF x =- 12725 THEN
            sigmoid_f := 4;
        ELSIF x =- 12724 THEN
            sigmoid_f := 4;
        ELSIF x =- 12723 THEN
            sigmoid_f := 4;
        ELSIF x =- 12722 THEN
            sigmoid_f := 4;
        ELSIF x =- 12721 THEN
            sigmoid_f := 4;
        ELSIF x =- 12720 THEN
            sigmoid_f := 4;
        ELSIF x =- 12719 THEN
            sigmoid_f := 4;
        ELSIF x =- 12718 THEN
            sigmoid_f := 4;
        ELSIF x =- 12717 THEN
            sigmoid_f := 4;
        ELSIF x =- 12716 THEN
            sigmoid_f := 4;
        ELSIF x =- 12715 THEN
            sigmoid_f := 4;
        ELSIF x =- 12714 THEN
            sigmoid_f := 4;
        ELSIF x =- 12713 THEN
            sigmoid_f := 4;
        ELSIF x =- 12712 THEN
            sigmoid_f := 4;
        ELSIF x =- 12711 THEN
            sigmoid_f := 4;
        ELSIF x =- 12710 THEN
            sigmoid_f := 4;
        ELSIF x =- 12709 THEN
            sigmoid_f := 4;
        ELSIF x =- 12708 THEN
            sigmoid_f := 4;
        ELSIF x =- 12707 THEN
            sigmoid_f := 4;
        ELSIF x =- 12706 THEN
            sigmoid_f := 4;
        ELSIF x =- 12705 THEN
            sigmoid_f := 4;
        ELSIF x =- 12704 THEN
            sigmoid_f := 4;
        ELSIF x =- 12703 THEN
            sigmoid_f := 4;
        ELSIF x =- 12702 THEN
            sigmoid_f := 4;
        ELSIF x =- 12701 THEN
            sigmoid_f := 4;
        ELSIF x =- 12700 THEN
            sigmoid_f := 4;
        ELSIF x =- 12699 THEN
            sigmoid_f := 4;
        ELSIF x =- 12698 THEN
            sigmoid_f := 4;
        ELSIF x =- 12697 THEN
            sigmoid_f := 4;
        ELSIF x =- 12696 THEN
            sigmoid_f := 4;
        ELSIF x =- 12695 THEN
            sigmoid_f := 4;
        ELSIF x =- 12694 THEN
            sigmoid_f := 4;
        ELSIF x =- 12693 THEN
            sigmoid_f := 4;
        ELSIF x =- 12692 THEN
            sigmoid_f := 4;
        ELSIF x =- 12691 THEN
            sigmoid_f := 4;
        ELSIF x =- 12690 THEN
            sigmoid_f := 4;
        ELSIF x =- 12689 THEN
            sigmoid_f := 4;
        ELSIF x =- 12688 THEN
            sigmoid_f := 4;
        ELSIF x =- 12687 THEN
            sigmoid_f := 4;
        ELSIF x =- 12686 THEN
            sigmoid_f := 4;
        ELSIF x =- 12685 THEN
            sigmoid_f := 4;
        ELSIF x =- 12684 THEN
            sigmoid_f := 4;
        ELSIF x =- 12683 THEN
            sigmoid_f := 4;
        ELSIF x =- 12682 THEN
            sigmoid_f := 4;
        ELSIF x =- 12681 THEN
            sigmoid_f := 4;
        ELSIF x =- 12680 THEN
            sigmoid_f := 4;
        ELSIF x =- 12679 THEN
            sigmoid_f := 4;
        ELSIF x =- 12678 THEN
            sigmoid_f := 4;
        ELSIF x =- 12677 THEN
            sigmoid_f := 4;
        ELSIF x =- 12676 THEN
            sigmoid_f := 4;
        ELSIF x =- 12675 THEN
            sigmoid_f := 4;
        ELSIF x =- 12674 THEN
            sigmoid_f := 4;
        ELSIF x =- 12673 THEN
            sigmoid_f := 4;
        ELSIF x =- 12672 THEN
            sigmoid_f := 4;
        ELSIF x =- 12671 THEN
            sigmoid_f := 4;
        ELSIF x =- 12670 THEN
            sigmoid_f := 4;
        ELSIF x =- 12669 THEN
            sigmoid_f := 4;
        ELSIF x =- 12668 THEN
            sigmoid_f := 4;
        ELSIF x =- 12667 THEN
            sigmoid_f := 4;
        ELSIF x =- 12666 THEN
            sigmoid_f := 4;
        ELSIF x =- 12665 THEN
            sigmoid_f := 4;
        ELSIF x =- 12664 THEN
            sigmoid_f := 4;
        ELSIF x =- 12663 THEN
            sigmoid_f := 4;
        ELSIF x =- 12662 THEN
            sigmoid_f := 4;
        ELSIF x =- 12661 THEN
            sigmoid_f := 4;
        ELSIF x =- 12660 THEN
            sigmoid_f := 4;
        ELSIF x =- 12659 THEN
            sigmoid_f := 4;
        ELSIF x =- 12658 THEN
            sigmoid_f := 4;
        ELSIF x =- 12657 THEN
            sigmoid_f := 4;
        ELSIF x =- 12656 THEN
            sigmoid_f := 4;
        ELSIF x =- 12655 THEN
            sigmoid_f := 4;
        ELSIF x =- 12654 THEN
            sigmoid_f := 4;
        ELSIF x =- 12653 THEN
            sigmoid_f := 4;
        ELSIF x =- 12652 THEN
            sigmoid_f := 4;
        ELSIF x =- 12651 THEN
            sigmoid_f := 4;
        ELSIF x =- 12650 THEN
            sigmoid_f := 4;
        ELSIF x =- 12649 THEN
            sigmoid_f := 4;
        ELSIF x =- 12648 THEN
            sigmoid_f := 4;
        ELSIF x =- 12647 THEN
            sigmoid_f := 4;
        ELSIF x =- 12646 THEN
            sigmoid_f := 4;
        ELSIF x =- 12645 THEN
            sigmoid_f := 4;
        ELSIF x =- 12644 THEN
            sigmoid_f := 4;
        ELSIF x =- 12643 THEN
            sigmoid_f := 4;
        ELSIF x =- 12642 THEN
            sigmoid_f := 4;
        ELSIF x =- 12641 THEN
            sigmoid_f := 4;
        ELSIF x =- 12640 THEN
            sigmoid_f := 4;
        ELSIF x =- 12639 THEN
            sigmoid_f := 4;
        ELSIF x =- 12638 THEN
            sigmoid_f := 4;
        ELSIF x =- 12637 THEN
            sigmoid_f := 4;
        ELSIF x =- 12636 THEN
            sigmoid_f := 4;
        ELSIF x =- 12635 THEN
            sigmoid_f := 4;
        ELSIF x =- 12634 THEN
            sigmoid_f := 4;
        ELSIF x =- 12633 THEN
            sigmoid_f := 4;
        ELSIF x =- 12632 THEN
            sigmoid_f := 4;
        ELSIF x =- 12631 THEN
            sigmoid_f := 4;
        ELSIF x =- 12630 THEN
            sigmoid_f := 4;
        ELSIF x =- 12629 THEN
            sigmoid_f := 4;
        ELSIF x =- 12628 THEN
            sigmoid_f := 4;
        ELSIF x =- 12627 THEN
            sigmoid_f := 4;
        ELSIF x =- 12626 THEN
            sigmoid_f := 4;
        ELSIF x =- 12625 THEN
            sigmoid_f := 4;
        ELSIF x =- 12624 THEN
            sigmoid_f := 4;
        ELSIF x =- 12623 THEN
            sigmoid_f := 4;
        ELSIF x =- 12622 THEN
            sigmoid_f := 4;
        ELSIF x =- 12621 THEN
            sigmoid_f := 4;
        ELSIF x =- 12620 THEN
            sigmoid_f := 4;
        ELSIF x =- 12619 THEN
            sigmoid_f := 4;
        ELSIF x =- 12618 THEN
            sigmoid_f := 4;
        ELSIF x =- 12617 THEN
            sigmoid_f := 4;
        ELSIF x =- 12616 THEN
            sigmoid_f := 4;
        ELSIF x =- 12615 THEN
            sigmoid_f := 4;
        ELSIF x =- 12614 THEN
            sigmoid_f := 4;
        ELSIF x =- 12613 THEN
            sigmoid_f := 4;
        ELSIF x =- 12612 THEN
            sigmoid_f := 4;
        ELSIF x =- 12611 THEN
            sigmoid_f := 4;
        ELSIF x =- 12610 THEN
            sigmoid_f := 4;
        ELSIF x =- 12609 THEN
            sigmoid_f := 4;
        ELSIF x =- 12608 THEN
            sigmoid_f := 4;
        ELSIF x =- 12607 THEN
            sigmoid_f := 4;
        ELSIF x =- 12606 THEN
            sigmoid_f := 4;
        ELSIF x =- 12605 THEN
            sigmoid_f := 4;
        ELSIF x =- 12604 THEN
            sigmoid_f := 4;
        ELSIF x =- 12603 THEN
            sigmoid_f := 4;
        ELSIF x =- 12602 THEN
            sigmoid_f := 4;
        ELSIF x =- 12601 THEN
            sigmoid_f := 4;
        ELSIF x =- 12600 THEN
            sigmoid_f := 4;
        ELSIF x =- 12599 THEN
            sigmoid_f := 4;
        ELSIF x =- 12598 THEN
            sigmoid_f := 4;
        ELSIF x =- 12597 THEN
            sigmoid_f := 4;
        ELSIF x =- 12596 THEN
            sigmoid_f := 4;
        ELSIF x =- 12595 THEN
            sigmoid_f := 4;
        ELSIF x =- 12594 THEN
            sigmoid_f := 4;
        ELSIF x =- 12593 THEN
            sigmoid_f := 4;
        ELSIF x =- 12592 THEN
            sigmoid_f := 4;
        ELSIF x =- 12591 THEN
            sigmoid_f := 4;
        ELSIF x =- 12590 THEN
            sigmoid_f := 4;
        ELSIF x =- 12589 THEN
            sigmoid_f := 4;
        ELSIF x =- 12588 THEN
            sigmoid_f := 4;
        ELSIF x =- 12587 THEN
            sigmoid_f := 4;
        ELSIF x =- 12586 THEN
            sigmoid_f := 4;
        ELSIF x =- 12585 THEN
            sigmoid_f := 4;
        ELSIF x =- 12584 THEN
            sigmoid_f := 4;
        ELSIF x =- 12583 THEN
            sigmoid_f := 4;
        ELSIF x =- 12582 THEN
            sigmoid_f := 4;
        ELSIF x =- 12581 THEN
            sigmoid_f := 4;
        ELSIF x =- 12580 THEN
            sigmoid_f := 4;
        ELSIF x =- 12579 THEN
            sigmoid_f := 4;
        ELSIF x =- 12578 THEN
            sigmoid_f := 4;
        ELSIF x =- 12577 THEN
            sigmoid_f := 4;
        ELSIF x =- 12576 THEN
            sigmoid_f := 4;
        ELSIF x =- 12575 THEN
            sigmoid_f := 4;
        ELSIF x =- 12574 THEN
            sigmoid_f := 4;
        ELSIF x =- 12573 THEN
            sigmoid_f := 4;
        ELSIF x =- 12572 THEN
            sigmoid_f := 4;
        ELSIF x =- 12571 THEN
            sigmoid_f := 4;
        ELSIF x =- 12570 THEN
            sigmoid_f := 4;
        ELSIF x =- 12569 THEN
            sigmoid_f := 4;
        ELSIF x =- 12568 THEN
            sigmoid_f := 4;
        ELSIF x =- 12567 THEN
            sigmoid_f := 4;
        ELSIF x =- 12566 THEN
            sigmoid_f := 4;
        ELSIF x =- 12565 THEN
            sigmoid_f := 4;
        ELSIF x =- 12564 THEN
            sigmoid_f := 4;
        ELSIF x =- 12563 THEN
            sigmoid_f := 4;
        ELSIF x =- 12562 THEN
            sigmoid_f := 4;
        ELSIF x =- 12561 THEN
            sigmoid_f := 4;
        ELSIF x =- 12560 THEN
            sigmoid_f := 4;
        ELSIF x =- 12559 THEN
            sigmoid_f := 4;
        ELSIF x =- 12558 THEN
            sigmoid_f := 4;
        ELSIF x =- 12557 THEN
            sigmoid_f := 4;
        ELSIF x =- 12556 THEN
            sigmoid_f := 4;
        ELSIF x =- 12555 THEN
            sigmoid_f := 4;
        ELSIF x =- 12554 THEN
            sigmoid_f := 4;
        ELSIF x =- 12553 THEN
            sigmoid_f := 4;
        ELSIF x =- 12552 THEN
            sigmoid_f := 4;
        ELSIF x =- 12551 THEN
            sigmoid_f := 4;
        ELSIF x =- 12550 THEN
            sigmoid_f := 4;
        ELSIF x =- 12549 THEN
            sigmoid_f := 4;
        ELSIF x =- 12548 THEN
            sigmoid_f := 4;
        ELSIF x =- 12547 THEN
            sigmoid_f := 4;
        ELSIF x =- 12546 THEN
            sigmoid_f := 4;
        ELSIF x =- 12545 THEN
            sigmoid_f := 4;
        ELSIF x =- 12544 THEN
            sigmoid_f := 4;
        ELSIF x =- 12543 THEN
            sigmoid_f := 4;
        ELSIF x =- 12542 THEN
            sigmoid_f := 4;
        ELSIF x =- 12541 THEN
            sigmoid_f := 4;
        ELSIF x =- 12540 THEN
            sigmoid_f := 4;
        ELSIF x =- 12539 THEN
            sigmoid_f := 4;
        ELSIF x =- 12538 THEN
            sigmoid_f := 4;
        ELSIF x =- 12537 THEN
            sigmoid_f := 4;
        ELSIF x =- 12536 THEN
            sigmoid_f := 4;
        ELSIF x =- 12535 THEN
            sigmoid_f := 4;
        ELSIF x =- 12534 THEN
            sigmoid_f := 4;
        ELSIF x =- 12533 THEN
            sigmoid_f := 4;
        ELSIF x =- 12532 THEN
            sigmoid_f := 4;
        ELSIF x =- 12531 THEN
            sigmoid_f := 4;
        ELSIF x =- 12530 THEN
            sigmoid_f := 4;
        ELSIF x =- 12529 THEN
            sigmoid_f := 4;
        ELSIF x =- 12528 THEN
            sigmoid_f := 4;
        ELSIF x =- 12527 THEN
            sigmoid_f := 4;
        ELSIF x =- 12526 THEN
            sigmoid_f := 4;
        ELSIF x =- 12525 THEN
            sigmoid_f := 4;
        ELSIF x =- 12524 THEN
            sigmoid_f := 4;
        ELSIF x =- 12523 THEN
            sigmoid_f := 4;
        ELSIF x =- 12522 THEN
            sigmoid_f := 4;
        ELSIF x =- 12521 THEN
            sigmoid_f := 4;
        ELSIF x =- 12520 THEN
            sigmoid_f := 4;
        ELSIF x =- 12519 THEN
            sigmoid_f := 4;
        ELSIF x =- 12518 THEN
            sigmoid_f := 4;
        ELSIF x =- 12517 THEN
            sigmoid_f := 4;
        ELSIF x =- 12516 THEN
            sigmoid_f := 4;
        ELSIF x =- 12515 THEN
            sigmoid_f := 4;
        ELSIF x =- 12514 THEN
            sigmoid_f := 4;
        ELSIF x =- 12513 THEN
            sigmoid_f := 4;
        ELSIF x =- 12512 THEN
            sigmoid_f := 4;
        ELSIF x =- 12511 THEN
            sigmoid_f := 4;
        ELSIF x =- 12510 THEN
            sigmoid_f := 4;
        ELSIF x =- 12509 THEN
            sigmoid_f := 4;
        ELSIF x =- 12508 THEN
            sigmoid_f := 4;
        ELSIF x =- 12507 THEN
            sigmoid_f := 4;
        ELSIF x =- 12506 THEN
            sigmoid_f := 4;
        ELSIF x =- 12505 THEN
            sigmoid_f := 4;
        ELSIF x =- 12504 THEN
            sigmoid_f := 4;
        ELSIF x =- 12503 THEN
            sigmoid_f := 4;
        ELSIF x =- 12502 THEN
            sigmoid_f := 4;
        ELSIF x =- 12501 THEN
            sigmoid_f := 4;
        ELSIF x =- 12500 THEN
            sigmoid_f := 4;
        ELSIF x =- 12499 THEN
            sigmoid_f := 4;
        ELSIF x =- 12498 THEN
            sigmoid_f := 4;
        ELSIF x =- 12497 THEN
            sigmoid_f := 4;
        ELSIF x =- 12496 THEN
            sigmoid_f := 4;
        ELSIF x =- 12495 THEN
            sigmoid_f := 4;
        ELSIF x =- 12494 THEN
            sigmoid_f := 4;
        ELSIF x =- 12493 THEN
            sigmoid_f := 4;
        ELSIF x =- 12492 THEN
            sigmoid_f := 4;
        ELSIF x =- 12491 THEN
            sigmoid_f := 4;
        ELSIF x =- 12490 THEN
            sigmoid_f := 4;
        ELSIF x =- 12489 THEN
            sigmoid_f := 4;
        ELSIF x =- 12488 THEN
            sigmoid_f := 4;
        ELSIF x =- 12487 THEN
            sigmoid_f := 4;
        ELSIF x =- 12486 THEN
            sigmoid_f := 4;
        ELSIF x =- 12485 THEN
            sigmoid_f := 4;
        ELSIF x =- 12484 THEN
            sigmoid_f := 4;
        ELSIF x =- 12483 THEN
            sigmoid_f := 4;
        ELSIF x =- 12482 THEN
            sigmoid_f := 4;
        ELSIF x =- 12481 THEN
            sigmoid_f := 4;
        ELSIF x =- 12480 THEN
            sigmoid_f := 4;
        ELSIF x =- 12479 THEN
            sigmoid_f := 4;
        ELSIF x =- 12478 THEN
            sigmoid_f := 4;
        ELSIF x =- 12477 THEN
            sigmoid_f := 4;
        ELSIF x =- 12476 THEN
            sigmoid_f := 4;
        ELSIF x =- 12475 THEN
            sigmoid_f := 4;
        ELSIF x =- 12474 THEN
            sigmoid_f := 4;
        ELSIF x =- 12473 THEN
            sigmoid_f := 4;
        ELSIF x =- 12472 THEN
            sigmoid_f := 4;
        ELSIF x =- 12471 THEN
            sigmoid_f := 4;
        ELSIF x =- 12470 THEN
            sigmoid_f := 4;
        ELSIF x =- 12469 THEN
            sigmoid_f := 4;
        ELSIF x =- 12468 THEN
            sigmoid_f := 4;
        ELSIF x =- 12467 THEN
            sigmoid_f := 4;
        ELSIF x =- 12466 THEN
            sigmoid_f := 4;
        ELSIF x =- 12465 THEN
            sigmoid_f := 4;
        ELSIF x =- 12464 THEN
            sigmoid_f := 4;
        ELSIF x =- 12463 THEN
            sigmoid_f := 4;
        ELSIF x =- 12462 THEN
            sigmoid_f := 4;
        ELSIF x =- 12461 THEN
            sigmoid_f := 4;
        ELSIF x =- 12460 THEN
            sigmoid_f := 4;
        ELSIF x =- 12459 THEN
            sigmoid_f := 4;
        ELSIF x =- 12458 THEN
            sigmoid_f := 4;
        ELSIF x =- 12457 THEN
            sigmoid_f := 4;
        ELSIF x =- 12456 THEN
            sigmoid_f := 4;
        ELSIF x =- 12455 THEN
            sigmoid_f := 4;
        ELSIF x =- 12454 THEN
            sigmoid_f := 4;
        ELSIF x =- 12453 THEN
            sigmoid_f := 4;
        ELSIF x =- 12452 THEN
            sigmoid_f := 4;
        ELSIF x =- 12451 THEN
            sigmoid_f := 4;
        ELSIF x =- 12450 THEN
            sigmoid_f := 4;
        ELSIF x =- 12449 THEN
            sigmoid_f := 4;
        ELSIF x =- 12448 THEN
            sigmoid_f := 4;
        ELSIF x =- 12447 THEN
            sigmoid_f := 4;
        ELSIF x =- 12446 THEN
            sigmoid_f := 4;
        ELSIF x =- 12445 THEN
            sigmoid_f := 4;
        ELSIF x =- 12444 THEN
            sigmoid_f := 4;
        ELSIF x =- 12443 THEN
            sigmoid_f := 4;
        ELSIF x =- 12442 THEN
            sigmoid_f := 4;
        ELSIF x =- 12441 THEN
            sigmoid_f := 4;
        ELSIF x =- 12440 THEN
            sigmoid_f := 4;
        ELSIF x =- 12439 THEN
            sigmoid_f := 4;
        ELSIF x =- 12438 THEN
            sigmoid_f := 4;
        ELSIF x =- 12437 THEN
            sigmoid_f := 4;
        ELSIF x =- 12436 THEN
            sigmoid_f := 4;
        ELSIF x =- 12435 THEN
            sigmoid_f := 4;
        ELSIF x =- 12434 THEN
            sigmoid_f := 4;
        ELSIF x =- 12433 THEN
            sigmoid_f := 4;
        ELSIF x =- 12432 THEN
            sigmoid_f := 4;
        ELSIF x =- 12431 THEN
            sigmoid_f := 4;
        ELSIF x =- 12430 THEN
            sigmoid_f := 4;
        ELSIF x =- 12429 THEN
            sigmoid_f := 4;
        ELSIF x =- 12428 THEN
            sigmoid_f := 4;
        ELSIF x =- 12427 THEN
            sigmoid_f := 4;
        ELSIF x =- 12426 THEN
            sigmoid_f := 4;
        ELSIF x =- 12425 THEN
            sigmoid_f := 4;
        ELSIF x =- 12424 THEN
            sigmoid_f := 4;
        ELSIF x =- 12423 THEN
            sigmoid_f := 4;
        ELSIF x =- 12422 THEN
            sigmoid_f := 4;
        ELSIF x =- 12421 THEN
            sigmoid_f := 4;
        ELSIF x =- 12420 THEN
            sigmoid_f := 4;
        ELSIF x =- 12419 THEN
            sigmoid_f := 4;
        ELSIF x =- 12418 THEN
            sigmoid_f := 4;
        ELSIF x =- 12417 THEN
            sigmoid_f := 4;
        ELSIF x =- 12416 THEN
            sigmoid_f := 4;
        ELSIF x =- 12415 THEN
            sigmoid_f := 4;
        ELSIF x =- 12414 THEN
            sigmoid_f := 4;
        ELSIF x =- 12413 THEN
            sigmoid_f := 4;
        ELSIF x =- 12412 THEN
            sigmoid_f := 4;
        ELSIF x =- 12411 THEN
            sigmoid_f := 4;
        ELSIF x =- 12410 THEN
            sigmoid_f := 4;
        ELSIF x =- 12409 THEN
            sigmoid_f := 4;
        ELSIF x =- 12408 THEN
            sigmoid_f := 4;
        ELSIF x =- 12407 THEN
            sigmoid_f := 4;
        ELSIF x =- 12406 THEN
            sigmoid_f := 4;
        ELSIF x =- 12405 THEN
            sigmoid_f := 4;
        ELSIF x =- 12404 THEN
            sigmoid_f := 4;
        ELSIF x =- 12403 THEN
            sigmoid_f := 4;
        ELSIF x =- 12402 THEN
            sigmoid_f := 4;
        ELSIF x =- 12401 THEN
            sigmoid_f := 4;
        ELSIF x =- 12400 THEN
            sigmoid_f := 4;
        ELSIF x =- 12399 THEN
            sigmoid_f := 4;
        ELSIF x =- 12398 THEN
            sigmoid_f := 4;
        ELSIF x =- 12397 THEN
            sigmoid_f := 4;
        ELSIF x =- 12396 THEN
            sigmoid_f := 4;
        ELSIF x =- 12395 THEN
            sigmoid_f := 4;
        ELSIF x =- 12394 THEN
            sigmoid_f := 4;
        ELSIF x =- 12393 THEN
            sigmoid_f := 4;
        ELSIF x =- 12392 THEN
            sigmoid_f := 4;
        ELSIF x =- 12391 THEN
            sigmoid_f := 4;
        ELSIF x =- 12390 THEN
            sigmoid_f := 4;
        ELSIF x =- 12389 THEN
            sigmoid_f := 4;
        ELSIF x =- 12388 THEN
            sigmoid_f := 4;
        ELSIF x =- 12387 THEN
            sigmoid_f := 4;
        ELSIF x =- 12386 THEN
            sigmoid_f := 4;
        ELSIF x =- 12385 THEN
            sigmoid_f := 4;
        ELSIF x =- 12384 THEN
            sigmoid_f := 4;
        ELSIF x =- 12383 THEN
            sigmoid_f := 4;
        ELSIF x =- 12382 THEN
            sigmoid_f := 4;
        ELSIF x =- 12381 THEN
            sigmoid_f := 4;
        ELSIF x =- 12380 THEN
            sigmoid_f := 4;
        ELSIF x =- 12379 THEN
            sigmoid_f := 4;
        ELSIF x =- 12378 THEN
            sigmoid_f := 4;
        ELSIF x =- 12377 THEN
            sigmoid_f := 4;
        ELSIF x =- 12376 THEN
            sigmoid_f := 4;
        ELSIF x =- 12375 THEN
            sigmoid_f := 4;
        ELSIF x =- 12374 THEN
            sigmoid_f := 4;
        ELSIF x =- 12373 THEN
            sigmoid_f := 4;
        ELSIF x =- 12372 THEN
            sigmoid_f := 4;
        ELSIF x =- 12371 THEN
            sigmoid_f := 4;
        ELSIF x =- 12370 THEN
            sigmoid_f := 4;
        ELSIF x =- 12369 THEN
            sigmoid_f := 4;
        ELSIF x =- 12368 THEN
            sigmoid_f := 4;
        ELSIF x =- 12367 THEN
            sigmoid_f := 4;
        ELSIF x =- 12366 THEN
            sigmoid_f := 4;
        ELSIF x =- 12365 THEN
            sigmoid_f := 4;
        ELSIF x =- 12364 THEN
            sigmoid_f := 4;
        ELSIF x =- 12363 THEN
            sigmoid_f := 4;
        ELSIF x =- 12362 THEN
            sigmoid_f := 4;
        ELSIF x =- 12361 THEN
            sigmoid_f := 4;
        ELSIF x =- 12360 THEN
            sigmoid_f := 4;
        ELSIF x =- 12359 THEN
            sigmoid_f := 4;
        ELSIF x =- 12358 THEN
            sigmoid_f := 4;
        ELSIF x =- 12357 THEN
            sigmoid_f := 4;
        ELSIF x =- 12356 THEN
            sigmoid_f := 4;
        ELSIF x =- 12355 THEN
            sigmoid_f := 4;
        ELSIF x =- 12354 THEN
            sigmoid_f := 4;
        ELSIF x =- 12353 THEN
            sigmoid_f := 4;
        ELSIF x =- 12352 THEN
            sigmoid_f := 4;
        ELSIF x =- 12351 THEN
            sigmoid_f := 4;
        ELSIF x =- 12350 THEN
            sigmoid_f := 4;
        ELSIF x =- 12349 THEN
            sigmoid_f := 4;
        ELSIF x =- 12348 THEN
            sigmoid_f := 4;
        ELSIF x =- 12347 THEN
            sigmoid_f := 4;
        ELSIF x =- 12346 THEN
            sigmoid_f := 4;
        ELSIF x =- 12345 THEN
            sigmoid_f := 4;
        ELSIF x =- 12344 THEN
            sigmoid_f := 4;
        ELSIF x =- 12343 THEN
            sigmoid_f := 4;
        ELSIF x =- 12342 THEN
            sigmoid_f := 4;
        ELSIF x =- 12341 THEN
            sigmoid_f := 4;
        ELSIF x =- 12340 THEN
            sigmoid_f := 4;
        ELSIF x =- 12339 THEN
            sigmoid_f := 4;
        ELSIF x =- 12338 THEN
            sigmoid_f := 4;
        ELSIF x =- 12337 THEN
            sigmoid_f := 4;
        ELSIF x =- 12336 THEN
            sigmoid_f := 4;
        ELSIF x =- 12335 THEN
            sigmoid_f := 4;
        ELSIF x =- 12334 THEN
            sigmoid_f := 4;
        ELSIF x =- 12333 THEN
            sigmoid_f := 4;
        ELSIF x =- 12332 THEN
            sigmoid_f := 4;
        ELSIF x =- 12331 THEN
            sigmoid_f := 4;
        ELSIF x =- 12330 THEN
            sigmoid_f := 4;
        ELSIF x =- 12329 THEN
            sigmoid_f := 4;
        ELSIF x =- 12328 THEN
            sigmoid_f := 4;
        ELSIF x =- 12327 THEN
            sigmoid_f := 4;
        ELSIF x =- 12326 THEN
            sigmoid_f := 4;
        ELSIF x =- 12325 THEN
            sigmoid_f := 4;
        ELSIF x =- 12324 THEN
            sigmoid_f := 4;
        ELSIF x =- 12323 THEN
            sigmoid_f := 4;
        ELSIF x =- 12322 THEN
            sigmoid_f := 4;
        ELSIF x =- 12321 THEN
            sigmoid_f := 4;
        ELSIF x =- 12320 THEN
            sigmoid_f := 4;
        ELSIF x =- 12319 THEN
            sigmoid_f := 4;
        ELSIF x =- 12318 THEN
            sigmoid_f := 4;
        ELSIF x =- 12317 THEN
            sigmoid_f := 4;
        ELSIF x =- 12316 THEN
            sigmoid_f := 4;
        ELSIF x =- 12315 THEN
            sigmoid_f := 4;
        ELSIF x =- 12314 THEN
            sigmoid_f := 4;
        ELSIF x =- 12313 THEN
            sigmoid_f := 4;
        ELSIF x =- 12312 THEN
            sigmoid_f := 4;
        ELSIF x =- 12311 THEN
            sigmoid_f := 4;
        ELSIF x =- 12310 THEN
            sigmoid_f := 4;
        ELSIF x =- 12309 THEN
            sigmoid_f := 4;
        ELSIF x =- 12308 THEN
            sigmoid_f := 4;
        ELSIF x =- 12307 THEN
            sigmoid_f := 4;
        ELSIF x =- 12306 THEN
            sigmoid_f := 4;
        ELSIF x =- 12305 THEN
            sigmoid_f := 4;
        ELSIF x =- 12304 THEN
            sigmoid_f := 4;
        ELSIF x =- 12303 THEN
            sigmoid_f := 4;
        ELSIF x =- 12302 THEN
            sigmoid_f := 4;
        ELSIF x =- 12301 THEN
            sigmoid_f := 4;
        ELSIF x =- 12300 THEN
            sigmoid_f := 4;
        ELSIF x =- 12299 THEN
            sigmoid_f := 4;
        ELSIF x =- 12298 THEN
            sigmoid_f := 4;
        ELSIF x =- 12297 THEN
            sigmoid_f := 4;
        ELSIF x =- 12296 THEN
            sigmoid_f := 4;
        ELSIF x =- 12295 THEN
            sigmoid_f := 4;
        ELSIF x =- 12294 THEN
            sigmoid_f := 4;
        ELSIF x =- 12293 THEN
            sigmoid_f := 4;
        ELSIF x =- 12292 THEN
            sigmoid_f := 4;
        ELSIF x =- 12291 THEN
            sigmoid_f := 4;
        ELSIF x =- 12290 THEN
            sigmoid_f := 4;
        ELSIF x =- 12289 THEN
            sigmoid_f := 4;
        ELSIF x =- 12288 THEN
            sigmoid_f := 4;
        ELSIF x =- 12287 THEN
            sigmoid_f := 6;
        ELSIF x =- 12286 THEN
            sigmoid_f := 6;
        ELSIF x =- 12285 THEN
            sigmoid_f := 6;
        ELSIF x =- 12284 THEN
            sigmoid_f := 6;
        ELSIF x =- 12283 THEN
            sigmoid_f := 6;
        ELSIF x =- 12282 THEN
            sigmoid_f := 6;
        ELSIF x =- 12281 THEN
            sigmoid_f := 6;
        ELSIF x =- 12280 THEN
            sigmoid_f := 6;
        ELSIF x =- 12279 THEN
            sigmoid_f := 6;
        ELSIF x =- 12278 THEN
            sigmoid_f := 6;
        ELSIF x =- 12277 THEN
            sigmoid_f := 6;
        ELSIF x =- 12276 THEN
            sigmoid_f := 6;
        ELSIF x =- 12275 THEN
            sigmoid_f := 6;
        ELSIF x =- 12274 THEN
            sigmoid_f := 6;
        ELSIF x =- 12273 THEN
            sigmoid_f := 6;
        ELSIF x =- 12272 THEN
            sigmoid_f := 6;
        ELSIF x =- 12271 THEN
            sigmoid_f := 6;
        ELSIF x =- 12270 THEN
            sigmoid_f := 6;
        ELSIF x =- 12269 THEN
            sigmoid_f := 6;
        ELSIF x =- 12268 THEN
            sigmoid_f := 6;
        ELSIF x =- 12267 THEN
            sigmoid_f := 6;
        ELSIF x =- 12266 THEN
            sigmoid_f := 6;
        ELSIF x =- 12265 THEN
            sigmoid_f := 6;
        ELSIF x =- 12264 THEN
            sigmoid_f := 6;
        ELSIF x =- 12263 THEN
            sigmoid_f := 6;
        ELSIF x =- 12262 THEN
            sigmoid_f := 6;
        ELSIF x =- 12261 THEN
            sigmoid_f := 6;
        ELSIF x =- 12260 THEN
            sigmoid_f := 6;
        ELSIF x =- 12259 THEN
            sigmoid_f := 6;
        ELSIF x =- 12258 THEN
            sigmoid_f := 6;
        ELSIF x =- 12257 THEN
            sigmoid_f := 6;
        ELSIF x =- 12256 THEN
            sigmoid_f := 6;
        ELSIF x =- 12255 THEN
            sigmoid_f := 6;
        ELSIF x =- 12254 THEN
            sigmoid_f := 6;
        ELSIF x =- 12253 THEN
            sigmoid_f := 6;
        ELSIF x =- 12252 THEN
            sigmoid_f := 6;
        ELSIF x =- 12251 THEN
            sigmoid_f := 6;
        ELSIF x =- 12250 THEN
            sigmoid_f := 6;
        ELSIF x =- 12249 THEN
            sigmoid_f := 6;
        ELSIF x =- 12248 THEN
            sigmoid_f := 6;
        ELSIF x =- 12247 THEN
            sigmoid_f := 6;
        ELSIF x =- 12246 THEN
            sigmoid_f := 6;
        ELSIF x =- 12245 THEN
            sigmoid_f := 6;
        ELSIF x =- 12244 THEN
            sigmoid_f := 6;
        ELSIF x =- 12243 THEN
            sigmoid_f := 6;
        ELSIF x =- 12242 THEN
            sigmoid_f := 6;
        ELSIF x =- 12241 THEN
            sigmoid_f := 6;
        ELSIF x =- 12240 THEN
            sigmoid_f := 6;
        ELSIF x =- 12239 THEN
            sigmoid_f := 6;
        ELSIF x =- 12238 THEN
            sigmoid_f := 6;
        ELSIF x =- 12237 THEN
            sigmoid_f := 6;
        ELSIF x =- 12236 THEN
            sigmoid_f := 6;
        ELSIF x =- 12235 THEN
            sigmoid_f := 6;
        ELSIF x =- 12234 THEN
            sigmoid_f := 6;
        ELSIF x =- 12233 THEN
            sigmoid_f := 6;
        ELSIF x =- 12232 THEN
            sigmoid_f := 6;
        ELSIF x =- 12231 THEN
            sigmoid_f := 6;
        ELSIF x =- 12230 THEN
            sigmoid_f := 6;
        ELSIF x =- 12229 THEN
            sigmoid_f := 6;
        ELSIF x =- 12228 THEN
            sigmoid_f := 6;
        ELSIF x =- 12227 THEN
            sigmoid_f := 6;
        ELSIF x =- 12226 THEN
            sigmoid_f := 6;
        ELSIF x =- 12225 THEN
            sigmoid_f := 6;
        ELSIF x =- 12224 THEN
            sigmoid_f := 6;
        ELSIF x =- 12223 THEN
            sigmoid_f := 6;
        ELSIF x =- 12222 THEN
            sigmoid_f := 6;
        ELSIF x =- 12221 THEN
            sigmoid_f := 6;
        ELSIF x =- 12220 THEN
            sigmoid_f := 6;
        ELSIF x =- 12219 THEN
            sigmoid_f := 6;
        ELSIF x =- 12218 THEN
            sigmoid_f := 6;
        ELSIF x =- 12217 THEN
            sigmoid_f := 6;
        ELSIF x =- 12216 THEN
            sigmoid_f := 6;
        ELSIF x =- 12215 THEN
            sigmoid_f := 6;
        ELSIF x =- 12214 THEN
            sigmoid_f := 6;
        ELSIF x =- 12213 THEN
            sigmoid_f := 6;
        ELSIF x =- 12212 THEN
            sigmoid_f := 6;
        ELSIF x =- 12211 THEN
            sigmoid_f := 6;
        ELSIF x =- 12210 THEN
            sigmoid_f := 6;
        ELSIF x =- 12209 THEN
            sigmoid_f := 6;
        ELSIF x =- 12208 THEN
            sigmoid_f := 6;
        ELSIF x =- 12207 THEN
            sigmoid_f := 6;
        ELSIF x =- 12206 THEN
            sigmoid_f := 6;
        ELSIF x =- 12205 THEN
            sigmoid_f := 6;
        ELSIF x =- 12204 THEN
            sigmoid_f := 6;
        ELSIF x =- 12203 THEN
            sigmoid_f := 6;
        ELSIF x =- 12202 THEN
            sigmoid_f := 6;
        ELSIF x =- 12201 THEN
            sigmoid_f := 6;
        ELSIF x =- 12200 THEN
            sigmoid_f := 6;
        ELSIF x =- 12199 THEN
            sigmoid_f := 6;
        ELSIF x =- 12198 THEN
            sigmoid_f := 6;
        ELSIF x =- 12197 THEN
            sigmoid_f := 6;
        ELSIF x =- 12196 THEN
            sigmoid_f := 6;
        ELSIF x =- 12195 THEN
            sigmoid_f := 6;
        ELSIF x =- 12194 THEN
            sigmoid_f := 6;
        ELSIF x =- 12193 THEN
            sigmoid_f := 6;
        ELSIF x =- 12192 THEN
            sigmoid_f := 6;
        ELSIF x =- 12191 THEN
            sigmoid_f := 6;
        ELSIF x =- 12190 THEN
            sigmoid_f := 6;
        ELSIF x =- 12189 THEN
            sigmoid_f := 6;
        ELSIF x =- 12188 THEN
            sigmoid_f := 6;
        ELSIF x =- 12187 THEN
            sigmoid_f := 6;
        ELSIF x =- 12186 THEN
            sigmoid_f := 6;
        ELSIF x =- 12185 THEN
            sigmoid_f := 6;
        ELSIF x =- 12184 THEN
            sigmoid_f := 6;
        ELSIF x =- 12183 THEN
            sigmoid_f := 6;
        ELSIF x =- 12182 THEN
            sigmoid_f := 6;
        ELSIF x =- 12181 THEN
            sigmoid_f := 6;
        ELSIF x =- 12180 THEN
            sigmoid_f := 6;
        ELSIF x =- 12179 THEN
            sigmoid_f := 6;
        ELSIF x =- 12178 THEN
            sigmoid_f := 6;
        ELSIF x =- 12177 THEN
            sigmoid_f := 6;
        ELSIF x =- 12176 THEN
            sigmoid_f := 6;
        ELSIF x =- 12175 THEN
            sigmoid_f := 6;
        ELSIF x =- 12174 THEN
            sigmoid_f := 6;
        ELSIF x =- 12173 THEN
            sigmoid_f := 6;
        ELSIF x =- 12172 THEN
            sigmoid_f := 6;
        ELSIF x =- 12171 THEN
            sigmoid_f := 6;
        ELSIF x =- 12170 THEN
            sigmoid_f := 6;
        ELSIF x =- 12169 THEN
            sigmoid_f := 6;
        ELSIF x =- 12168 THEN
            sigmoid_f := 6;
        ELSIF x =- 12167 THEN
            sigmoid_f := 6;
        ELSIF x =- 12166 THEN
            sigmoid_f := 6;
        ELSIF x =- 12165 THEN
            sigmoid_f := 6;
        ELSIF x =- 12164 THEN
            sigmoid_f := 6;
        ELSIF x =- 12163 THEN
            sigmoid_f := 6;
        ELSIF x =- 12162 THEN
            sigmoid_f := 6;
        ELSIF x =- 12161 THEN
            sigmoid_f := 6;
        ELSIF x =- 12160 THEN
            sigmoid_f := 6;
        ELSIF x =- 12159 THEN
            sigmoid_f := 6;
        ELSIF x =- 12158 THEN
            sigmoid_f := 6;
        ELSIF x =- 12157 THEN
            sigmoid_f := 6;
        ELSIF x =- 12156 THEN
            sigmoid_f := 6;
        ELSIF x =- 12155 THEN
            sigmoid_f := 6;
        ELSIF x =- 12154 THEN
            sigmoid_f := 6;
        ELSIF x =- 12153 THEN
            sigmoid_f := 6;
        ELSIF x =- 12152 THEN
            sigmoid_f := 6;
        ELSIF x =- 12151 THEN
            sigmoid_f := 6;
        ELSIF x =- 12150 THEN
            sigmoid_f := 6;
        ELSIF x =- 12149 THEN
            sigmoid_f := 6;
        ELSIF x =- 12148 THEN
            sigmoid_f := 6;
        ELSIF x =- 12147 THEN
            sigmoid_f := 6;
        ELSIF x =- 12146 THEN
            sigmoid_f := 6;
        ELSIF x =- 12145 THEN
            sigmoid_f := 6;
        ELSIF x =- 12144 THEN
            sigmoid_f := 6;
        ELSIF x =- 12143 THEN
            sigmoid_f := 6;
        ELSIF x =- 12142 THEN
            sigmoid_f := 6;
        ELSIF x =- 12141 THEN
            sigmoid_f := 6;
        ELSIF x =- 12140 THEN
            sigmoid_f := 6;
        ELSIF x =- 12139 THEN
            sigmoid_f := 6;
        ELSIF x =- 12138 THEN
            sigmoid_f := 6;
        ELSIF x =- 12137 THEN
            sigmoid_f := 6;
        ELSIF x =- 12136 THEN
            sigmoid_f := 6;
        ELSIF x =- 12135 THEN
            sigmoid_f := 6;
        ELSIF x =- 12134 THEN
            sigmoid_f := 6;
        ELSIF x =- 12133 THEN
            sigmoid_f := 6;
        ELSIF x =- 12132 THEN
            sigmoid_f := 6;
        ELSIF x =- 12131 THEN
            sigmoid_f := 6;
        ELSIF x =- 12130 THEN
            sigmoid_f := 6;
        ELSIF x =- 12129 THEN
            sigmoid_f := 6;
        ELSIF x =- 12128 THEN
            sigmoid_f := 6;
        ELSIF x =- 12127 THEN
            sigmoid_f := 6;
        ELSIF x =- 12126 THEN
            sigmoid_f := 6;
        ELSIF x =- 12125 THEN
            sigmoid_f := 6;
        ELSIF x =- 12124 THEN
            sigmoid_f := 6;
        ELSIF x =- 12123 THEN
            sigmoid_f := 6;
        ELSIF x =- 12122 THEN
            sigmoid_f := 6;
        ELSIF x =- 12121 THEN
            sigmoid_f := 6;
        ELSIF x =- 12120 THEN
            sigmoid_f := 6;
        ELSIF x =- 12119 THEN
            sigmoid_f := 6;
        ELSIF x =- 12118 THEN
            sigmoid_f := 6;
        ELSIF x =- 12117 THEN
            sigmoid_f := 6;
        ELSIF x =- 12116 THEN
            sigmoid_f := 6;
        ELSIF x =- 12115 THEN
            sigmoid_f := 6;
        ELSIF x =- 12114 THEN
            sigmoid_f := 6;
        ELSIF x =- 12113 THEN
            sigmoid_f := 6;
        ELSIF x =- 12112 THEN
            sigmoid_f := 6;
        ELSIF x =- 12111 THEN
            sigmoid_f := 6;
        ELSIF x =- 12110 THEN
            sigmoid_f := 6;
        ELSIF x =- 12109 THEN
            sigmoid_f := 6;
        ELSIF x =- 12108 THEN
            sigmoid_f := 6;
        ELSIF x =- 12107 THEN
            sigmoid_f := 6;
        ELSIF x =- 12106 THEN
            sigmoid_f := 6;
        ELSIF x =- 12105 THEN
            sigmoid_f := 6;
        ELSIF x =- 12104 THEN
            sigmoid_f := 6;
        ELSIF x =- 12103 THEN
            sigmoid_f := 6;
        ELSIF x =- 12102 THEN
            sigmoid_f := 6;
        ELSIF x =- 12101 THEN
            sigmoid_f := 6;
        ELSIF x =- 12100 THEN
            sigmoid_f := 6;
        ELSIF x =- 12099 THEN
            sigmoid_f := 6;
        ELSIF x =- 12098 THEN
            sigmoid_f := 6;
        ELSIF x =- 12097 THEN
            sigmoid_f := 6;
        ELSIF x =- 12096 THEN
            sigmoid_f := 6;
        ELSIF x =- 12095 THEN
            sigmoid_f := 6;
        ELSIF x =- 12094 THEN
            sigmoid_f := 6;
        ELSIF x =- 12093 THEN
            sigmoid_f := 6;
        ELSIF x =- 12092 THEN
            sigmoid_f := 6;
        ELSIF x =- 12091 THEN
            sigmoid_f := 6;
        ELSIF x =- 12090 THEN
            sigmoid_f := 6;
        ELSIF x =- 12089 THEN
            sigmoid_f := 6;
        ELSIF x =- 12088 THEN
            sigmoid_f := 6;
        ELSIF x =- 12087 THEN
            sigmoid_f := 6;
        ELSIF x =- 12086 THEN
            sigmoid_f := 6;
        ELSIF x =- 12085 THEN
            sigmoid_f := 6;
        ELSIF x =- 12084 THEN
            sigmoid_f := 6;
        ELSIF x =- 12083 THEN
            sigmoid_f := 6;
        ELSIF x =- 12082 THEN
            sigmoid_f := 6;
        ELSIF x =- 12081 THEN
            sigmoid_f := 6;
        ELSIF x =- 12080 THEN
            sigmoid_f := 6;
        ELSIF x =- 12079 THEN
            sigmoid_f := 6;
        ELSIF x =- 12078 THEN
            sigmoid_f := 6;
        ELSIF x =- 12077 THEN
            sigmoid_f := 6;
        ELSIF x =- 12076 THEN
            sigmoid_f := 6;
        ELSIF x =- 12075 THEN
            sigmoid_f := 6;
        ELSIF x =- 12074 THEN
            sigmoid_f := 6;
        ELSIF x =- 12073 THEN
            sigmoid_f := 6;
        ELSIF x =- 12072 THEN
            sigmoid_f := 6;
        ELSIF x =- 12071 THEN
            sigmoid_f := 6;
        ELSIF x =- 12070 THEN
            sigmoid_f := 6;
        ELSIF x =- 12069 THEN
            sigmoid_f := 6;
        ELSIF x =- 12068 THEN
            sigmoid_f := 6;
        ELSIF x =- 12067 THEN
            sigmoid_f := 6;
        ELSIF x =- 12066 THEN
            sigmoid_f := 6;
        ELSIF x =- 12065 THEN
            sigmoid_f := 6;
        ELSIF x =- 12064 THEN
            sigmoid_f := 6;
        ELSIF x =- 12063 THEN
            sigmoid_f := 6;
        ELSIF x =- 12062 THEN
            sigmoid_f := 6;
        ELSIF x =- 12061 THEN
            sigmoid_f := 6;
        ELSIF x =- 12060 THEN
            sigmoid_f := 6;
        ELSIF x =- 12059 THEN
            sigmoid_f := 6;
        ELSIF x =- 12058 THEN
            sigmoid_f := 6;
        ELSIF x =- 12057 THEN
            sigmoid_f := 6;
        ELSIF x =- 12056 THEN
            sigmoid_f := 6;
        ELSIF x =- 12055 THEN
            sigmoid_f := 6;
        ELSIF x =- 12054 THEN
            sigmoid_f := 6;
        ELSIF x =- 12053 THEN
            sigmoid_f := 6;
        ELSIF x =- 12052 THEN
            sigmoid_f := 6;
        ELSIF x =- 12051 THEN
            sigmoid_f := 6;
        ELSIF x =- 12050 THEN
            sigmoid_f := 6;
        ELSIF x =- 12049 THEN
            sigmoid_f := 6;
        ELSIF x =- 12048 THEN
            sigmoid_f := 6;
        ELSIF x =- 12047 THEN
            sigmoid_f := 6;
        ELSIF x =- 12046 THEN
            sigmoid_f := 6;
        ELSIF x =- 12045 THEN
            sigmoid_f := 6;
        ELSIF x =- 12044 THEN
            sigmoid_f := 6;
        ELSIF x =- 12043 THEN
            sigmoid_f := 6;
        ELSIF x =- 12042 THEN
            sigmoid_f := 6;
        ELSIF x =- 12041 THEN
            sigmoid_f := 6;
        ELSIF x =- 12040 THEN
            sigmoid_f := 6;
        ELSIF x =- 12039 THEN
            sigmoid_f := 6;
        ELSIF x =- 12038 THEN
            sigmoid_f := 6;
        ELSIF x =- 12037 THEN
            sigmoid_f := 6;
        ELSIF x =- 12036 THEN
            sigmoid_f := 6;
        ELSIF x =- 12035 THEN
            sigmoid_f := 6;
        ELSIF x =- 12034 THEN
            sigmoid_f := 6;
        ELSIF x =- 12033 THEN
            sigmoid_f := 6;
        ELSIF x =- 12032 THEN
            sigmoid_f := 6;
        ELSIF x =- 12031 THEN
            sigmoid_f := 6;
        ELSIF x =- 12030 THEN
            sigmoid_f := 6;
        ELSIF x =- 12029 THEN
            sigmoid_f := 6;
        ELSIF x =- 12028 THEN
            sigmoid_f := 6;
        ELSIF x =- 12027 THEN
            sigmoid_f := 6;
        ELSIF x =- 12026 THEN
            sigmoid_f := 6;
        ELSIF x =- 12025 THEN
            sigmoid_f := 6;
        ELSIF x =- 12024 THEN
            sigmoid_f := 6;
        ELSIF x =- 12023 THEN
            sigmoid_f := 6;
        ELSIF x =- 12022 THEN
            sigmoid_f := 6;
        ELSIF x =- 12021 THEN
            sigmoid_f := 6;
        ELSIF x =- 12020 THEN
            sigmoid_f := 6;
        ELSIF x =- 12019 THEN
            sigmoid_f := 6;
        ELSIF x =- 12018 THEN
            sigmoid_f := 6;
        ELSIF x =- 12017 THEN
            sigmoid_f := 6;
        ELSIF x =- 12016 THEN
            sigmoid_f := 6;
        ELSIF x =- 12015 THEN
            sigmoid_f := 6;
        ELSIF x =- 12014 THEN
            sigmoid_f := 6;
        ELSIF x =- 12013 THEN
            sigmoid_f := 6;
        ELSIF x =- 12012 THEN
            sigmoid_f := 6;
        ELSIF x =- 12011 THEN
            sigmoid_f := 6;
        ELSIF x =- 12010 THEN
            sigmoid_f := 6;
        ELSIF x =- 12009 THEN
            sigmoid_f := 6;
        ELSIF x =- 12008 THEN
            sigmoid_f := 6;
        ELSIF x =- 12007 THEN
            sigmoid_f := 6;
        ELSIF x =- 12006 THEN
            sigmoid_f := 6;
        ELSIF x =- 12005 THEN
            sigmoid_f := 6;
        ELSIF x =- 12004 THEN
            sigmoid_f := 6;
        ELSIF x =- 12003 THEN
            sigmoid_f := 6;
        ELSIF x =- 12002 THEN
            sigmoid_f := 6;
        ELSIF x =- 12001 THEN
            sigmoid_f := 6;
        ELSIF x =- 12000 THEN
            sigmoid_f := 6;
        ELSIF x =- 11999 THEN
            sigmoid_f := 6;
        ELSIF x =- 11998 THEN
            sigmoid_f := 6;
        ELSIF x =- 11997 THEN
            sigmoid_f := 6;
        ELSIF x =- 11996 THEN
            sigmoid_f := 6;
        ELSIF x =- 11995 THEN
            sigmoid_f := 6;
        ELSIF x =- 11994 THEN
            sigmoid_f := 6;
        ELSIF x =- 11993 THEN
            sigmoid_f := 6;
        ELSIF x =- 11992 THEN
            sigmoid_f := 6;
        ELSIF x =- 11991 THEN
            sigmoid_f := 6;
        ELSIF x =- 11990 THEN
            sigmoid_f := 6;
        ELSIF x =- 11989 THEN
            sigmoid_f := 6;
        ELSIF x =- 11988 THEN
            sigmoid_f := 6;
        ELSIF x =- 11987 THEN
            sigmoid_f := 6;
        ELSIF x =- 11986 THEN
            sigmoid_f := 6;
        ELSIF x =- 11985 THEN
            sigmoid_f := 6;
        ELSIF x =- 11984 THEN
            sigmoid_f := 6;
        ELSIF x =- 11983 THEN
            sigmoid_f := 6;
        ELSIF x =- 11982 THEN
            sigmoid_f := 6;
        ELSIF x =- 11981 THEN
            sigmoid_f := 6;
        ELSIF x =- 11980 THEN
            sigmoid_f := 6;
        ELSIF x =- 11979 THEN
            sigmoid_f := 6;
        ELSIF x =- 11978 THEN
            sigmoid_f := 6;
        ELSIF x =- 11977 THEN
            sigmoid_f := 6;
        ELSIF x =- 11976 THEN
            sigmoid_f := 6;
        ELSIF x =- 11975 THEN
            sigmoid_f := 6;
        ELSIF x =- 11974 THEN
            sigmoid_f := 6;
        ELSIF x =- 11973 THEN
            sigmoid_f := 6;
        ELSIF x =- 11972 THEN
            sigmoid_f := 6;
        ELSIF x =- 11971 THEN
            sigmoid_f := 6;
        ELSIF x =- 11970 THEN
            sigmoid_f := 6;
        ELSIF x =- 11969 THEN
            sigmoid_f := 6;
        ELSIF x =- 11968 THEN
            sigmoid_f := 6;
        ELSIF x =- 11967 THEN
            sigmoid_f := 6;
        ELSIF x =- 11966 THEN
            sigmoid_f := 6;
        ELSIF x =- 11965 THEN
            sigmoid_f := 6;
        ELSIF x =- 11964 THEN
            sigmoid_f := 6;
        ELSIF x =- 11963 THEN
            sigmoid_f := 6;
        ELSIF x =- 11962 THEN
            sigmoid_f := 6;
        ELSIF x =- 11961 THEN
            sigmoid_f := 6;
        ELSIF x =- 11960 THEN
            sigmoid_f := 6;
        ELSIF x =- 11959 THEN
            sigmoid_f := 6;
        ELSIF x =- 11958 THEN
            sigmoid_f := 6;
        ELSIF x =- 11957 THEN
            sigmoid_f := 6;
        ELSIF x =- 11956 THEN
            sigmoid_f := 6;
        ELSIF x =- 11955 THEN
            sigmoid_f := 6;
        ELSIF x =- 11954 THEN
            sigmoid_f := 6;
        ELSIF x =- 11953 THEN
            sigmoid_f := 6;
        ELSIF x =- 11952 THEN
            sigmoid_f := 6;
        ELSIF x =- 11951 THEN
            sigmoid_f := 6;
        ELSIF x =- 11950 THEN
            sigmoid_f := 6;
        ELSIF x =- 11949 THEN
            sigmoid_f := 6;
        ELSIF x =- 11948 THEN
            sigmoid_f := 6;
        ELSIF x =- 11947 THEN
            sigmoid_f := 6;
        ELSIF x =- 11946 THEN
            sigmoid_f := 6;
        ELSIF x =- 11945 THEN
            sigmoid_f := 6;
        ELSIF x =- 11944 THEN
            sigmoid_f := 6;
        ELSIF x =- 11943 THEN
            sigmoid_f := 6;
        ELSIF x =- 11942 THEN
            sigmoid_f := 6;
        ELSIF x =- 11941 THEN
            sigmoid_f := 6;
        ELSIF x =- 11940 THEN
            sigmoid_f := 6;
        ELSIF x =- 11939 THEN
            sigmoid_f := 6;
        ELSIF x =- 11938 THEN
            sigmoid_f := 6;
        ELSIF x =- 11937 THEN
            sigmoid_f := 6;
        ELSIF x =- 11936 THEN
            sigmoid_f := 6;
        ELSIF x =- 11935 THEN
            sigmoid_f := 6;
        ELSIF x =- 11934 THEN
            sigmoid_f := 6;
        ELSIF x =- 11933 THEN
            sigmoid_f := 6;
        ELSIF x =- 11932 THEN
            sigmoid_f := 6;
        ELSIF x =- 11931 THEN
            sigmoid_f := 6;
        ELSIF x =- 11930 THEN
            sigmoid_f := 6;
        ELSIF x =- 11929 THEN
            sigmoid_f := 6;
        ELSIF x =- 11928 THEN
            sigmoid_f := 6;
        ELSIF x =- 11927 THEN
            sigmoid_f := 6;
        ELSIF x =- 11926 THEN
            sigmoid_f := 6;
        ELSIF x =- 11925 THEN
            sigmoid_f := 6;
        ELSIF x =- 11924 THEN
            sigmoid_f := 6;
        ELSIF x =- 11923 THEN
            sigmoid_f := 6;
        ELSIF x =- 11922 THEN
            sigmoid_f := 6;
        ELSIF x =- 11921 THEN
            sigmoid_f := 6;
        ELSIF x =- 11920 THEN
            sigmoid_f := 6;
        ELSIF x =- 11919 THEN
            sigmoid_f := 6;
        ELSIF x =- 11918 THEN
            sigmoid_f := 6;
        ELSIF x =- 11917 THEN
            sigmoid_f := 6;
        ELSIF x =- 11916 THEN
            sigmoid_f := 6;
        ELSIF x =- 11915 THEN
            sigmoid_f := 6;
        ELSIF x =- 11914 THEN
            sigmoid_f := 6;
        ELSIF x =- 11913 THEN
            sigmoid_f := 6;
        ELSIF x =- 11912 THEN
            sigmoid_f := 6;
        ELSIF x =- 11911 THEN
            sigmoid_f := 6;
        ELSIF x =- 11910 THEN
            sigmoid_f := 6;
        ELSIF x =- 11909 THEN
            sigmoid_f := 6;
        ELSIF x =- 11908 THEN
            sigmoid_f := 6;
        ELSIF x =- 11907 THEN
            sigmoid_f := 6;
        ELSIF x =- 11906 THEN
            sigmoid_f := 6;
        ELSIF x =- 11905 THEN
            sigmoid_f := 6;
        ELSIF x =- 11904 THEN
            sigmoid_f := 6;
        ELSIF x =- 11903 THEN
            sigmoid_f := 6;
        ELSIF x =- 11902 THEN
            sigmoid_f := 6;
        ELSIF x =- 11901 THEN
            sigmoid_f := 6;
        ELSIF x =- 11900 THEN
            sigmoid_f := 6;
        ELSIF x =- 11899 THEN
            sigmoid_f := 6;
        ELSIF x =- 11898 THEN
            sigmoid_f := 6;
        ELSIF x =- 11897 THEN
            sigmoid_f := 6;
        ELSIF x =- 11896 THEN
            sigmoid_f := 6;
        ELSIF x =- 11895 THEN
            sigmoid_f := 6;
        ELSIF x =- 11894 THEN
            sigmoid_f := 6;
        ELSIF x =- 11893 THEN
            sigmoid_f := 6;
        ELSIF x =- 11892 THEN
            sigmoid_f := 6;
        ELSIF x =- 11891 THEN
            sigmoid_f := 6;
        ELSIF x =- 11890 THEN
            sigmoid_f := 6;
        ELSIF x =- 11889 THEN
            sigmoid_f := 6;
        ELSIF x =- 11888 THEN
            sigmoid_f := 6;
        ELSIF x =- 11887 THEN
            sigmoid_f := 6;
        ELSIF x =- 11886 THEN
            sigmoid_f := 6;
        ELSIF x =- 11885 THEN
            sigmoid_f := 6;
        ELSIF x =- 11884 THEN
            sigmoid_f := 6;
        ELSIF x =- 11883 THEN
            sigmoid_f := 6;
        ELSIF x =- 11882 THEN
            sigmoid_f := 6;
        ELSIF x =- 11881 THEN
            sigmoid_f := 6;
        ELSIF x =- 11880 THEN
            sigmoid_f := 6;
        ELSIF x =- 11879 THEN
            sigmoid_f := 6;
        ELSIF x =- 11878 THEN
            sigmoid_f := 6;
        ELSIF x =- 11877 THEN
            sigmoid_f := 6;
        ELSIF x =- 11876 THEN
            sigmoid_f := 6;
        ELSIF x =- 11875 THEN
            sigmoid_f := 6;
        ELSIF x =- 11874 THEN
            sigmoid_f := 6;
        ELSIF x =- 11873 THEN
            sigmoid_f := 6;
        ELSIF x =- 11872 THEN
            sigmoid_f := 6;
        ELSIF x =- 11871 THEN
            sigmoid_f := 6;
        ELSIF x =- 11870 THEN
            sigmoid_f := 6;
        ELSIF x =- 11869 THEN
            sigmoid_f := 6;
        ELSIF x =- 11868 THEN
            sigmoid_f := 6;
        ELSIF x =- 11867 THEN
            sigmoid_f := 6;
        ELSIF x =- 11866 THEN
            sigmoid_f := 6;
        ELSIF x =- 11865 THEN
            sigmoid_f := 6;
        ELSIF x =- 11864 THEN
            sigmoid_f := 6;
        ELSIF x =- 11863 THEN
            sigmoid_f := 6;
        ELSIF x =- 11862 THEN
            sigmoid_f := 6;
        ELSIF x =- 11861 THEN
            sigmoid_f := 6;
        ELSIF x =- 11860 THEN
            sigmoid_f := 6;
        ELSIF x =- 11859 THEN
            sigmoid_f := 6;
        ELSIF x =- 11858 THEN
            sigmoid_f := 6;
        ELSIF x =- 11857 THEN
            sigmoid_f := 6;
        ELSIF x =- 11856 THEN
            sigmoid_f := 6;
        ELSIF x =- 11855 THEN
            sigmoid_f := 6;
        ELSIF x =- 11854 THEN
            sigmoid_f := 6;
        ELSIF x =- 11853 THEN
            sigmoid_f := 6;
        ELSIF x =- 11852 THEN
            sigmoid_f := 6;
        ELSIF x =- 11851 THEN
            sigmoid_f := 6;
        ELSIF x =- 11850 THEN
            sigmoid_f := 6;
        ELSIF x =- 11849 THEN
            sigmoid_f := 6;
        ELSIF x =- 11848 THEN
            sigmoid_f := 6;
        ELSIF x =- 11847 THEN
            sigmoid_f := 6;
        ELSIF x =- 11846 THEN
            sigmoid_f := 6;
        ELSIF x =- 11845 THEN
            sigmoid_f := 6;
        ELSIF x =- 11844 THEN
            sigmoid_f := 6;
        ELSIF x =- 11843 THEN
            sigmoid_f := 6;
        ELSIF x =- 11842 THEN
            sigmoid_f := 6;
        ELSIF x =- 11841 THEN
            sigmoid_f := 6;
        ELSIF x =- 11840 THEN
            sigmoid_f := 6;
        ELSIF x =- 11839 THEN
            sigmoid_f := 6;
        ELSIF x =- 11838 THEN
            sigmoid_f := 6;
        ELSIF x =- 11837 THEN
            sigmoid_f := 6;
        ELSIF x =- 11836 THEN
            sigmoid_f := 6;
        ELSIF x =- 11835 THEN
            sigmoid_f := 6;
        ELSIF x =- 11834 THEN
            sigmoid_f := 6;
        ELSIF x =- 11833 THEN
            sigmoid_f := 6;
        ELSIF x =- 11832 THEN
            sigmoid_f := 6;
        ELSIF x =- 11831 THEN
            sigmoid_f := 6;
        ELSIF x =- 11830 THEN
            sigmoid_f := 6;
        ELSIF x =- 11829 THEN
            sigmoid_f := 6;
        ELSIF x =- 11828 THEN
            sigmoid_f := 6;
        ELSIF x =- 11827 THEN
            sigmoid_f := 6;
        ELSIF x =- 11826 THEN
            sigmoid_f := 6;
        ELSIF x =- 11825 THEN
            sigmoid_f := 6;
        ELSIF x =- 11824 THEN
            sigmoid_f := 6;
        ELSIF x =- 11823 THEN
            sigmoid_f := 6;
        ELSIF x =- 11822 THEN
            sigmoid_f := 6;
        ELSIF x =- 11821 THEN
            sigmoid_f := 6;
        ELSIF x =- 11820 THEN
            sigmoid_f := 6;
        ELSIF x =- 11819 THEN
            sigmoid_f := 6;
        ELSIF x =- 11818 THEN
            sigmoid_f := 6;
        ELSIF x =- 11817 THEN
            sigmoid_f := 6;
        ELSIF x =- 11816 THEN
            sigmoid_f := 6;
        ELSIF x =- 11815 THEN
            sigmoid_f := 6;
        ELSIF x =- 11814 THEN
            sigmoid_f := 6;
        ELSIF x =- 11813 THEN
            sigmoid_f := 6;
        ELSIF x =- 11812 THEN
            sigmoid_f := 6;
        ELSIF x =- 11811 THEN
            sigmoid_f := 6;
        ELSIF x =- 11810 THEN
            sigmoid_f := 6;
        ELSIF x =- 11809 THEN
            sigmoid_f := 6;
        ELSIF x =- 11808 THEN
            sigmoid_f := 6;
        ELSIF x =- 11807 THEN
            sigmoid_f := 6;
        ELSIF x =- 11806 THEN
            sigmoid_f := 6;
        ELSIF x =- 11805 THEN
            sigmoid_f := 6;
        ELSIF x =- 11804 THEN
            sigmoid_f := 6;
        ELSIF x =- 11803 THEN
            sigmoid_f := 6;
        ELSIF x =- 11802 THEN
            sigmoid_f := 6;
        ELSIF x =- 11801 THEN
            sigmoid_f := 6;
        ELSIF x =- 11800 THEN
            sigmoid_f := 6;
        ELSIF x =- 11799 THEN
            sigmoid_f := 6;
        ELSIF x =- 11798 THEN
            sigmoid_f := 6;
        ELSIF x =- 11797 THEN
            sigmoid_f := 6;
        ELSIF x =- 11796 THEN
            sigmoid_f := 6;
        ELSIF x =- 11795 THEN
            sigmoid_f := 6;
        ELSIF x =- 11794 THEN
            sigmoid_f := 6;
        ELSIF x =- 11793 THEN
            sigmoid_f := 6;
        ELSIF x =- 11792 THEN
            sigmoid_f := 6;
        ELSIF x =- 11791 THEN
            sigmoid_f := 6;
        ELSIF x =- 11790 THEN
            sigmoid_f := 6;
        ELSIF x =- 11789 THEN
            sigmoid_f := 6;
        ELSIF x =- 11788 THEN
            sigmoid_f := 6;
        ELSIF x =- 11787 THEN
            sigmoid_f := 6;
        ELSIF x =- 11786 THEN
            sigmoid_f := 6;
        ELSIF x =- 11785 THEN
            sigmoid_f := 6;
        ELSIF x =- 11784 THEN
            sigmoid_f := 6;
        ELSIF x =- 11783 THEN
            sigmoid_f := 6;
        ELSIF x =- 11782 THEN
            sigmoid_f := 6;
        ELSIF x =- 11781 THEN
            sigmoid_f := 6;
        ELSIF x =- 11780 THEN
            sigmoid_f := 6;
        ELSIF x =- 11779 THEN
            sigmoid_f := 6;
        ELSIF x =- 11778 THEN
            sigmoid_f := 6;
        ELSIF x =- 11777 THEN
            sigmoid_f := 6;
        ELSIF x =- 11776 THEN
            sigmoid_f := 6;
        ELSIF x =- 11775 THEN
            sigmoid_f := 6;
        ELSIF x =- 11774 THEN
            sigmoid_f := 6;
        ELSIF x =- 11773 THEN
            sigmoid_f := 6;
        ELSIF x =- 11772 THEN
            sigmoid_f := 6;
        ELSIF x =- 11771 THEN
            sigmoid_f := 6;
        ELSIF x =- 11770 THEN
            sigmoid_f := 6;
        ELSIF x =- 11769 THEN
            sigmoid_f := 6;
        ELSIF x =- 11768 THEN
            sigmoid_f := 6;
        ELSIF x =- 11767 THEN
            sigmoid_f := 6;
        ELSIF x =- 11766 THEN
            sigmoid_f := 6;
        ELSIF x =- 11765 THEN
            sigmoid_f := 6;
        ELSIF x =- 11764 THEN
            sigmoid_f := 6;
        ELSIF x =- 11763 THEN
            sigmoid_f := 6;
        ELSIF x =- 11762 THEN
            sigmoid_f := 6;
        ELSIF x =- 11761 THEN
            sigmoid_f := 6;
        ELSIF x =- 11760 THEN
            sigmoid_f := 6;
        ELSIF x =- 11759 THEN
            sigmoid_f := 6;
        ELSIF x =- 11758 THEN
            sigmoid_f := 6;
        ELSIF x =- 11757 THEN
            sigmoid_f := 6;
        ELSIF x =- 11756 THEN
            sigmoid_f := 6;
        ELSIF x =- 11755 THEN
            sigmoid_f := 6;
        ELSIF x =- 11754 THEN
            sigmoid_f := 6;
        ELSIF x =- 11753 THEN
            sigmoid_f := 6;
        ELSIF x =- 11752 THEN
            sigmoid_f := 6;
        ELSIF x =- 11751 THEN
            sigmoid_f := 6;
        ELSIF x =- 11750 THEN
            sigmoid_f := 6;
        ELSIF x =- 11749 THEN
            sigmoid_f := 6;
        ELSIF x =- 11748 THEN
            sigmoid_f := 6;
        ELSIF x =- 11747 THEN
            sigmoid_f := 6;
        ELSIF x =- 11746 THEN
            sigmoid_f := 6;
        ELSIF x =- 11745 THEN
            sigmoid_f := 6;
        ELSIF x =- 11744 THEN
            sigmoid_f := 6;
        ELSIF x =- 11743 THEN
            sigmoid_f := 6;
        ELSIF x =- 11742 THEN
            sigmoid_f := 6;
        ELSIF x =- 11741 THEN
            sigmoid_f := 6;
        ELSIF x =- 11740 THEN
            sigmoid_f := 6;
        ELSIF x =- 11739 THEN
            sigmoid_f := 6;
        ELSIF x =- 11738 THEN
            sigmoid_f := 6;
        ELSIF x =- 11737 THEN
            sigmoid_f := 6;
        ELSIF x =- 11736 THEN
            sigmoid_f := 6;
        ELSIF x =- 11735 THEN
            sigmoid_f := 6;
        ELSIF x =- 11734 THEN
            sigmoid_f := 6;
        ELSIF x =- 11733 THEN
            sigmoid_f := 6;
        ELSIF x =- 11732 THEN
            sigmoid_f := 6;
        ELSIF x =- 11731 THEN
            sigmoid_f := 6;
        ELSIF x =- 11730 THEN
            sigmoid_f := 6;
        ELSIF x =- 11729 THEN
            sigmoid_f := 6;
        ELSIF x =- 11728 THEN
            sigmoid_f := 6;
        ELSIF x =- 11727 THEN
            sigmoid_f := 6;
        ELSIF x =- 11726 THEN
            sigmoid_f := 6;
        ELSIF x =- 11725 THEN
            sigmoid_f := 6;
        ELSIF x =- 11724 THEN
            sigmoid_f := 6;
        ELSIF x =- 11723 THEN
            sigmoid_f := 6;
        ELSIF x =- 11722 THEN
            sigmoid_f := 6;
        ELSIF x =- 11721 THEN
            sigmoid_f := 6;
        ELSIF x =- 11720 THEN
            sigmoid_f := 6;
        ELSIF x =- 11719 THEN
            sigmoid_f := 6;
        ELSIF x =- 11718 THEN
            sigmoid_f := 6;
        ELSIF x =- 11717 THEN
            sigmoid_f := 6;
        ELSIF x =- 11716 THEN
            sigmoid_f := 6;
        ELSIF x =- 11715 THEN
            sigmoid_f := 6;
        ELSIF x =- 11714 THEN
            sigmoid_f := 6;
        ELSIF x =- 11713 THEN
            sigmoid_f := 6;
        ELSIF x =- 11712 THEN
            sigmoid_f := 6;
        ELSIF x =- 11711 THEN
            sigmoid_f := 6;
        ELSIF x =- 11710 THEN
            sigmoid_f := 6;
        ELSIF x =- 11709 THEN
            sigmoid_f := 6;
        ELSIF x =- 11708 THEN
            sigmoid_f := 6;
        ELSIF x =- 11707 THEN
            sigmoid_f := 6;
        ELSIF x =- 11706 THEN
            sigmoid_f := 6;
        ELSIF x =- 11705 THEN
            sigmoid_f := 6;
        ELSIF x =- 11704 THEN
            sigmoid_f := 6;
        ELSIF x =- 11703 THEN
            sigmoid_f := 6;
        ELSIF x =- 11702 THEN
            sigmoid_f := 6;
        ELSIF x =- 11701 THEN
            sigmoid_f := 6;
        ELSIF x =- 11700 THEN
            sigmoid_f := 6;
        ELSIF x =- 11699 THEN
            sigmoid_f := 6;
        ELSIF x =- 11698 THEN
            sigmoid_f := 6;
        ELSIF x =- 11697 THEN
            sigmoid_f := 6;
        ELSIF x =- 11696 THEN
            sigmoid_f := 6;
        ELSIF x =- 11695 THEN
            sigmoid_f := 6;
        ELSIF x =- 11694 THEN
            sigmoid_f := 6;
        ELSIF x =- 11693 THEN
            sigmoid_f := 6;
        ELSIF x =- 11692 THEN
            sigmoid_f := 6;
        ELSIF x =- 11691 THEN
            sigmoid_f := 6;
        ELSIF x =- 11690 THEN
            sigmoid_f := 6;
        ELSIF x =- 11689 THEN
            sigmoid_f := 6;
        ELSIF x =- 11688 THEN
            sigmoid_f := 6;
        ELSIF x =- 11687 THEN
            sigmoid_f := 6;
        ELSIF x =- 11686 THEN
            sigmoid_f := 6;
        ELSIF x =- 11685 THEN
            sigmoid_f := 6;
        ELSIF x =- 11684 THEN
            sigmoid_f := 6;
        ELSIF x =- 11683 THEN
            sigmoid_f := 6;
        ELSIF x =- 11682 THEN
            sigmoid_f := 6;
        ELSIF x =- 11681 THEN
            sigmoid_f := 6;
        ELSIF x =- 11680 THEN
            sigmoid_f := 6;
        ELSIF x =- 11679 THEN
            sigmoid_f := 6;
        ELSIF x =- 11678 THEN
            sigmoid_f := 6;
        ELSIF x =- 11677 THEN
            sigmoid_f := 6;
        ELSIF x =- 11676 THEN
            sigmoid_f := 6;
        ELSIF x =- 11675 THEN
            sigmoid_f := 6;
        ELSIF x =- 11674 THEN
            sigmoid_f := 6;
        ELSIF x =- 11673 THEN
            sigmoid_f := 6;
        ELSIF x =- 11672 THEN
            sigmoid_f := 6;
        ELSIF x =- 11671 THEN
            sigmoid_f := 6;
        ELSIF x =- 11670 THEN
            sigmoid_f := 6;
        ELSIF x =- 11669 THEN
            sigmoid_f := 6;
        ELSIF x =- 11668 THEN
            sigmoid_f := 6;
        ELSIF x =- 11667 THEN
            sigmoid_f := 6;
        ELSIF x =- 11666 THEN
            sigmoid_f := 6;
        ELSIF x =- 11665 THEN
            sigmoid_f := 6;
        ELSIF x =- 11664 THEN
            sigmoid_f := 6;
        ELSIF x =- 11663 THEN
            sigmoid_f := 6;
        ELSIF x =- 11662 THEN
            sigmoid_f := 6;
        ELSIF x =- 11661 THEN
            sigmoid_f := 6;
        ELSIF x =- 11660 THEN
            sigmoid_f := 6;
        ELSIF x =- 11659 THEN
            sigmoid_f := 6;
        ELSIF x =- 11658 THEN
            sigmoid_f := 6;
        ELSIF x =- 11657 THEN
            sigmoid_f := 6;
        ELSIF x =- 11656 THEN
            sigmoid_f := 6;
        ELSIF x =- 11655 THEN
            sigmoid_f := 6;
        ELSIF x =- 11654 THEN
            sigmoid_f := 6;
        ELSIF x =- 11653 THEN
            sigmoid_f := 6;
        ELSIF x =- 11652 THEN
            sigmoid_f := 6;
        ELSIF x =- 11651 THEN
            sigmoid_f := 6;
        ELSIF x =- 11650 THEN
            sigmoid_f := 6;
        ELSIF x =- 11649 THEN
            sigmoid_f := 6;
        ELSIF x =- 11648 THEN
            sigmoid_f := 6;
        ELSIF x =- 11647 THEN
            sigmoid_f := 6;
        ELSIF x =- 11646 THEN
            sigmoid_f := 6;
        ELSIF x =- 11645 THEN
            sigmoid_f := 6;
        ELSIF x =- 11644 THEN
            sigmoid_f := 6;
        ELSIF x =- 11643 THEN
            sigmoid_f := 6;
        ELSIF x =- 11642 THEN
            sigmoid_f := 6;
        ELSIF x =- 11641 THEN
            sigmoid_f := 6;
        ELSIF x =- 11640 THEN
            sigmoid_f := 6;
        ELSIF x =- 11639 THEN
            sigmoid_f := 6;
        ELSIF x =- 11638 THEN
            sigmoid_f := 6;
        ELSIF x =- 11637 THEN
            sigmoid_f := 6;
        ELSIF x =- 11636 THEN
            sigmoid_f := 6;
        ELSIF x =- 11635 THEN
            sigmoid_f := 6;
        ELSIF x =- 11634 THEN
            sigmoid_f := 6;
        ELSIF x =- 11633 THEN
            sigmoid_f := 6;
        ELSIF x =- 11632 THEN
            sigmoid_f := 6;
        ELSIF x =- 11631 THEN
            sigmoid_f := 6;
        ELSIF x =- 11630 THEN
            sigmoid_f := 6;
        ELSIF x =- 11629 THEN
            sigmoid_f := 6;
        ELSIF x =- 11628 THEN
            sigmoid_f := 6;
        ELSIF x =- 11627 THEN
            sigmoid_f := 6;
        ELSIF x =- 11626 THEN
            sigmoid_f := 6;
        ELSIF x =- 11625 THEN
            sigmoid_f := 6;
        ELSIF x =- 11624 THEN
            sigmoid_f := 6;
        ELSIF x =- 11623 THEN
            sigmoid_f := 6;
        ELSIF x =- 11622 THEN
            sigmoid_f := 6;
        ELSIF x =- 11621 THEN
            sigmoid_f := 6;
        ELSIF x =- 11620 THEN
            sigmoid_f := 6;
        ELSIF x =- 11619 THEN
            sigmoid_f := 6;
        ELSIF x =- 11618 THEN
            sigmoid_f := 6;
        ELSIF x =- 11617 THEN
            sigmoid_f := 6;
        ELSIF x =- 11616 THEN
            sigmoid_f := 6;
        ELSIF x =- 11615 THEN
            sigmoid_f := 6;
        ELSIF x =- 11614 THEN
            sigmoid_f := 6;
        ELSIF x =- 11613 THEN
            sigmoid_f := 6;
        ELSIF x =- 11612 THEN
            sigmoid_f := 6;
        ELSIF x =- 11611 THEN
            sigmoid_f := 6;
        ELSIF x =- 11610 THEN
            sigmoid_f := 6;
        ELSIF x =- 11609 THEN
            sigmoid_f := 6;
        ELSIF x =- 11608 THEN
            sigmoid_f := 6;
        ELSIF x =- 11607 THEN
            sigmoid_f := 6;
        ELSIF x =- 11606 THEN
            sigmoid_f := 6;
        ELSIF x =- 11605 THEN
            sigmoid_f := 7;
        ELSIF x =- 11604 THEN
            sigmoid_f := 7;
        ELSIF x =- 11603 THEN
            sigmoid_f := 7;
        ELSIF x =- 11602 THEN
            sigmoid_f := 7;
        ELSIF x =- 11601 THEN
            sigmoid_f := 7;
        ELSIF x =- 11600 THEN
            sigmoid_f := 7;
        ELSIF x =- 11599 THEN
            sigmoid_f := 7;
        ELSIF x =- 11598 THEN
            sigmoid_f := 7;
        ELSIF x =- 11597 THEN
            sigmoid_f := 7;
        ELSIF x =- 11596 THEN
            sigmoid_f := 7;
        ELSIF x =- 11595 THEN
            sigmoid_f := 7;
        ELSIF x =- 11594 THEN
            sigmoid_f := 7;
        ELSIF x =- 11593 THEN
            sigmoid_f := 7;
        ELSIF x =- 11592 THEN
            sigmoid_f := 7;
        ELSIF x =- 11591 THEN
            sigmoid_f := 7;
        ELSIF x =- 11590 THEN
            sigmoid_f := 7;
        ELSIF x =- 11589 THEN
            sigmoid_f := 7;
        ELSIF x =- 11588 THEN
            sigmoid_f := 7;
        ELSIF x =- 11587 THEN
            sigmoid_f := 7;
        ELSIF x =- 11586 THEN
            sigmoid_f := 7;
        ELSIF x =- 11585 THEN
            sigmoid_f := 7;
        ELSIF x =- 11584 THEN
            sigmoid_f := 7;
        ELSIF x =- 11583 THEN
            sigmoid_f := 7;
        ELSIF x =- 11582 THEN
            sigmoid_f := 7;
        ELSIF x =- 11581 THEN
            sigmoid_f := 7;
        ELSIF x =- 11580 THEN
            sigmoid_f := 7;
        ELSIF x =- 11579 THEN
            sigmoid_f := 7;
        ELSIF x =- 11578 THEN
            sigmoid_f := 7;
        ELSIF x =- 11577 THEN
            sigmoid_f := 7;
        ELSIF x =- 11576 THEN
            sigmoid_f := 7;
        ELSIF x =- 11575 THEN
            sigmoid_f := 7;
        ELSIF x =- 11574 THEN
            sigmoid_f := 7;
        ELSIF x =- 11573 THEN
            sigmoid_f := 7;
        ELSIF x =- 11572 THEN
            sigmoid_f := 7;
        ELSIF x =- 11571 THEN
            sigmoid_f := 7;
        ELSIF x =- 11570 THEN
            sigmoid_f := 7;
        ELSIF x =- 11569 THEN
            sigmoid_f := 7;
        ELSIF x =- 11568 THEN
            sigmoid_f := 7;
        ELSIF x =- 11567 THEN
            sigmoid_f := 7;
        ELSIF x =- 11566 THEN
            sigmoid_f := 7;
        ELSIF x =- 11565 THEN
            sigmoid_f := 7;
        ELSIF x =- 11564 THEN
            sigmoid_f := 7;
        ELSIF x =- 11563 THEN
            sigmoid_f := 7;
        ELSIF x =- 11562 THEN
            sigmoid_f := 7;
        ELSIF x =- 11561 THEN
            sigmoid_f := 7;
        ELSIF x =- 11560 THEN
            sigmoid_f := 7;
        ELSIF x =- 11559 THEN
            sigmoid_f := 7;
        ELSIF x =- 11558 THEN
            sigmoid_f := 7;
        ELSIF x =- 11557 THEN
            sigmoid_f := 7;
        ELSIF x =- 11556 THEN
            sigmoid_f := 7;
        ELSIF x =- 11555 THEN
            sigmoid_f := 7;
        ELSIF x =- 11554 THEN
            sigmoid_f := 7;
        ELSIF x =- 11553 THEN
            sigmoid_f := 7;
        ELSIF x =- 11552 THEN
            sigmoid_f := 7;
        ELSIF x =- 11551 THEN
            sigmoid_f := 7;
        ELSIF x =- 11550 THEN
            sigmoid_f := 7;
        ELSIF x =- 11549 THEN
            sigmoid_f := 7;
        ELSIF x =- 11548 THEN
            sigmoid_f := 7;
        ELSIF x =- 11547 THEN
            sigmoid_f := 7;
        ELSIF x =- 11546 THEN
            sigmoid_f := 7;
        ELSIF x =- 11545 THEN
            sigmoid_f := 7;
        ELSIF x =- 11544 THEN
            sigmoid_f := 7;
        ELSIF x =- 11543 THEN
            sigmoid_f := 7;
        ELSIF x =- 11542 THEN
            sigmoid_f := 7;
        ELSIF x =- 11541 THEN
            sigmoid_f := 7;
        ELSIF x =- 11540 THEN
            sigmoid_f := 7;
        ELSIF x =- 11539 THEN
            sigmoid_f := 7;
        ELSIF x =- 11538 THEN
            sigmoid_f := 7;
        ELSIF x =- 11537 THEN
            sigmoid_f := 7;
        ELSIF x =- 11536 THEN
            sigmoid_f := 7;
        ELSIF x =- 11535 THEN
            sigmoid_f := 7;
        ELSIF x =- 11534 THEN
            sigmoid_f := 7;
        ELSIF x =- 11533 THEN
            sigmoid_f := 7;
        ELSIF x =- 11532 THEN
            sigmoid_f := 7;
        ELSIF x =- 11531 THEN
            sigmoid_f := 7;
        ELSIF x =- 11530 THEN
            sigmoid_f := 7;
        ELSIF x =- 11529 THEN
            sigmoid_f := 7;
        ELSIF x =- 11528 THEN
            sigmoid_f := 7;
        ELSIF x =- 11527 THEN
            sigmoid_f := 7;
        ELSIF x =- 11526 THEN
            sigmoid_f := 7;
        ELSIF x =- 11525 THEN
            sigmoid_f := 7;
        ELSIF x =- 11524 THEN
            sigmoid_f := 7;
        ELSIF x =- 11523 THEN
            sigmoid_f := 7;
        ELSIF x =- 11522 THEN
            sigmoid_f := 7;
        ELSIF x =- 11521 THEN
            sigmoid_f := 7;
        ELSIF x =- 11520 THEN
            sigmoid_f := 7;
        ELSIF x =- 11519 THEN
            sigmoid_f := 7;
        ELSIF x =- 11518 THEN
            sigmoid_f := 7;
        ELSIF x =- 11517 THEN
            sigmoid_f := 7;
        ELSIF x =- 11516 THEN
            sigmoid_f := 7;
        ELSIF x =- 11515 THEN
            sigmoid_f := 7;
        ELSIF x =- 11514 THEN
            sigmoid_f := 7;
        ELSIF x =- 11513 THEN
            sigmoid_f := 7;
        ELSIF x =- 11512 THEN
            sigmoid_f := 7;
        ELSIF x =- 11511 THEN
            sigmoid_f := 7;
        ELSIF x =- 11510 THEN
            sigmoid_f := 7;
        ELSIF x =- 11509 THEN
            sigmoid_f := 7;
        ELSIF x =- 11508 THEN
            sigmoid_f := 7;
        ELSIF x =- 11507 THEN
            sigmoid_f := 7;
        ELSIF x =- 11506 THEN
            sigmoid_f := 7;
        ELSIF x =- 11505 THEN
            sigmoid_f := 7;
        ELSIF x =- 11504 THEN
            sigmoid_f := 7;
        ELSIF x =- 11503 THEN
            sigmoid_f := 7;
        ELSIF x =- 11502 THEN
            sigmoid_f := 7;
        ELSIF x =- 11501 THEN
            sigmoid_f := 7;
        ELSIF x =- 11500 THEN
            sigmoid_f := 7;
        ELSIF x =- 11499 THEN
            sigmoid_f := 7;
        ELSIF x =- 11498 THEN
            sigmoid_f := 7;
        ELSIF x =- 11497 THEN
            sigmoid_f := 7;
        ELSIF x =- 11496 THEN
            sigmoid_f := 7;
        ELSIF x =- 11495 THEN
            sigmoid_f := 7;
        ELSIF x =- 11494 THEN
            sigmoid_f := 7;
        ELSIF x =- 11493 THEN
            sigmoid_f := 7;
        ELSIF x =- 11492 THEN
            sigmoid_f := 7;
        ELSIF x =- 11491 THEN
            sigmoid_f := 7;
        ELSIF x =- 11490 THEN
            sigmoid_f := 7;
        ELSIF x =- 11489 THEN
            sigmoid_f := 7;
        ELSIF x =- 11488 THEN
            sigmoid_f := 7;
        ELSIF x =- 11487 THEN
            sigmoid_f := 7;
        ELSIF x =- 11486 THEN
            sigmoid_f := 7;
        ELSIF x =- 11485 THEN
            sigmoid_f := 7;
        ELSIF x =- 11484 THEN
            sigmoid_f := 7;
        ELSIF x =- 11483 THEN
            sigmoid_f := 7;
        ELSIF x =- 11482 THEN
            sigmoid_f := 7;
        ELSIF x =- 11481 THEN
            sigmoid_f := 7;
        ELSIF x =- 11480 THEN
            sigmoid_f := 7;
        ELSIF x =- 11479 THEN
            sigmoid_f := 7;
        ELSIF x =- 11478 THEN
            sigmoid_f := 7;
        ELSIF x =- 11477 THEN
            sigmoid_f := 7;
        ELSIF x =- 11476 THEN
            sigmoid_f := 7;
        ELSIF x =- 11475 THEN
            sigmoid_f := 7;
        ELSIF x =- 11474 THEN
            sigmoid_f := 7;
        ELSIF x =- 11473 THEN
            sigmoid_f := 7;
        ELSIF x =- 11472 THEN
            sigmoid_f := 7;
        ELSIF x =- 11471 THEN
            sigmoid_f := 7;
        ELSIF x =- 11470 THEN
            sigmoid_f := 7;
        ELSIF x =- 11469 THEN
            sigmoid_f := 7;
        ELSIF x =- 11468 THEN
            sigmoid_f := 7;
        ELSIF x =- 11467 THEN
            sigmoid_f := 7;
        ELSIF x =- 11466 THEN
            sigmoid_f := 7;
        ELSIF x =- 11465 THEN
            sigmoid_f := 7;
        ELSIF x =- 11464 THEN
            sigmoid_f := 7;
        ELSIF x =- 11463 THEN
            sigmoid_f := 7;
        ELSIF x =- 11462 THEN
            sigmoid_f := 7;
        ELSIF x =- 11461 THEN
            sigmoid_f := 7;
        ELSIF x =- 11460 THEN
            sigmoid_f := 7;
        ELSIF x =- 11459 THEN
            sigmoid_f := 7;
        ELSIF x =- 11458 THEN
            sigmoid_f := 7;
        ELSIF x =- 11457 THEN
            sigmoid_f := 7;
        ELSIF x =- 11456 THEN
            sigmoid_f := 7;
        ELSIF x =- 11455 THEN
            sigmoid_f := 7;
        ELSIF x =- 11454 THEN
            sigmoid_f := 7;
        ELSIF x =- 11453 THEN
            sigmoid_f := 7;
        ELSIF x =- 11452 THEN
            sigmoid_f := 7;
        ELSIF x =- 11451 THEN
            sigmoid_f := 7;
        ELSIF x =- 11450 THEN
            sigmoid_f := 7;
        ELSIF x =- 11449 THEN
            sigmoid_f := 7;
        ELSIF x =- 11448 THEN
            sigmoid_f := 7;
        ELSIF x =- 11447 THEN
            sigmoid_f := 7;
        ELSIF x =- 11446 THEN
            sigmoid_f := 7;
        ELSIF x =- 11445 THEN
            sigmoid_f := 7;
        ELSIF x =- 11444 THEN
            sigmoid_f := 7;
        ELSIF x =- 11443 THEN
            sigmoid_f := 7;
        ELSIF x =- 11442 THEN
            sigmoid_f := 7;
        ELSIF x =- 11441 THEN
            sigmoid_f := 7;
        ELSIF x =- 11440 THEN
            sigmoid_f := 7;
        ELSIF x =- 11439 THEN
            sigmoid_f := 7;
        ELSIF x =- 11438 THEN
            sigmoid_f := 7;
        ELSIF x =- 11437 THEN
            sigmoid_f := 7;
        ELSIF x =- 11436 THEN
            sigmoid_f := 7;
        ELSIF x =- 11435 THEN
            sigmoid_f := 7;
        ELSIF x =- 11434 THEN
            sigmoid_f := 7;
        ELSIF x =- 11433 THEN
            sigmoid_f := 7;
        ELSIF x =- 11432 THEN
            sigmoid_f := 7;
        ELSIF x =- 11431 THEN
            sigmoid_f := 7;
        ELSIF x =- 11430 THEN
            sigmoid_f := 7;
        ELSIF x =- 11429 THEN
            sigmoid_f := 7;
        ELSIF x =- 11428 THEN
            sigmoid_f := 7;
        ELSIF x =- 11427 THEN
            sigmoid_f := 7;
        ELSIF x =- 11426 THEN
            sigmoid_f := 7;
        ELSIF x =- 11425 THEN
            sigmoid_f := 7;
        ELSIF x =- 11424 THEN
            sigmoid_f := 7;
        ELSIF x =- 11423 THEN
            sigmoid_f := 7;
        ELSIF x =- 11422 THEN
            sigmoid_f := 7;
        ELSIF x =- 11421 THEN
            sigmoid_f := 7;
        ELSIF x =- 11420 THEN
            sigmoid_f := 7;
        ELSIF x =- 11419 THEN
            sigmoid_f := 7;
        ELSIF x =- 11418 THEN
            sigmoid_f := 7;
        ELSIF x =- 11417 THEN
            sigmoid_f := 7;
        ELSIF x =- 11416 THEN
            sigmoid_f := 7;
        ELSIF x =- 11415 THEN
            sigmoid_f := 7;
        ELSIF x =- 11414 THEN
            sigmoid_f := 7;
        ELSIF x =- 11413 THEN
            sigmoid_f := 7;
        ELSIF x =- 11412 THEN
            sigmoid_f := 7;
        ELSIF x =- 11411 THEN
            sigmoid_f := 7;
        ELSIF x =- 11410 THEN
            sigmoid_f := 7;
        ELSIF x =- 11409 THEN
            sigmoid_f := 7;
        ELSIF x =- 11408 THEN
            sigmoid_f := 7;
        ELSIF x =- 11407 THEN
            sigmoid_f := 7;
        ELSIF x =- 11406 THEN
            sigmoid_f := 7;
        ELSIF x =- 11405 THEN
            sigmoid_f := 7;
        ELSIF x =- 11404 THEN
            sigmoid_f := 7;
        ELSIF x =- 11403 THEN
            sigmoid_f := 7;
        ELSIF x =- 11402 THEN
            sigmoid_f := 7;
        ELSIF x =- 11401 THEN
            sigmoid_f := 7;
        ELSIF x =- 11400 THEN
            sigmoid_f := 7;
        ELSIF x =- 11399 THEN
            sigmoid_f := 7;
        ELSIF x =- 11398 THEN
            sigmoid_f := 7;
        ELSIF x =- 11397 THEN
            sigmoid_f := 7;
        ELSIF x =- 11396 THEN
            sigmoid_f := 7;
        ELSIF x =- 11395 THEN
            sigmoid_f := 7;
        ELSIF x =- 11394 THEN
            sigmoid_f := 7;
        ELSIF x =- 11393 THEN
            sigmoid_f := 7;
        ELSIF x =- 11392 THEN
            sigmoid_f := 7;
        ELSIF x =- 11391 THEN
            sigmoid_f := 7;
        ELSIF x =- 11390 THEN
            sigmoid_f := 7;
        ELSIF x =- 11389 THEN
            sigmoid_f := 7;
        ELSIF x =- 11388 THEN
            sigmoid_f := 7;
        ELSIF x =- 11387 THEN
            sigmoid_f := 7;
        ELSIF x =- 11386 THEN
            sigmoid_f := 7;
        ELSIF x =- 11385 THEN
            sigmoid_f := 7;
        ELSIF x =- 11384 THEN
            sigmoid_f := 7;
        ELSIF x =- 11383 THEN
            sigmoid_f := 7;
        ELSIF x =- 11382 THEN
            sigmoid_f := 7;
        ELSIF x =- 11381 THEN
            sigmoid_f := 7;
        ELSIF x =- 11380 THEN
            sigmoid_f := 7;
        ELSIF x =- 11379 THEN
            sigmoid_f := 7;
        ELSIF x =- 11378 THEN
            sigmoid_f := 7;
        ELSIF x =- 11377 THEN
            sigmoid_f := 8;
        ELSIF x =- 11376 THEN
            sigmoid_f := 8;
        ELSIF x =- 11375 THEN
            sigmoid_f := 8;
        ELSIF x =- 11374 THEN
            sigmoid_f := 8;
        ELSIF x =- 11373 THEN
            sigmoid_f := 8;
        ELSIF x =- 11372 THEN
            sigmoid_f := 8;
        ELSIF x =- 11371 THEN
            sigmoid_f := 8;
        ELSIF x =- 11370 THEN
            sigmoid_f := 8;
        ELSIF x =- 11369 THEN
            sigmoid_f := 8;
        ELSIF x =- 11368 THEN
            sigmoid_f := 8;
        ELSIF x =- 11367 THEN
            sigmoid_f := 8;
        ELSIF x =- 11366 THEN
            sigmoid_f := 8;
        ELSIF x =- 11365 THEN
            sigmoid_f := 8;
        ELSIF x =- 11364 THEN
            sigmoid_f := 8;
        ELSIF x =- 11363 THEN
            sigmoid_f := 8;
        ELSIF x =- 11362 THEN
            sigmoid_f := 8;
        ELSIF x =- 11361 THEN
            sigmoid_f := 8;
        ELSIF x =- 11360 THEN
            sigmoid_f := 8;
        ELSIF x =- 11359 THEN
            sigmoid_f := 8;
        ELSIF x =- 11358 THEN
            sigmoid_f := 8;
        ELSIF x =- 11357 THEN
            sigmoid_f := 8;
        ELSIF x =- 11356 THEN
            sigmoid_f := 8;
        ELSIF x =- 11355 THEN
            sigmoid_f := 8;
        ELSIF x =- 11354 THEN
            sigmoid_f := 8;
        ELSIF x =- 11353 THEN
            sigmoid_f := 8;
        ELSIF x =- 11352 THEN
            sigmoid_f := 8;
        ELSIF x =- 11351 THEN
            sigmoid_f := 8;
        ELSIF x =- 11350 THEN
            sigmoid_f := 8;
        ELSIF x =- 11349 THEN
            sigmoid_f := 8;
        ELSIF x =- 11348 THEN
            sigmoid_f := 8;
        ELSIF x =- 11347 THEN
            sigmoid_f := 8;
        ELSIF x =- 11346 THEN
            sigmoid_f := 8;
        ELSIF x =- 11345 THEN
            sigmoid_f := 8;
        ELSIF x =- 11344 THEN
            sigmoid_f := 8;
        ELSIF x =- 11343 THEN
            sigmoid_f := 8;
        ELSIF x =- 11342 THEN
            sigmoid_f := 8;
        ELSIF x =- 11341 THEN
            sigmoid_f := 8;
        ELSIF x =- 11340 THEN
            sigmoid_f := 8;
        ELSIF x =- 11339 THEN
            sigmoid_f := 8;
        ELSIF x =- 11338 THEN
            sigmoid_f := 8;
        ELSIF x =- 11337 THEN
            sigmoid_f := 8;
        ELSIF x =- 11336 THEN
            sigmoid_f := 8;
        ELSIF x =- 11335 THEN
            sigmoid_f := 8;
        ELSIF x =- 11334 THEN
            sigmoid_f := 8;
        ELSIF x =- 11333 THEN
            sigmoid_f := 8;
        ELSIF x =- 11332 THEN
            sigmoid_f := 8;
        ELSIF x =- 11331 THEN
            sigmoid_f := 8;
        ELSIF x =- 11330 THEN
            sigmoid_f := 8;
        ELSIF x =- 11329 THEN
            sigmoid_f := 8;
        ELSIF x =- 11328 THEN
            sigmoid_f := 8;
        ELSIF x =- 11327 THEN
            sigmoid_f := 8;
        ELSIF x =- 11326 THEN
            sigmoid_f := 8;
        ELSIF x =- 11325 THEN
            sigmoid_f := 8;
        ELSIF x =- 11324 THEN
            sigmoid_f := 8;
        ELSIF x =- 11323 THEN
            sigmoid_f := 8;
        ELSIF x =- 11322 THEN
            sigmoid_f := 8;
        ELSIF x =- 11321 THEN
            sigmoid_f := 8;
        ELSIF x =- 11320 THEN
            sigmoid_f := 8;
        ELSIF x =- 11319 THEN
            sigmoid_f := 8;
        ELSIF x =- 11318 THEN
            sigmoid_f := 8;
        ELSIF x =- 11317 THEN
            sigmoid_f := 8;
        ELSIF x =- 11316 THEN
            sigmoid_f := 8;
        ELSIF x =- 11315 THEN
            sigmoid_f := 8;
        ELSIF x =- 11314 THEN
            sigmoid_f := 8;
        ELSIF x =- 11313 THEN
            sigmoid_f := 8;
        ELSIF x =- 11312 THEN
            sigmoid_f := 8;
        ELSIF x =- 11311 THEN
            sigmoid_f := 8;
        ELSIF x =- 11310 THEN
            sigmoid_f := 8;
        ELSIF x =- 11309 THEN
            sigmoid_f := 8;
        ELSIF x =- 11308 THEN
            sigmoid_f := 8;
        ELSIF x =- 11307 THEN
            sigmoid_f := 8;
        ELSIF x =- 11306 THEN
            sigmoid_f := 8;
        ELSIF x =- 11305 THEN
            sigmoid_f := 8;
        ELSIF x =- 11304 THEN
            sigmoid_f := 8;
        ELSIF x =- 11303 THEN
            sigmoid_f := 8;
        ELSIF x =- 11302 THEN
            sigmoid_f := 8;
        ELSIF x =- 11301 THEN
            sigmoid_f := 8;
        ELSIF x =- 11300 THEN
            sigmoid_f := 8;
        ELSIF x =- 11299 THEN
            sigmoid_f := 8;
        ELSIF x =- 11298 THEN
            sigmoid_f := 8;
        ELSIF x =- 11297 THEN
            sigmoid_f := 8;
        ELSIF x =- 11296 THEN
            sigmoid_f := 8;
        ELSIF x =- 11295 THEN
            sigmoid_f := 8;
        ELSIF x =- 11294 THEN
            sigmoid_f := 8;
        ELSIF x =- 11293 THEN
            sigmoid_f := 8;
        ELSIF x =- 11292 THEN
            sigmoid_f := 8;
        ELSIF x =- 11291 THEN
            sigmoid_f := 8;
        ELSIF x =- 11290 THEN
            sigmoid_f := 8;
        ELSIF x =- 11289 THEN
            sigmoid_f := 8;
        ELSIF x =- 11288 THEN
            sigmoid_f := 8;
        ELSIF x =- 11287 THEN
            sigmoid_f := 8;
        ELSIF x =- 11286 THEN
            sigmoid_f := 8;
        ELSIF x =- 11285 THEN
            sigmoid_f := 8;
        ELSIF x =- 11284 THEN
            sigmoid_f := 8;
        ELSIF x =- 11283 THEN
            sigmoid_f := 8;
        ELSIF x =- 11282 THEN
            sigmoid_f := 8;
        ELSIF x =- 11281 THEN
            sigmoid_f := 8;
        ELSIF x =- 11280 THEN
            sigmoid_f := 8;
        ELSIF x =- 11279 THEN
            sigmoid_f := 8;
        ELSIF x =- 11278 THEN
            sigmoid_f := 8;
        ELSIF x =- 11277 THEN
            sigmoid_f := 8;
        ELSIF x =- 11276 THEN
            sigmoid_f := 8;
        ELSIF x =- 11275 THEN
            sigmoid_f := 8;
        ELSIF x =- 11274 THEN
            sigmoid_f := 8;
        ELSIF x =- 11273 THEN
            sigmoid_f := 8;
        ELSIF x =- 11272 THEN
            sigmoid_f := 8;
        ELSIF x =- 11271 THEN
            sigmoid_f := 8;
        ELSIF x =- 11270 THEN
            sigmoid_f := 8;
        ELSIF x =- 11269 THEN
            sigmoid_f := 8;
        ELSIF x =- 11268 THEN
            sigmoid_f := 8;
        ELSIF x =- 11267 THEN
            sigmoid_f := 8;
        ELSIF x =- 11266 THEN
            sigmoid_f := 8;
        ELSIF x =- 11265 THEN
            sigmoid_f := 8;
        ELSIF x =- 11264 THEN
            sigmoid_f := 8;
        ELSIF x =- 11263 THEN
            sigmoid_f := 8;
        ELSIF x =- 11262 THEN
            sigmoid_f := 8;
        ELSIF x =- 11261 THEN
            sigmoid_f := 8;
        ELSIF x =- 11260 THEN
            sigmoid_f := 8;
        ELSIF x =- 11259 THEN
            sigmoid_f := 8;
        ELSIF x =- 11258 THEN
            sigmoid_f := 8;
        ELSIF x =- 11257 THEN
            sigmoid_f := 8;
        ELSIF x =- 11256 THEN
            sigmoid_f := 8;
        ELSIF x =- 11255 THEN
            sigmoid_f := 8;
        ELSIF x =- 11254 THEN
            sigmoid_f := 8;
        ELSIF x =- 11253 THEN
            sigmoid_f := 8;
        ELSIF x =- 11252 THEN
            sigmoid_f := 8;
        ELSIF x =- 11251 THEN
            sigmoid_f := 8;
        ELSIF x =- 11250 THEN
            sigmoid_f := 8;
        ELSIF x =- 11249 THEN
            sigmoid_f := 8;
        ELSIF x =- 11248 THEN
            sigmoid_f := 8;
        ELSIF x =- 11247 THEN
            sigmoid_f := 8;
        ELSIF x =- 11246 THEN
            sigmoid_f := 8;
        ELSIF x =- 11245 THEN
            sigmoid_f := 8;
        ELSIF x =- 11244 THEN
            sigmoid_f := 8;
        ELSIF x =- 11243 THEN
            sigmoid_f := 8;
        ELSIF x =- 11242 THEN
            sigmoid_f := 8;
        ELSIF x =- 11241 THEN
            sigmoid_f := 8;
        ELSIF x =- 11240 THEN
            sigmoid_f := 8;
        ELSIF x =- 11239 THEN
            sigmoid_f := 8;
        ELSIF x =- 11238 THEN
            sigmoid_f := 8;
        ELSIF x =- 11237 THEN
            sigmoid_f := 8;
        ELSIF x =- 11236 THEN
            sigmoid_f := 8;
        ELSIF x =- 11235 THEN
            sigmoid_f := 8;
        ELSIF x =- 11234 THEN
            sigmoid_f := 8;
        ELSIF x =- 11233 THEN
            sigmoid_f := 8;
        ELSIF x =- 11232 THEN
            sigmoid_f := 8;
        ELSIF x =- 11231 THEN
            sigmoid_f := 8;
        ELSIF x =- 11230 THEN
            sigmoid_f := 8;
        ELSIF x =- 11229 THEN
            sigmoid_f := 8;
        ELSIF x =- 11228 THEN
            sigmoid_f := 8;
        ELSIF x =- 11227 THEN
            sigmoid_f := 8;
        ELSIF x =- 11226 THEN
            sigmoid_f := 8;
        ELSIF x =- 11225 THEN
            sigmoid_f := 8;
        ELSIF x =- 11224 THEN
            sigmoid_f := 8;
        ELSIF x =- 11223 THEN
            sigmoid_f := 8;
        ELSIF x =- 11222 THEN
            sigmoid_f := 8;
        ELSIF x =- 11221 THEN
            sigmoid_f := 8;
        ELSIF x =- 11220 THEN
            sigmoid_f := 8;
        ELSIF x =- 11219 THEN
            sigmoid_f := 8;
        ELSIF x =- 11218 THEN
            sigmoid_f := 8;
        ELSIF x =- 11217 THEN
            sigmoid_f := 8;
        ELSIF x =- 11216 THEN
            sigmoid_f := 8;
        ELSIF x =- 11215 THEN
            sigmoid_f := 8;
        ELSIF x =- 11214 THEN
            sigmoid_f := 8;
        ELSIF x =- 11213 THEN
            sigmoid_f := 8;
        ELSIF x =- 11212 THEN
            sigmoid_f := 8;
        ELSIF x =- 11211 THEN
            sigmoid_f := 8;
        ELSIF x =- 11210 THEN
            sigmoid_f := 8;
        ELSIF x =- 11209 THEN
            sigmoid_f := 8;
        ELSIF x =- 11208 THEN
            sigmoid_f := 8;
        ELSIF x =- 11207 THEN
            sigmoid_f := 8;
        ELSIF x =- 11206 THEN
            sigmoid_f := 8;
        ELSIF x =- 11205 THEN
            sigmoid_f := 8;
        ELSIF x =- 11204 THEN
            sigmoid_f := 8;
        ELSIF x =- 11203 THEN
            sigmoid_f := 8;
        ELSIF x =- 11202 THEN
            sigmoid_f := 8;
        ELSIF x =- 11201 THEN
            sigmoid_f := 8;
        ELSIF x =- 11200 THEN
            sigmoid_f := 8;
        ELSIF x =- 11199 THEN
            sigmoid_f := 8;
        ELSIF x =- 11198 THEN
            sigmoid_f := 8;
        ELSIF x =- 11197 THEN
            sigmoid_f := 8;
        ELSIF x =- 11196 THEN
            sigmoid_f := 8;
        ELSIF x =- 11195 THEN
            sigmoid_f := 8;
        ELSIF x =- 11194 THEN
            sigmoid_f := 8;
        ELSIF x =- 11193 THEN
            sigmoid_f := 8;
        ELSIF x =- 11192 THEN
            sigmoid_f := 8;
        ELSIF x =- 11191 THEN
            sigmoid_f := 8;
        ELSIF x =- 11190 THEN
            sigmoid_f := 8;
        ELSIF x =- 11189 THEN
            sigmoid_f := 8;
        ELSIF x =- 11188 THEN
            sigmoid_f := 8;
        ELSIF x =- 11187 THEN
            sigmoid_f := 8;
        ELSIF x =- 11186 THEN
            sigmoid_f := 8;
        ELSIF x =- 11185 THEN
            sigmoid_f := 8;
        ELSIF x =- 11184 THEN
            sigmoid_f := 8;
        ELSIF x =- 11183 THEN
            sigmoid_f := 8;
        ELSIF x =- 11182 THEN
            sigmoid_f := 8;
        ELSIF x =- 11181 THEN
            sigmoid_f := 8;
        ELSIF x =- 11180 THEN
            sigmoid_f := 8;
        ELSIF x =- 11179 THEN
            sigmoid_f := 8;
        ELSIF x =- 11178 THEN
            sigmoid_f := 8;
        ELSIF x =- 11177 THEN
            sigmoid_f := 8;
        ELSIF x =- 11176 THEN
            sigmoid_f := 8;
        ELSIF x =- 11175 THEN
            sigmoid_f := 8;
        ELSIF x =- 11174 THEN
            sigmoid_f := 8;
        ELSIF x =- 11173 THEN
            sigmoid_f := 8;
        ELSIF x =- 11172 THEN
            sigmoid_f := 8;
        ELSIF x =- 11171 THEN
            sigmoid_f := 8;
        ELSIF x =- 11170 THEN
            sigmoid_f := 8;
        ELSIF x =- 11169 THEN
            sigmoid_f := 8;
        ELSIF x =- 11168 THEN
            sigmoid_f := 8;
        ELSIF x =- 11167 THEN
            sigmoid_f := 8;
        ELSIF x =- 11166 THEN
            sigmoid_f := 8;
        ELSIF x =- 11165 THEN
            sigmoid_f := 8;
        ELSIF x =- 11164 THEN
            sigmoid_f := 8;
        ELSIF x =- 11163 THEN
            sigmoid_f := 8;
        ELSIF x =- 11162 THEN
            sigmoid_f := 8;
        ELSIF x =- 11161 THEN
            sigmoid_f := 8;
        ELSIF x =- 11160 THEN
            sigmoid_f := 8;
        ELSIF x =- 11159 THEN
            sigmoid_f := 8;
        ELSIF x =- 11158 THEN
            sigmoid_f := 8;
        ELSIF x =- 11157 THEN
            sigmoid_f := 8;
        ELSIF x =- 11156 THEN
            sigmoid_f := 8;
        ELSIF x =- 11155 THEN
            sigmoid_f := 8;
        ELSIF x =- 11154 THEN
            sigmoid_f := 8;
        ELSIF x =- 11153 THEN
            sigmoid_f := 8;
        ELSIF x =- 11152 THEN
            sigmoid_f := 8;
        ELSIF x =- 11151 THEN
            sigmoid_f := 8;
        ELSIF x =- 11150 THEN
            sigmoid_f := 8;
        ELSIF x =- 11149 THEN
            sigmoid_f := 8;
        ELSIF x =- 11148 THEN
            sigmoid_f := 8;
        ELSIF x =- 11147 THEN
            sigmoid_f := 8;
        ELSIF x =- 11146 THEN
            sigmoid_f := 8;
        ELSIF x =- 11145 THEN
            sigmoid_f := 8;
        ELSIF x =- 11144 THEN
            sigmoid_f := 8;
        ELSIF x =- 11143 THEN
            sigmoid_f := 8;
        ELSIF x =- 11142 THEN
            sigmoid_f := 8;
        ELSIF x =- 11141 THEN
            sigmoid_f := 8;
        ELSIF x =- 11140 THEN
            sigmoid_f := 8;
        ELSIF x =- 11139 THEN
            sigmoid_f := 8;
        ELSIF x =- 11138 THEN
            sigmoid_f := 8;
        ELSIF x =- 11137 THEN
            sigmoid_f := 8;
        ELSIF x =- 11136 THEN
            sigmoid_f := 8;
        ELSIF x =- 11135 THEN
            sigmoid_f := 8;
        ELSIF x =- 11134 THEN
            sigmoid_f := 8;
        ELSIF x =- 11133 THEN
            sigmoid_f := 8;
        ELSIF x =- 11132 THEN
            sigmoid_f := 8;
        ELSIF x =- 11131 THEN
            sigmoid_f := 8;
        ELSIF x =- 11130 THEN
            sigmoid_f := 8;
        ELSIF x =- 11129 THEN
            sigmoid_f := 8;
        ELSIF x =- 11128 THEN
            sigmoid_f := 8;
        ELSIF x =- 11127 THEN
            sigmoid_f := 8;
        ELSIF x =- 11126 THEN
            sigmoid_f := 8;
        ELSIF x =- 11125 THEN
            sigmoid_f := 8;
        ELSIF x =- 11124 THEN
            sigmoid_f := 8;
        ELSIF x =- 11123 THEN
            sigmoid_f := 8;
        ELSIF x =- 11122 THEN
            sigmoid_f := 8;
        ELSIF x =- 11121 THEN
            sigmoid_f := 8;
        ELSIF x =- 11120 THEN
            sigmoid_f := 8;
        ELSIF x =- 11119 THEN
            sigmoid_f := 8;
        ELSIF x =- 11118 THEN
            sigmoid_f := 8;
        ELSIF x =- 11117 THEN
            sigmoid_f := 8;
        ELSIF x =- 11116 THEN
            sigmoid_f := 8;
        ELSIF x =- 11115 THEN
            sigmoid_f := 8;
        ELSIF x =- 11114 THEN
            sigmoid_f := 8;
        ELSIF x =- 11113 THEN
            sigmoid_f := 8;
        ELSIF x =- 11112 THEN
            sigmoid_f := 8;
        ELSIF x =- 11111 THEN
            sigmoid_f := 8;
        ELSIF x =- 11110 THEN
            sigmoid_f := 8;
        ELSIF x =- 11109 THEN
            sigmoid_f := 8;
        ELSIF x =- 11108 THEN
            sigmoid_f := 8;
        ELSIF x =- 11107 THEN
            sigmoid_f := 8;
        ELSIF x =- 11106 THEN
            sigmoid_f := 8;
        ELSIF x =- 11105 THEN
            sigmoid_f := 8;
        ELSIF x =- 11104 THEN
            sigmoid_f := 8;
        ELSIF x =- 11103 THEN
            sigmoid_f := 8;
        ELSIF x =- 11102 THEN
            sigmoid_f := 8;
        ELSIF x =- 11101 THEN
            sigmoid_f := 8;
        ELSIF x =- 11100 THEN
            sigmoid_f := 8;
        ELSIF x =- 11099 THEN
            sigmoid_f := 8;
        ELSIF x =- 11098 THEN
            sigmoid_f := 8;
        ELSIF x =- 11097 THEN
            sigmoid_f := 8;
        ELSIF x =- 11096 THEN
            sigmoid_f := 8;
        ELSIF x =- 11095 THEN
            sigmoid_f := 8;
        ELSIF x =- 11094 THEN
            sigmoid_f := 8;
        ELSIF x =- 11093 THEN
            sigmoid_f := 9;
        ELSIF x =- 11092 THEN
            sigmoid_f := 9;
        ELSIF x =- 11091 THEN
            sigmoid_f := 9;
        ELSIF x =- 11090 THEN
            sigmoid_f := 9;
        ELSIF x =- 11089 THEN
            sigmoid_f := 9;
        ELSIF x =- 11088 THEN
            sigmoid_f := 9;
        ELSIF x =- 11087 THEN
            sigmoid_f := 9;
        ELSIF x =- 11086 THEN
            sigmoid_f := 9;
        ELSIF x =- 11085 THEN
            sigmoid_f := 9;
        ELSIF x =- 11084 THEN
            sigmoid_f := 9;
        ELSIF x =- 11083 THEN
            sigmoid_f := 9;
        ELSIF x =- 11082 THEN
            sigmoid_f := 9;
        ELSIF x =- 11081 THEN
            sigmoid_f := 9;
        ELSIF x =- 11080 THEN
            sigmoid_f := 9;
        ELSIF x =- 11079 THEN
            sigmoid_f := 9;
        ELSIF x =- 11078 THEN
            sigmoid_f := 9;
        ELSIF x =- 11077 THEN
            sigmoid_f := 9;
        ELSIF x =- 11076 THEN
            sigmoid_f := 9;
        ELSIF x =- 11075 THEN
            sigmoid_f := 9;
        ELSIF x =- 11074 THEN
            sigmoid_f := 9;
        ELSIF x =- 11073 THEN
            sigmoid_f := 9;
        ELSIF x =- 11072 THEN
            sigmoid_f := 9;
        ELSIF x =- 11071 THEN
            sigmoid_f := 9;
        ELSIF x =- 11070 THEN
            sigmoid_f := 9;
        ELSIF x =- 11069 THEN
            sigmoid_f := 9;
        ELSIF x =- 11068 THEN
            sigmoid_f := 9;
        ELSIF x =- 11067 THEN
            sigmoid_f := 9;
        ELSIF x =- 11066 THEN
            sigmoid_f := 9;
        ELSIF x =- 11065 THEN
            sigmoid_f := 9;
        ELSIF x =- 11064 THEN
            sigmoid_f := 9;
        ELSIF x =- 11063 THEN
            sigmoid_f := 9;
        ELSIF x =- 11062 THEN
            sigmoid_f := 9;
        ELSIF x =- 11061 THEN
            sigmoid_f := 9;
        ELSIF x =- 11060 THEN
            sigmoid_f := 9;
        ELSIF x =- 11059 THEN
            sigmoid_f := 9;
        ELSIF x =- 11058 THEN
            sigmoid_f := 9;
        ELSIF x =- 11057 THEN
            sigmoid_f := 9;
        ELSIF x =- 11056 THEN
            sigmoid_f := 9;
        ELSIF x =- 11055 THEN
            sigmoid_f := 9;
        ELSIF x =- 11054 THEN
            sigmoid_f := 9;
        ELSIF x =- 11053 THEN
            sigmoid_f := 9;
        ELSIF x =- 11052 THEN
            sigmoid_f := 9;
        ELSIF x =- 11051 THEN
            sigmoid_f := 9;
        ELSIF x =- 11050 THEN
            sigmoid_f := 9;
        ELSIF x =- 11049 THEN
            sigmoid_f := 9;
        ELSIF x =- 11048 THEN
            sigmoid_f := 9;
        ELSIF x =- 11047 THEN
            sigmoid_f := 9;
        ELSIF x =- 11046 THEN
            sigmoid_f := 9;
        ELSIF x =- 11045 THEN
            sigmoid_f := 9;
        ELSIF x =- 11044 THEN
            sigmoid_f := 9;
        ELSIF x =- 11043 THEN
            sigmoid_f := 9;
        ELSIF x =- 11042 THEN
            sigmoid_f := 9;
        ELSIF x =- 11041 THEN
            sigmoid_f := 9;
        ELSIF x =- 11040 THEN
            sigmoid_f := 9;
        ELSIF x =- 11039 THEN
            sigmoid_f := 9;
        ELSIF x =- 11038 THEN
            sigmoid_f := 9;
        ELSIF x =- 11037 THEN
            sigmoid_f := 9;
        ELSIF x =- 11036 THEN
            sigmoid_f := 9;
        ELSIF x =- 11035 THEN
            sigmoid_f := 9;
        ELSIF x =- 11034 THEN
            sigmoid_f := 9;
        ELSIF x =- 11033 THEN
            sigmoid_f := 9;
        ELSIF x =- 11032 THEN
            sigmoid_f := 9;
        ELSIF x =- 11031 THEN
            sigmoid_f := 9;
        ELSIF x =- 11030 THEN
            sigmoid_f := 9;
        ELSIF x =- 11029 THEN
            sigmoid_f := 9;
        ELSIF x =- 11028 THEN
            sigmoid_f := 9;
        ELSIF x =- 11027 THEN
            sigmoid_f := 9;
        ELSIF x =- 11026 THEN
            sigmoid_f := 9;
        ELSIF x =- 11025 THEN
            sigmoid_f := 9;
        ELSIF x =- 11024 THEN
            sigmoid_f := 9;
        ELSIF x =- 11023 THEN
            sigmoid_f := 9;
        ELSIF x =- 11022 THEN
            sigmoid_f := 9;
        ELSIF x =- 11021 THEN
            sigmoid_f := 9;
        ELSIF x =- 11020 THEN
            sigmoid_f := 9;
        ELSIF x =- 11019 THEN
            sigmoid_f := 9;
        ELSIF x =- 11018 THEN
            sigmoid_f := 9;
        ELSIF x =- 11017 THEN
            sigmoid_f := 9;
        ELSIF x =- 11016 THEN
            sigmoid_f := 9;
        ELSIF x =- 11015 THEN
            sigmoid_f := 9;
        ELSIF x =- 11014 THEN
            sigmoid_f := 9;
        ELSIF x =- 11013 THEN
            sigmoid_f := 9;
        ELSIF x =- 11012 THEN
            sigmoid_f := 9;
        ELSIF x =- 11011 THEN
            sigmoid_f := 9;
        ELSIF x =- 11010 THEN
            sigmoid_f := 9;
        ELSIF x =- 11009 THEN
            sigmoid_f := 9;
        ELSIF x =- 11008 THEN
            sigmoid_f := 9;
        ELSIF x =- 11007 THEN
            sigmoid_f := 9;
        ELSIF x =- 11006 THEN
            sigmoid_f := 9;
        ELSIF x =- 11005 THEN
            sigmoid_f := 9;
        ELSIF x =- 11004 THEN
            sigmoid_f := 9;
        ELSIF x =- 11003 THEN
            sigmoid_f := 9;
        ELSIF x =- 11002 THEN
            sigmoid_f := 9;
        ELSIF x =- 11001 THEN
            sigmoid_f := 9;
        ELSIF x =- 11000 THEN
            sigmoid_f := 9;
        ELSIF x =- 10999 THEN
            sigmoid_f := 9;
        ELSIF x =- 10998 THEN
            sigmoid_f := 9;
        ELSIF x =- 10997 THEN
            sigmoid_f := 9;
        ELSIF x =- 10996 THEN
            sigmoid_f := 9;
        ELSIF x =- 10995 THEN
            sigmoid_f := 9;
        ELSIF x =- 10994 THEN
            sigmoid_f := 9;
        ELSIF x =- 10993 THEN
            sigmoid_f := 9;
        ELSIF x =- 10992 THEN
            sigmoid_f := 9;
        ELSIF x =- 10991 THEN
            sigmoid_f := 9;
        ELSIF x =- 10990 THEN
            sigmoid_f := 9;
        ELSIF x =- 10989 THEN
            sigmoid_f := 9;
        ELSIF x =- 10988 THEN
            sigmoid_f := 9;
        ELSIF x =- 10987 THEN
            sigmoid_f := 9;
        ELSIF x =- 10986 THEN
            sigmoid_f := 9;
        ELSIF x =- 10985 THEN
            sigmoid_f := 9;
        ELSIF x =- 10984 THEN
            sigmoid_f := 9;
        ELSIF x =- 10983 THEN
            sigmoid_f := 9;
        ELSIF x =- 10982 THEN
            sigmoid_f := 9;
        ELSIF x =- 10981 THEN
            sigmoid_f := 9;
        ELSIF x =- 10980 THEN
            sigmoid_f := 9;
        ELSIF x =- 10979 THEN
            sigmoid_f := 9;
        ELSIF x =- 10978 THEN
            sigmoid_f := 9;
        ELSIF x =- 10977 THEN
            sigmoid_f := 9;
        ELSIF x =- 10976 THEN
            sigmoid_f := 9;
        ELSIF x =- 10975 THEN
            sigmoid_f := 9;
        ELSIF x =- 10974 THEN
            sigmoid_f := 9;
        ELSIF x =- 10973 THEN
            sigmoid_f := 9;
        ELSIF x =- 10972 THEN
            sigmoid_f := 9;
        ELSIF x =- 10971 THEN
            sigmoid_f := 9;
        ELSIF x =- 10970 THEN
            sigmoid_f := 9;
        ELSIF x =- 10969 THEN
            sigmoid_f := 9;
        ELSIF x =- 10968 THEN
            sigmoid_f := 9;
        ELSIF x =- 10967 THEN
            sigmoid_f := 9;
        ELSIF x =- 10966 THEN
            sigmoid_f := 9;
        ELSIF x =- 10965 THEN
            sigmoid_f := 9;
        ELSIF x =- 10964 THEN
            sigmoid_f := 9;
        ELSIF x =- 10963 THEN
            sigmoid_f := 9;
        ELSIF x =- 10962 THEN
            sigmoid_f := 9;
        ELSIF x =- 10961 THEN
            sigmoid_f := 9;
        ELSIF x =- 10960 THEN
            sigmoid_f := 9;
        ELSIF x =- 10959 THEN
            sigmoid_f := 9;
        ELSIF x =- 10958 THEN
            sigmoid_f := 9;
        ELSIF x =- 10957 THEN
            sigmoid_f := 9;
        ELSIF x =- 10956 THEN
            sigmoid_f := 9;
        ELSIF x =- 10955 THEN
            sigmoid_f := 9;
        ELSIF x =- 10954 THEN
            sigmoid_f := 9;
        ELSIF x =- 10953 THEN
            sigmoid_f := 9;
        ELSIF x =- 10952 THEN
            sigmoid_f := 9;
        ELSIF x =- 10951 THEN
            sigmoid_f := 9;
        ELSIF x =- 10950 THEN
            sigmoid_f := 9;
        ELSIF x =- 10949 THEN
            sigmoid_f := 9;
        ELSIF x =- 10948 THEN
            sigmoid_f := 9;
        ELSIF x =- 10947 THEN
            sigmoid_f := 9;
        ELSIF x =- 10946 THEN
            sigmoid_f := 9;
        ELSIF x =- 10945 THEN
            sigmoid_f := 9;
        ELSIF x =- 10944 THEN
            sigmoid_f := 9;
        ELSIF x =- 10943 THEN
            sigmoid_f := 9;
        ELSIF x =- 10942 THEN
            sigmoid_f := 9;
        ELSIF x =- 10941 THEN
            sigmoid_f := 9;
        ELSIF x =- 10940 THEN
            sigmoid_f := 9;
        ELSIF x =- 10939 THEN
            sigmoid_f := 9;
        ELSIF x =- 10938 THEN
            sigmoid_f := 9;
        ELSIF x =- 10937 THEN
            sigmoid_f := 9;
        ELSIF x =- 10936 THEN
            sigmoid_f := 9;
        ELSIF x =- 10935 THEN
            sigmoid_f := 9;
        ELSIF x =- 10934 THEN
            sigmoid_f := 9;
        ELSIF x =- 10933 THEN
            sigmoid_f := 9;
        ELSIF x =- 10932 THEN
            sigmoid_f := 9;
        ELSIF x =- 10931 THEN
            sigmoid_f := 9;
        ELSIF x =- 10930 THEN
            sigmoid_f := 9;
        ELSIF x =- 10929 THEN
            sigmoid_f := 9;
        ELSIF x =- 10928 THEN
            sigmoid_f := 9;
        ELSIF x =- 10927 THEN
            sigmoid_f := 9;
        ELSIF x =- 10926 THEN
            sigmoid_f := 9;
        ELSIF x =- 10925 THEN
            sigmoid_f := 9;
        ELSIF x =- 10924 THEN
            sigmoid_f := 9;
        ELSIF x =- 10923 THEN
            sigmoid_f := 9;
        ELSIF x =- 10922 THEN
            sigmoid_f := 10;
        ELSIF x =- 10921 THEN
            sigmoid_f := 10;
        ELSIF x =- 10920 THEN
            sigmoid_f := 10;
        ELSIF x =- 10919 THEN
            sigmoid_f := 10;
        ELSIF x =- 10918 THEN
            sigmoid_f := 10;
        ELSIF x =- 10917 THEN
            sigmoid_f := 10;
        ELSIF x =- 10916 THEN
            sigmoid_f := 10;
        ELSIF x =- 10915 THEN
            sigmoid_f := 10;
        ELSIF x =- 10914 THEN
            sigmoid_f := 10;
        ELSIF x =- 10913 THEN
            sigmoid_f := 10;
        ELSIF x =- 10912 THEN
            sigmoid_f := 10;
        ELSIF x =- 10911 THEN
            sigmoid_f := 10;
        ELSIF x =- 10910 THEN
            sigmoid_f := 10;
        ELSIF x =- 10909 THEN
            sigmoid_f := 10;
        ELSIF x =- 10908 THEN
            sigmoid_f := 10;
        ELSIF x =- 10907 THEN
            sigmoid_f := 10;
        ELSIF x =- 10906 THEN
            sigmoid_f := 10;
        ELSIF x =- 10905 THEN
            sigmoid_f := 10;
        ELSIF x =- 10904 THEN
            sigmoid_f := 10;
        ELSIF x =- 10903 THEN
            sigmoid_f := 10;
        ELSIF x =- 10902 THEN
            sigmoid_f := 10;
        ELSIF x =- 10901 THEN
            sigmoid_f := 10;
        ELSIF x =- 10900 THEN
            sigmoid_f := 10;
        ELSIF x =- 10899 THEN
            sigmoid_f := 10;
        ELSIF x =- 10898 THEN
            sigmoid_f := 10;
        ELSIF x =- 10897 THEN
            sigmoid_f := 10;
        ELSIF x =- 10896 THEN
            sigmoid_f := 10;
        ELSIF x =- 10895 THEN
            sigmoid_f := 10;
        ELSIF x =- 10894 THEN
            sigmoid_f := 10;
        ELSIF x =- 10893 THEN
            sigmoid_f := 10;
        ELSIF x =- 10892 THEN
            sigmoid_f := 10;
        ELSIF x =- 10891 THEN
            sigmoid_f := 10;
        ELSIF x =- 10890 THEN
            sigmoid_f := 10;
        ELSIF x =- 10889 THEN
            sigmoid_f := 10;
        ELSIF x =- 10888 THEN
            sigmoid_f := 10;
        ELSIF x =- 10887 THEN
            sigmoid_f := 10;
        ELSIF x =- 10886 THEN
            sigmoid_f := 10;
        ELSIF x =- 10885 THEN
            sigmoid_f := 10;
        ELSIF x =- 10884 THEN
            sigmoid_f := 10;
        ELSIF x =- 10883 THEN
            sigmoid_f := 10;
        ELSIF x =- 10882 THEN
            sigmoid_f := 10;
        ELSIF x =- 10881 THEN
            sigmoid_f := 10;
        ELSIF x =- 10880 THEN
            sigmoid_f := 10;
        ELSIF x =- 10879 THEN
            sigmoid_f := 10;
        ELSIF x =- 10878 THEN
            sigmoid_f := 10;
        ELSIF x =- 10877 THEN
            sigmoid_f := 10;
        ELSIF x =- 10876 THEN
            sigmoid_f := 10;
        ELSIF x =- 10875 THEN
            sigmoid_f := 10;
        ELSIF x =- 10874 THEN
            sigmoid_f := 10;
        ELSIF x =- 10873 THEN
            sigmoid_f := 10;
        ELSIF x =- 10872 THEN
            sigmoid_f := 10;
        ELSIF x =- 10871 THEN
            sigmoid_f := 10;
        ELSIF x =- 10870 THEN
            sigmoid_f := 10;
        ELSIF x =- 10869 THEN
            sigmoid_f := 10;
        ELSIF x =- 10868 THEN
            sigmoid_f := 10;
        ELSIF x =- 10867 THEN
            sigmoid_f := 10;
        ELSIF x =- 10866 THEN
            sigmoid_f := 10;
        ELSIF x =- 10865 THEN
            sigmoid_f := 10;
        ELSIF x =- 10864 THEN
            sigmoid_f := 10;
        ELSIF x =- 10863 THEN
            sigmoid_f := 10;
        ELSIF x =- 10862 THEN
            sigmoid_f := 10;
        ELSIF x =- 10861 THEN
            sigmoid_f := 10;
        ELSIF x =- 10860 THEN
            sigmoid_f := 10;
        ELSIF x =- 10859 THEN
            sigmoid_f := 10;
        ELSIF x =- 10858 THEN
            sigmoid_f := 10;
        ELSIF x =- 10857 THEN
            sigmoid_f := 10;
        ELSIF x =- 10856 THEN
            sigmoid_f := 10;
        ELSIF x =- 10855 THEN
            sigmoid_f := 10;
        ELSIF x =- 10854 THEN
            sigmoid_f := 10;
        ELSIF x =- 10853 THEN
            sigmoid_f := 10;
        ELSIF x =- 10852 THEN
            sigmoid_f := 10;
        ELSIF x =- 10851 THEN
            sigmoid_f := 10;
        ELSIF x =- 10850 THEN
            sigmoid_f := 10;
        ELSIF x =- 10849 THEN
            sigmoid_f := 10;
        ELSIF x =- 10848 THEN
            sigmoid_f := 10;
        ELSIF x =- 10847 THEN
            sigmoid_f := 10;
        ELSIF x =- 10846 THEN
            sigmoid_f := 10;
        ELSIF x =- 10845 THEN
            sigmoid_f := 10;
        ELSIF x =- 10844 THEN
            sigmoid_f := 10;
        ELSIF x =- 10843 THEN
            sigmoid_f := 10;
        ELSIF x =- 10842 THEN
            sigmoid_f := 10;
        ELSIF x =- 10841 THEN
            sigmoid_f := 10;
        ELSIF x =- 10840 THEN
            sigmoid_f := 10;
        ELSIF x =- 10839 THEN
            sigmoid_f := 10;
        ELSIF x =- 10838 THEN
            sigmoid_f := 10;
        ELSIF x =- 10837 THEN
            sigmoid_f := 10;
        ELSIF x =- 10836 THEN
            sigmoid_f := 10;
        ELSIF x =- 10835 THEN
            sigmoid_f := 10;
        ELSIF x =- 10834 THEN
            sigmoid_f := 10;
        ELSIF x =- 10833 THEN
            sigmoid_f := 10;
        ELSIF x =- 10832 THEN
            sigmoid_f := 10;
        ELSIF x =- 10831 THEN
            sigmoid_f := 10;
        ELSIF x =- 10830 THEN
            sigmoid_f := 10;
        ELSIF x =- 10829 THEN
            sigmoid_f := 10;
        ELSIF x =- 10828 THEN
            sigmoid_f := 10;
        ELSIF x =- 10827 THEN
            sigmoid_f := 10;
        ELSIF x =- 10826 THEN
            sigmoid_f := 10;
        ELSIF x =- 10825 THEN
            sigmoid_f := 10;
        ELSIF x =- 10824 THEN
            sigmoid_f := 10;
        ELSIF x =- 10823 THEN
            sigmoid_f := 10;
        ELSIF x =- 10822 THEN
            sigmoid_f := 10;
        ELSIF x =- 10821 THEN
            sigmoid_f := 10;
        ELSIF x =- 10820 THEN
            sigmoid_f := 10;
        ELSIF x =- 10819 THEN
            sigmoid_f := 10;
        ELSIF x =- 10818 THEN
            sigmoid_f := 10;
        ELSIF x =- 10817 THEN
            sigmoid_f := 10;
        ELSIF x =- 10816 THEN
            sigmoid_f := 10;
        ELSIF x =- 10815 THEN
            sigmoid_f := 10;
        ELSIF x =- 10814 THEN
            sigmoid_f := 10;
        ELSIF x =- 10813 THEN
            sigmoid_f := 10;
        ELSIF x =- 10812 THEN
            sigmoid_f := 10;
        ELSIF x =- 10811 THEN
            sigmoid_f := 10;
        ELSIF x =- 10810 THEN
            sigmoid_f := 10;
        ELSIF x =- 10809 THEN
            sigmoid_f := 10;
        ELSIF x =- 10808 THEN
            sigmoid_f := 10;
        ELSIF x =- 10807 THEN
            sigmoid_f := 10;
        ELSIF x =- 10806 THEN
            sigmoid_f := 10;
        ELSIF x =- 10805 THEN
            sigmoid_f := 10;
        ELSIF x =- 10804 THEN
            sigmoid_f := 10;
        ELSIF x =- 10803 THEN
            sigmoid_f := 10;
        ELSIF x =- 10802 THEN
            sigmoid_f := 10;
        ELSIF x =- 10801 THEN
            sigmoid_f := 10;
        ELSIF x =- 10800 THEN
            sigmoid_f := 10;
        ELSIF x =- 10799 THEN
            sigmoid_f := 10;
        ELSIF x =- 10798 THEN
            sigmoid_f := 10;
        ELSIF x =- 10797 THEN
            sigmoid_f := 10;
        ELSIF x =- 10796 THEN
            sigmoid_f := 10;
        ELSIF x =- 10795 THEN
            sigmoid_f := 10;
        ELSIF x =- 10794 THEN
            sigmoid_f := 10;
        ELSIF x =- 10793 THEN
            sigmoid_f := 10;
        ELSIF x =- 10792 THEN
            sigmoid_f := 10;
        ELSIF x =- 10791 THEN
            sigmoid_f := 10;
        ELSIF x =- 10790 THEN
            sigmoid_f := 10;
        ELSIF x =- 10789 THEN
            sigmoid_f := 10;
        ELSIF x =- 10788 THEN
            sigmoid_f := 10;
        ELSIF x =- 10787 THEN
            sigmoid_f := 10;
        ELSIF x =- 10786 THEN
            sigmoid_f := 10;
        ELSIF x =- 10785 THEN
            sigmoid_f := 10;
        ELSIF x =- 10784 THEN
            sigmoid_f := 10;
        ELSIF x =- 10783 THEN
            sigmoid_f := 10;
        ELSIF x =- 10782 THEN
            sigmoid_f := 10;
        ELSIF x =- 10781 THEN
            sigmoid_f := 10;
        ELSIF x =- 10780 THEN
            sigmoid_f := 10;
        ELSIF x =- 10779 THEN
            sigmoid_f := 10;
        ELSIF x =- 10778 THEN
            sigmoid_f := 10;
        ELSIF x =- 10777 THEN
            sigmoid_f := 10;
        ELSIF x =- 10776 THEN
            sigmoid_f := 10;
        ELSIF x =- 10775 THEN
            sigmoid_f := 10;
        ELSIF x =- 10774 THEN
            sigmoid_f := 10;
        ELSIF x =- 10773 THEN
            sigmoid_f := 10;
        ELSIF x =- 10772 THEN
            sigmoid_f := 10;
        ELSIF x =- 10771 THEN
            sigmoid_f := 10;
        ELSIF x =- 10770 THEN
            sigmoid_f := 10;
        ELSIF x =- 10769 THEN
            sigmoid_f := 10;
        ELSIF x =- 10768 THEN
            sigmoid_f := 10;
        ELSIF x =- 10767 THEN
            sigmoid_f := 10;
        ELSIF x =- 10766 THEN
            sigmoid_f := 10;
        ELSIF x =- 10765 THEN
            sigmoid_f := 10;
        ELSIF x =- 10764 THEN
            sigmoid_f := 10;
        ELSIF x =- 10763 THEN
            sigmoid_f := 10;
        ELSIF x =- 10762 THEN
            sigmoid_f := 10;
        ELSIF x =- 10761 THEN
            sigmoid_f := 10;
        ELSIF x =- 10760 THEN
            sigmoid_f := 10;
        ELSIF x =- 10759 THEN
            sigmoid_f := 10;
        ELSIF x =- 10758 THEN
            sigmoid_f := 10;
        ELSIF x =- 10757 THEN
            sigmoid_f := 10;
        ELSIF x =- 10756 THEN
            sigmoid_f := 10;
        ELSIF x =- 10755 THEN
            sigmoid_f := 10;
        ELSIF x =- 10754 THEN
            sigmoid_f := 10;
        ELSIF x =- 10753 THEN
            sigmoid_f := 10;
        ELSIF x =- 10752 THEN
            sigmoid_f := 11;
        ELSIF x =- 10751 THEN
            sigmoid_f := 10;
        ELSIF x =- 10750 THEN
            sigmoid_f := 10;
        ELSIF x =- 10749 THEN
            sigmoid_f := 10;
        ELSIF x =- 10748 THEN
            sigmoid_f := 10;
        ELSIF x =- 10747 THEN
            sigmoid_f := 10;
        ELSIF x =- 10746 THEN
            sigmoid_f := 10;
        ELSIF x =- 10745 THEN
            sigmoid_f := 10;
        ELSIF x =- 10744 THEN
            sigmoid_f := 10;
        ELSIF x =- 10743 THEN
            sigmoid_f := 10;
        ELSIF x =- 10742 THEN
            sigmoid_f := 10;
        ELSIF x =- 10741 THEN
            sigmoid_f := 10;
        ELSIF x =- 10740 THEN
            sigmoid_f := 10;
        ELSIF x =- 10739 THEN
            sigmoid_f := 10;
        ELSIF x =- 10738 THEN
            sigmoid_f := 10;
        ELSIF x =- 10737 THEN
            sigmoid_f := 10;
        ELSIF x =- 10736 THEN
            sigmoid_f := 10;
        ELSIF x =- 10735 THEN
            sigmoid_f := 10;
        ELSIF x =- 10734 THEN
            sigmoid_f := 10;
        ELSIF x =- 10733 THEN
            sigmoid_f := 10;
        ELSIF x =- 10732 THEN
            sigmoid_f := 10;
        ELSIF x =- 10731 THEN
            sigmoid_f := 10;
        ELSIF x =- 10730 THEN
            sigmoid_f := 10;
        ELSIF x =- 10729 THEN
            sigmoid_f := 10;
        ELSIF x =- 10728 THEN
            sigmoid_f := 10;
        ELSIF x =- 10727 THEN
            sigmoid_f := 10;
        ELSIF x =- 10726 THEN
            sigmoid_f := 10;
        ELSIF x =- 10725 THEN
            sigmoid_f := 10;
        ELSIF x =- 10724 THEN
            sigmoid_f := 10;
        ELSIF x =- 10723 THEN
            sigmoid_f := 10;
        ELSIF x =- 10722 THEN
            sigmoid_f := 10;
        ELSIF x =- 10721 THEN
            sigmoid_f := 10;
        ELSIF x =- 10720 THEN
            sigmoid_f := 10;
        ELSIF x =- 10719 THEN
            sigmoid_f := 10;
        ELSIF x =- 10718 THEN
            sigmoid_f := 10;
        ELSIF x =- 10717 THEN
            sigmoid_f := 10;
        ELSIF x =- 10716 THEN
            sigmoid_f := 10;
        ELSIF x =- 10715 THEN
            sigmoid_f := 10;
        ELSIF x =- 10714 THEN
            sigmoid_f := 10;
        ELSIF x =- 10713 THEN
            sigmoid_f := 10;
        ELSIF x =- 10712 THEN
            sigmoid_f := 10;
        ELSIF x =- 10711 THEN
            sigmoid_f := 10;
        ELSIF x =- 10710 THEN
            sigmoid_f := 10;
        ELSIF x =- 10709 THEN
            sigmoid_f := 10;
        ELSIF x =- 10708 THEN
            sigmoid_f := 10;
        ELSIF x =- 10707 THEN
            sigmoid_f := 10;
        ELSIF x =- 10706 THEN
            sigmoid_f := 10;
        ELSIF x =- 10705 THEN
            sigmoid_f := 10;
        ELSIF x =- 10704 THEN
            sigmoid_f := 10;
        ELSIF x =- 10703 THEN
            sigmoid_f := 10;
        ELSIF x =- 10702 THEN
            sigmoid_f := 10;
        ELSIF x =- 10701 THEN
            sigmoid_f := 10;
        ELSIF x =- 10700 THEN
            sigmoid_f := 10;
        ELSIF x =- 10699 THEN
            sigmoid_f := 10;
        ELSIF x =- 10698 THEN
            sigmoid_f := 10;
        ELSIF x =- 10697 THEN
            sigmoid_f := 10;
        ELSIF x =- 10696 THEN
            sigmoid_f := 10;
        ELSIF x =- 10695 THEN
            sigmoid_f := 10;
        ELSIF x =- 10694 THEN
            sigmoid_f := 10;
        ELSIF x =- 10693 THEN
            sigmoid_f := 10;
        ELSIF x =- 10692 THEN
            sigmoid_f := 10;
        ELSIF x =- 10691 THEN
            sigmoid_f := 10;
        ELSIF x =- 10690 THEN
            sigmoid_f := 10;
        ELSIF x =- 10689 THEN
            sigmoid_f := 10;
        ELSIF x =- 10688 THEN
            sigmoid_f := 10;
        ELSIF x =- 10687 THEN
            sigmoid_f := 10;
        ELSIF x =- 10686 THEN
            sigmoid_f := 10;
        ELSIF x =- 10685 THEN
            sigmoid_f := 10;
        ELSIF x =- 10684 THEN
            sigmoid_f := 10;
        ELSIF x =- 10683 THEN
            sigmoid_f := 10;
        ELSIF x =- 10682 THEN
            sigmoid_f := 10;
        ELSIF x =- 10681 THEN
            sigmoid_f := 10;
        ELSIF x =- 10680 THEN
            sigmoid_f := 10;
        ELSIF x =- 10679 THEN
            sigmoid_f := 10;
        ELSIF x =- 10678 THEN
            sigmoid_f := 11;
        ELSIF x =- 10677 THEN
            sigmoid_f := 11;
        ELSIF x =- 10676 THEN
            sigmoid_f := 11;
        ELSIF x =- 10675 THEN
            sigmoid_f := 11;
        ELSIF x =- 10674 THEN
            sigmoid_f := 11;
        ELSIF x =- 10673 THEN
            sigmoid_f := 11;
        ELSIF x =- 10672 THEN
            sigmoid_f := 11;
        ELSIF x =- 10671 THEN
            sigmoid_f := 11;
        ELSIF x =- 10670 THEN
            sigmoid_f := 11;
        ELSIF x =- 10669 THEN
            sigmoid_f := 11;
        ELSIF x =- 10668 THEN
            sigmoid_f := 11;
        ELSIF x =- 10667 THEN
            sigmoid_f := 11;
        ELSIF x =- 10666 THEN
            sigmoid_f := 11;
        ELSIF x =- 10665 THEN
            sigmoid_f := 11;
        ELSIF x =- 10664 THEN
            sigmoid_f := 11;
        ELSIF x =- 10663 THEN
            sigmoid_f := 11;
        ELSIF x =- 10662 THEN
            sigmoid_f := 11;
        ELSIF x =- 10661 THEN
            sigmoid_f := 11;
        ELSIF x =- 10660 THEN
            sigmoid_f := 11;
        ELSIF x =- 10659 THEN
            sigmoid_f := 11;
        ELSIF x =- 10658 THEN
            sigmoid_f := 11;
        ELSIF x =- 10657 THEN
            sigmoid_f := 11;
        ELSIF x =- 10656 THEN
            sigmoid_f := 11;
        ELSIF x =- 10655 THEN
            sigmoid_f := 11;
        ELSIF x =- 10654 THEN
            sigmoid_f := 11;
        ELSIF x =- 10653 THEN
            sigmoid_f := 11;
        ELSIF x =- 10652 THEN
            sigmoid_f := 11;
        ELSIF x =- 10651 THEN
            sigmoid_f := 11;
        ELSIF x =- 10650 THEN
            sigmoid_f := 11;
        ELSIF x =- 10649 THEN
            sigmoid_f := 11;
        ELSIF x =- 10648 THEN
            sigmoid_f := 11;
        ELSIF x =- 10647 THEN
            sigmoid_f := 11;
        ELSIF x =- 10646 THEN
            sigmoid_f := 11;
        ELSIF x =- 10645 THEN
            sigmoid_f := 11;
        ELSIF x =- 10644 THEN
            sigmoid_f := 11;
        ELSIF x =- 10643 THEN
            sigmoid_f := 11;
        ELSIF x =- 10642 THEN
            sigmoid_f := 11;
        ELSIF x =- 10641 THEN
            sigmoid_f := 11;
        ELSIF x =- 10640 THEN
            sigmoid_f := 11;
        ELSIF x =- 10639 THEN
            sigmoid_f := 11;
        ELSIF x =- 10638 THEN
            sigmoid_f := 11;
        ELSIF x =- 10637 THEN
            sigmoid_f := 11;
        ELSIF x =- 10636 THEN
            sigmoid_f := 11;
        ELSIF x =- 10635 THEN
            sigmoid_f := 11;
        ELSIF x =- 10634 THEN
            sigmoid_f := 11;
        ELSIF x =- 10633 THEN
            sigmoid_f := 11;
        ELSIF x =- 10632 THEN
            sigmoid_f := 11;
        ELSIF x =- 10631 THEN
            sigmoid_f := 11;
        ELSIF x =- 10630 THEN
            sigmoid_f := 11;
        ELSIF x =- 10629 THEN
            sigmoid_f := 11;
        ELSIF x =- 10628 THEN
            sigmoid_f := 11;
        ELSIF x =- 10627 THEN
            sigmoid_f := 11;
        ELSIF x =- 10626 THEN
            sigmoid_f := 11;
        ELSIF x =- 10625 THEN
            sigmoid_f := 11;
        ELSIF x =- 10624 THEN
            sigmoid_f := 11;
        ELSIF x =- 10623 THEN
            sigmoid_f := 11;
        ELSIF x =- 10622 THEN
            sigmoid_f := 11;
        ELSIF x =- 10621 THEN
            sigmoid_f := 11;
        ELSIF x =- 10620 THEN
            sigmoid_f := 11;
        ELSIF x =- 10619 THEN
            sigmoid_f := 11;
        ELSIF x =- 10618 THEN
            sigmoid_f := 11;
        ELSIF x =- 10617 THEN
            sigmoid_f := 11;
        ELSIF x =- 10616 THEN
            sigmoid_f := 11;
        ELSIF x =- 10615 THEN
            sigmoid_f := 11;
        ELSIF x =- 10614 THEN
            sigmoid_f := 11;
        ELSIF x =- 10613 THEN
            sigmoid_f := 11;
        ELSIF x =- 10612 THEN
            sigmoid_f := 11;
        ELSIF x =- 10611 THEN
            sigmoid_f := 11;
        ELSIF x =- 10610 THEN
            sigmoid_f := 11;
        ELSIF x =- 10609 THEN
            sigmoid_f := 11;
        ELSIF x =- 10608 THEN
            sigmoid_f := 11;
        ELSIF x =- 10607 THEN
            sigmoid_f := 11;
        ELSIF x =- 10606 THEN
            sigmoid_f := 11;
        ELSIF x =- 10605 THEN
            sigmoid_f := 11;
        ELSIF x =- 10604 THEN
            sigmoid_f := 11;
        ELSIF x =- 10603 THEN
            sigmoid_f := 11;
        ELSIF x =- 10602 THEN
            sigmoid_f := 11;
        ELSIF x =- 10601 THEN
            sigmoid_f := 11;
        ELSIF x =- 10600 THEN
            sigmoid_f := 11;
        ELSIF x =- 10599 THEN
            sigmoid_f := 11;
        ELSIF x =- 10598 THEN
            sigmoid_f := 11;
        ELSIF x =- 10597 THEN
            sigmoid_f := 11;
        ELSIF x =- 10596 THEN
            sigmoid_f := 11;
        ELSIF x =- 10595 THEN
            sigmoid_f := 11;
        ELSIF x =- 10594 THEN
            sigmoid_f := 11;
        ELSIF x =- 10593 THEN
            sigmoid_f := 11;
        ELSIF x =- 10592 THEN
            sigmoid_f := 11;
        ELSIF x =- 10591 THEN
            sigmoid_f := 11;
        ELSIF x =- 10590 THEN
            sigmoid_f := 11;
        ELSIF x =- 10589 THEN
            sigmoid_f := 11;
        ELSIF x =- 10588 THEN
            sigmoid_f := 11;
        ELSIF x =- 10587 THEN
            sigmoid_f := 11;
        ELSIF x =- 10586 THEN
            sigmoid_f := 11;
        ELSIF x =- 10585 THEN
            sigmoid_f := 11;
        ELSIF x =- 10584 THEN
            sigmoid_f := 11;
        ELSIF x =- 10583 THEN
            sigmoid_f := 11;
        ELSIF x =- 10582 THEN
            sigmoid_f := 11;
        ELSIF x =- 10581 THEN
            sigmoid_f := 11;
        ELSIF x =- 10580 THEN
            sigmoid_f := 11;
        ELSIF x =- 10579 THEN
            sigmoid_f := 11;
        ELSIF x =- 10578 THEN
            sigmoid_f := 11;
        ELSIF x =- 10577 THEN
            sigmoid_f := 11;
        ELSIF x =- 10576 THEN
            sigmoid_f := 11;
        ELSIF x =- 10575 THEN
            sigmoid_f := 11;
        ELSIF x =- 10574 THEN
            sigmoid_f := 11;
        ELSIF x =- 10573 THEN
            sigmoid_f := 11;
        ELSIF x =- 10572 THEN
            sigmoid_f := 11;
        ELSIF x =- 10571 THEN
            sigmoid_f := 11;
        ELSIF x =- 10570 THEN
            sigmoid_f := 11;
        ELSIF x =- 10569 THEN
            sigmoid_f := 11;
        ELSIF x =- 10568 THEN
            sigmoid_f := 11;
        ELSIF x =- 10567 THEN
            sigmoid_f := 11;
        ELSIF x =- 10566 THEN
            sigmoid_f := 11;
        ELSIF x =- 10565 THEN
            sigmoid_f := 11;
        ELSIF x =- 10564 THEN
            sigmoid_f := 11;
        ELSIF x =- 10563 THEN
            sigmoid_f := 11;
        ELSIF x =- 10562 THEN
            sigmoid_f := 11;
        ELSIF x =- 10561 THEN
            sigmoid_f := 11;
        ELSIF x =- 10560 THEN
            sigmoid_f := 11;
        ELSIF x =- 10559 THEN
            sigmoid_f := 11;
        ELSIF x =- 10558 THEN
            sigmoid_f := 11;
        ELSIF x =- 10557 THEN
            sigmoid_f := 11;
        ELSIF x =- 10556 THEN
            sigmoid_f := 11;
        ELSIF x =- 10555 THEN
            sigmoid_f := 11;
        ELSIF x =- 10554 THEN
            sigmoid_f := 11;
        ELSIF x =- 10553 THEN
            sigmoid_f := 11;
        ELSIF x =- 10552 THEN
            sigmoid_f := 11;
        ELSIF x =- 10551 THEN
            sigmoid_f := 11;
        ELSIF x =- 10550 THEN
            sigmoid_f := 11;
        ELSIF x =- 10549 THEN
            sigmoid_f := 11;
        ELSIF x =- 10548 THEN
            sigmoid_f := 11;
        ELSIF x =- 10547 THEN
            sigmoid_f := 11;
        ELSIF x =- 10546 THEN
            sigmoid_f := 11;
        ELSIF x =- 10545 THEN
            sigmoid_f := 11;
        ELSIF x =- 10544 THEN
            sigmoid_f := 11;
        ELSIF x =- 10543 THEN
            sigmoid_f := 11;
        ELSIF x =- 10542 THEN
            sigmoid_f := 11;
        ELSIF x =- 10541 THEN
            sigmoid_f := 11;
        ELSIF x =- 10540 THEN
            sigmoid_f := 11;
        ELSIF x =- 10539 THEN
            sigmoid_f := 11;
        ELSIF x =- 10538 THEN
            sigmoid_f := 11;
        ELSIF x =- 10537 THEN
            sigmoid_f := 11;
        ELSIF x =- 10536 THEN
            sigmoid_f := 11;
        ELSIF x =- 10535 THEN
            sigmoid_f := 11;
        ELSIF x =- 10534 THEN
            sigmoid_f := 11;
        ELSIF x =- 10533 THEN
            sigmoid_f := 11;
        ELSIF x =- 10532 THEN
            sigmoid_f := 12;
        ELSIF x =- 10531 THEN
            sigmoid_f := 12;
        ELSIF x =- 10530 THEN
            sigmoid_f := 12;
        ELSIF x =- 10529 THEN
            sigmoid_f := 12;
        ELSIF x =- 10528 THEN
            sigmoid_f := 12;
        ELSIF x =- 10527 THEN
            sigmoid_f := 12;
        ELSIF x =- 10526 THEN
            sigmoid_f := 12;
        ELSIF x =- 10525 THEN
            sigmoid_f := 12;
        ELSIF x =- 10524 THEN
            sigmoid_f := 12;
        ELSIF x =- 10523 THEN
            sigmoid_f := 12;
        ELSIF x =- 10522 THEN
            sigmoid_f := 12;
        ELSIF x =- 10521 THEN
            sigmoid_f := 12;
        ELSIF x =- 10520 THEN
            sigmoid_f := 12;
        ELSIF x =- 10519 THEN
            sigmoid_f := 12;
        ELSIF x =- 10518 THEN
            sigmoid_f := 12;
        ELSIF x =- 10517 THEN
            sigmoid_f := 12;
        ELSIF x =- 10516 THEN
            sigmoid_f := 12;
        ELSIF x =- 10515 THEN
            sigmoid_f := 12;
        ELSIF x =- 10514 THEN
            sigmoid_f := 12;
        ELSIF x =- 10513 THEN
            sigmoid_f := 12;
        ELSIF x =- 10512 THEN
            sigmoid_f := 12;
        ELSIF x =- 10511 THEN
            sigmoid_f := 12;
        ELSIF x =- 10510 THEN
            sigmoid_f := 12;
        ELSIF x =- 10509 THEN
            sigmoid_f := 12;
        ELSIF x =- 10508 THEN
            sigmoid_f := 12;
        ELSIF x =- 10507 THEN
            sigmoid_f := 12;
        ELSIF x =- 10506 THEN
            sigmoid_f := 12;
        ELSIF x =- 10505 THEN
            sigmoid_f := 12;
        ELSIF x =- 10504 THEN
            sigmoid_f := 12;
        ELSIF x =- 10503 THEN
            sigmoid_f := 12;
        ELSIF x =- 10502 THEN
            sigmoid_f := 12;
        ELSIF x =- 10501 THEN
            sigmoid_f := 12;
        ELSIF x =- 10500 THEN
            sigmoid_f := 12;
        ELSIF x =- 10499 THEN
            sigmoid_f := 12;
        ELSIF x =- 10498 THEN
            sigmoid_f := 12;
        ELSIF x =- 10497 THEN
            sigmoid_f := 12;
        ELSIF x =- 10496 THEN
            sigmoid_f := 12;
        ELSIF x =- 10495 THEN
            sigmoid_f := 12;
        ELSIF x =- 10494 THEN
            sigmoid_f := 12;
        ELSIF x =- 10493 THEN
            sigmoid_f := 12;
        ELSIF x =- 10492 THEN
            sigmoid_f := 12;
        ELSIF x =- 10491 THEN
            sigmoid_f := 12;
        ELSIF x =- 10490 THEN
            sigmoid_f := 12;
        ELSIF x =- 10489 THEN
            sigmoid_f := 12;
        ELSIF x =- 10488 THEN
            sigmoid_f := 12;
        ELSIF x =- 10487 THEN
            sigmoid_f := 12;
        ELSIF x =- 10486 THEN
            sigmoid_f := 12;
        ELSIF x =- 10485 THEN
            sigmoid_f := 12;
        ELSIF x =- 10484 THEN
            sigmoid_f := 12;
        ELSIF x =- 10483 THEN
            sigmoid_f := 12;
        ELSIF x =- 10482 THEN
            sigmoid_f := 12;
        ELSIF x =- 10481 THEN
            sigmoid_f := 12;
        ELSIF x =- 10480 THEN
            sigmoid_f := 12;
        ELSIF x =- 10479 THEN
            sigmoid_f := 12;
        ELSIF x =- 10478 THEN
            sigmoid_f := 12;
        ELSIF x =- 10477 THEN
            sigmoid_f := 12;
        ELSIF x =- 10476 THEN
            sigmoid_f := 12;
        ELSIF x =- 10475 THEN
            sigmoid_f := 12;
        ELSIF x =- 10474 THEN
            sigmoid_f := 12;
        ELSIF x =- 10473 THEN
            sigmoid_f := 12;
        ELSIF x =- 10472 THEN
            sigmoid_f := 12;
        ELSIF x =- 10471 THEN
            sigmoid_f := 12;
        ELSIF x =- 10470 THEN
            sigmoid_f := 12;
        ELSIF x =- 10469 THEN
            sigmoid_f := 12;
        ELSIF x =- 10468 THEN
            sigmoid_f := 12;
        ELSIF x =- 10467 THEN
            sigmoid_f := 12;
        ELSIF x =- 10466 THEN
            sigmoid_f := 12;
        ELSIF x =- 10465 THEN
            sigmoid_f := 12;
        ELSIF x =- 10464 THEN
            sigmoid_f := 12;
        ELSIF x =- 10463 THEN
            sigmoid_f := 12;
        ELSIF x =- 10462 THEN
            sigmoid_f := 12;
        ELSIF x =- 10461 THEN
            sigmoid_f := 12;
        ELSIF x =- 10460 THEN
            sigmoid_f := 12;
        ELSIF x =- 10459 THEN
            sigmoid_f := 12;
        ELSIF x =- 10458 THEN
            sigmoid_f := 12;
        ELSIF x =- 10457 THEN
            sigmoid_f := 12;
        ELSIF x =- 10456 THEN
            sigmoid_f := 12;
        ELSIF x =- 10455 THEN
            sigmoid_f := 12;
        ELSIF x =- 10454 THEN
            sigmoid_f := 12;
        ELSIF x =- 10453 THEN
            sigmoid_f := 12;
        ELSIF x =- 10452 THEN
            sigmoid_f := 12;
        ELSIF x =- 10451 THEN
            sigmoid_f := 12;
        ELSIF x =- 10450 THEN
            sigmoid_f := 12;
        ELSIF x =- 10449 THEN
            sigmoid_f := 12;
        ELSIF x =- 10448 THEN
            sigmoid_f := 12;
        ELSIF x =- 10447 THEN
            sigmoid_f := 12;
        ELSIF x =- 10446 THEN
            sigmoid_f := 12;
        ELSIF x =- 10445 THEN
            sigmoid_f := 12;
        ELSIF x =- 10444 THEN
            sigmoid_f := 12;
        ELSIF x =- 10443 THEN
            sigmoid_f := 12;
        ELSIF x =- 10442 THEN
            sigmoid_f := 12;
        ELSIF x =- 10441 THEN
            sigmoid_f := 12;
        ELSIF x =- 10440 THEN
            sigmoid_f := 12;
        ELSIF x =- 10439 THEN
            sigmoid_f := 12;
        ELSIF x =- 10438 THEN
            sigmoid_f := 12;
        ELSIF x =- 10437 THEN
            sigmoid_f := 12;
        ELSIF x =- 10436 THEN
            sigmoid_f := 12;
        ELSIF x =- 10435 THEN
            sigmoid_f := 12;
        ELSIF x =- 10434 THEN
            sigmoid_f := 12;
        ELSIF x =- 10433 THEN
            sigmoid_f := 12;
        ELSIF x =- 10432 THEN
            sigmoid_f := 12;
        ELSIF x =- 10431 THEN
            sigmoid_f := 12;
        ELSIF x =- 10430 THEN
            sigmoid_f := 12;
        ELSIF x =- 10429 THEN
            sigmoid_f := 12;
        ELSIF x =- 10428 THEN
            sigmoid_f := 12;
        ELSIF x =- 10427 THEN
            sigmoid_f := 12;
        ELSIF x =- 10426 THEN
            sigmoid_f := 12;
        ELSIF x =- 10425 THEN
            sigmoid_f := 12;
        ELSIF x =- 10424 THEN
            sigmoid_f := 12;
        ELSIF x =- 10423 THEN
            sigmoid_f := 12;
        ELSIF x =- 10422 THEN
            sigmoid_f := 12;
        ELSIF x =- 10421 THEN
            sigmoid_f := 12;
        ELSIF x =- 10420 THEN
            sigmoid_f := 12;
        ELSIF x =- 10419 THEN
            sigmoid_f := 12;
        ELSIF x =- 10418 THEN
            sigmoid_f := 12;
        ELSIF x =- 10417 THEN
            sigmoid_f := 12;
        ELSIF x =- 10416 THEN
            sigmoid_f := 12;
        ELSIF x =- 10415 THEN
            sigmoid_f := 12;
        ELSIF x =- 10414 THEN
            sigmoid_f := 12;
        ELSIF x =- 10413 THEN
            sigmoid_f := 12;
        ELSIF x =- 10412 THEN
            sigmoid_f := 12;
        ELSIF x =- 10411 THEN
            sigmoid_f := 12;
        ELSIF x =- 10410 THEN
            sigmoid_f := 12;
        ELSIF x =- 10409 THEN
            sigmoid_f := 12;
        ELSIF x =- 10408 THEN
            sigmoid_f := 12;
        ELSIF x =- 10407 THEN
            sigmoid_f := 12;
        ELSIF x =- 10406 THEN
            sigmoid_f := 12;
        ELSIF x =- 10405 THEN
            sigmoid_f := 12;
        ELSIF x =- 10404 THEN
            sigmoid_f := 12;
        ELSIF x =- 10403 THEN
            sigmoid_f := 12;
        ELSIF x =- 10402 THEN
            sigmoid_f := 12;
        ELSIF x =- 10401 THEN
            sigmoid_f := 12;
        ELSIF x =- 10400 THEN
            sigmoid_f := 12;
        ELSIF x =- 10399 THEN
            sigmoid_f := 12;
        ELSIF x =- 10398 THEN
            sigmoid_f := 12;
        ELSIF x =- 10397 THEN
            sigmoid_f := 12;
        ELSIF x =- 10396 THEN
            sigmoid_f := 12;
        ELSIF x =- 10395 THEN
            sigmoid_f := 12;
        ELSIF x =- 10394 THEN
            sigmoid_f := 12;
        ELSIF x =- 10393 THEN
            sigmoid_f := 12;
        ELSIF x =- 10392 THEN
            sigmoid_f := 12;
        ELSIF x =- 10391 THEN
            sigmoid_f := 12;
        ELSIF x =- 10390 THEN
            sigmoid_f := 12;
        ELSIF x =- 10389 THEN
            sigmoid_f := 12;
        ELSIF x =- 10388 THEN
            sigmoid_f := 12;
        ELSIF x =- 10387 THEN
            sigmoid_f := 12;
        ELSIF x =- 10386 THEN
            sigmoid_f := 13;
        ELSIF x =- 10385 THEN
            sigmoid_f := 13;
        ELSIF x =- 10384 THEN
            sigmoid_f := 13;
        ELSIF x =- 10383 THEN
            sigmoid_f := 13;
        ELSIF x =- 10382 THEN
            sigmoid_f := 13;
        ELSIF x =- 10381 THEN
            sigmoid_f := 13;
        ELSIF x =- 10380 THEN
            sigmoid_f := 13;
        ELSIF x =- 10379 THEN
            sigmoid_f := 13;
        ELSIF x =- 10378 THEN
            sigmoid_f := 13;
        ELSIF x =- 10377 THEN
            sigmoid_f := 13;
        ELSIF x =- 10376 THEN
            sigmoid_f := 13;
        ELSIF x =- 10375 THEN
            sigmoid_f := 13;
        ELSIF x =- 10374 THEN
            sigmoid_f := 13;
        ELSIF x =- 10373 THEN
            sigmoid_f := 13;
        ELSIF x =- 10372 THEN
            sigmoid_f := 13;
        ELSIF x =- 10371 THEN
            sigmoid_f := 13;
        ELSIF x =- 10370 THEN
            sigmoid_f := 13;
        ELSIF x =- 10369 THEN
            sigmoid_f := 13;
        ELSIF x =- 10368 THEN
            sigmoid_f := 13;
        ELSIF x =- 10367 THEN
            sigmoid_f := 13;
        ELSIF x =- 10366 THEN
            sigmoid_f := 13;
        ELSIF x =- 10365 THEN
            sigmoid_f := 13;
        ELSIF x =- 10364 THEN
            sigmoid_f := 13;
        ELSIF x =- 10363 THEN
            sigmoid_f := 13;
        ELSIF x =- 10362 THEN
            sigmoid_f := 13;
        ELSIF x =- 10361 THEN
            sigmoid_f := 13;
        ELSIF x =- 10360 THEN
            sigmoid_f := 13;
        ELSIF x =- 10359 THEN
            sigmoid_f := 13;
        ELSIF x =- 10358 THEN
            sigmoid_f := 13;
        ELSIF x =- 10357 THEN
            sigmoid_f := 13;
        ELSIF x =- 10356 THEN
            sigmoid_f := 13;
        ELSIF x =- 10355 THEN
            sigmoid_f := 13;
        ELSIF x =- 10354 THEN
            sigmoid_f := 13;
        ELSIF x =- 10353 THEN
            sigmoid_f := 13;
        ELSIF x =- 10352 THEN
            sigmoid_f := 13;
        ELSIF x =- 10351 THEN
            sigmoid_f := 13;
        ELSIF x =- 10350 THEN
            sigmoid_f := 13;
        ELSIF x =- 10349 THEN
            sigmoid_f := 13;
        ELSIF x =- 10348 THEN
            sigmoid_f := 13;
        ELSIF x =- 10347 THEN
            sigmoid_f := 13;
        ELSIF x =- 10346 THEN
            sigmoid_f := 13;
        ELSIF x =- 10345 THEN
            sigmoid_f := 13;
        ELSIF x =- 10344 THEN
            sigmoid_f := 13;
        ELSIF x =- 10343 THEN
            sigmoid_f := 13;
        ELSIF x =- 10342 THEN
            sigmoid_f := 13;
        ELSIF x =- 10341 THEN
            sigmoid_f := 13;
        ELSIF x =- 10340 THEN
            sigmoid_f := 13;
        ELSIF x =- 10339 THEN
            sigmoid_f := 13;
        ELSIF x =- 10338 THEN
            sigmoid_f := 13;
        ELSIF x =- 10337 THEN
            sigmoid_f := 13;
        ELSIF x =- 10336 THEN
            sigmoid_f := 13;
        ELSIF x =- 10335 THEN
            sigmoid_f := 13;
        ELSIF x =- 10334 THEN
            sigmoid_f := 13;
        ELSIF x =- 10333 THEN
            sigmoid_f := 13;
        ELSIF x =- 10332 THEN
            sigmoid_f := 13;
        ELSIF x =- 10331 THEN
            sigmoid_f := 13;
        ELSIF x =- 10330 THEN
            sigmoid_f := 13;
        ELSIF x =- 10329 THEN
            sigmoid_f := 13;
        ELSIF x =- 10328 THEN
            sigmoid_f := 13;
        ELSIF x =- 10327 THEN
            sigmoid_f := 13;
        ELSIF x =- 10326 THEN
            sigmoid_f := 13;
        ELSIF x =- 10325 THEN
            sigmoid_f := 13;
        ELSIF x =- 10324 THEN
            sigmoid_f := 13;
        ELSIF x =- 10323 THEN
            sigmoid_f := 13;
        ELSIF x =- 10322 THEN
            sigmoid_f := 13;
        ELSIF x =- 10321 THEN
            sigmoid_f := 13;
        ELSIF x =- 10320 THEN
            sigmoid_f := 13;
        ELSIF x =- 10319 THEN
            sigmoid_f := 13;
        ELSIF x =- 10318 THEN
            sigmoid_f := 13;
        ELSIF x =- 10317 THEN
            sigmoid_f := 13;
        ELSIF x =- 10316 THEN
            sigmoid_f := 13;
        ELSIF x =- 10315 THEN
            sigmoid_f := 13;
        ELSIF x =- 10314 THEN
            sigmoid_f := 13;
        ELSIF x =- 10313 THEN
            sigmoid_f := 13;
        ELSIF x =- 10312 THEN
            sigmoid_f := 13;
        ELSIF x =- 10311 THEN
            sigmoid_f := 13;
        ELSIF x =- 10310 THEN
            sigmoid_f := 13;
        ELSIF x =- 10309 THEN
            sigmoid_f := 13;
        ELSIF x =- 10308 THEN
            sigmoid_f := 13;
        ELSIF x =- 10307 THEN
            sigmoid_f := 13;
        ELSIF x =- 10306 THEN
            sigmoid_f := 13;
        ELSIF x =- 10305 THEN
            sigmoid_f := 13;
        ELSIF x =- 10304 THEN
            sigmoid_f := 13;
        ELSIF x =- 10303 THEN
            sigmoid_f := 13;
        ELSIF x =- 10302 THEN
            sigmoid_f := 13;
        ELSIF x =- 10301 THEN
            sigmoid_f := 13;
        ELSIF x =- 10300 THEN
            sigmoid_f := 13;
        ELSIF x =- 10299 THEN
            sigmoid_f := 13;
        ELSIF x =- 10298 THEN
            sigmoid_f := 13;
        ELSIF x =- 10297 THEN
            sigmoid_f := 13;
        ELSIF x =- 10296 THEN
            sigmoid_f := 13;
        ELSIF x =- 10295 THEN
            sigmoid_f := 13;
        ELSIF x =- 10294 THEN
            sigmoid_f := 13;
        ELSIF x =- 10293 THEN
            sigmoid_f := 13;
        ELSIF x =- 10292 THEN
            sigmoid_f := 13;
        ELSIF x =- 10291 THEN
            sigmoid_f := 13;
        ELSIF x =- 10290 THEN
            sigmoid_f := 13;
        ELSIF x =- 10289 THEN
            sigmoid_f := 13;
        ELSIF x =- 10288 THEN
            sigmoid_f := 13;
        ELSIF x =- 10287 THEN
            sigmoid_f := 13;
        ELSIF x =- 10286 THEN
            sigmoid_f := 13;
        ELSIF x =- 10285 THEN
            sigmoid_f := 13;
        ELSIF x =- 10284 THEN
            sigmoid_f := 13;
        ELSIF x =- 10283 THEN
            sigmoid_f := 13;
        ELSIF x =- 10282 THEN
            sigmoid_f := 13;
        ELSIF x =- 10281 THEN
            sigmoid_f := 13;
        ELSIF x =- 10280 THEN
            sigmoid_f := 13;
        ELSIF x =- 10279 THEN
            sigmoid_f := 13;
        ELSIF x =- 10278 THEN
            sigmoid_f := 13;
        ELSIF x =- 10277 THEN
            sigmoid_f := 13;
        ELSIF x =- 10276 THEN
            sigmoid_f := 13;
        ELSIF x =- 10275 THEN
            sigmoid_f := 13;
        ELSIF x =- 10274 THEN
            sigmoid_f := 13;
        ELSIF x =- 10273 THEN
            sigmoid_f := 13;
        ELSIF x =- 10272 THEN
            sigmoid_f := 13;
        ELSIF x =- 10271 THEN
            sigmoid_f := 13;
        ELSIF x =- 10270 THEN
            sigmoid_f := 13;
        ELSIF x =- 10269 THEN
            sigmoid_f := 13;
        ELSIF x =- 10268 THEN
            sigmoid_f := 13;
        ELSIF x =- 10267 THEN
            sigmoid_f := 13;
        ELSIF x =- 10266 THEN
            sigmoid_f := 13;
        ELSIF x =- 10265 THEN
            sigmoid_f := 13;
        ELSIF x =- 10264 THEN
            sigmoid_f := 13;
        ELSIF x =- 10263 THEN
            sigmoid_f := 13;
        ELSIF x =- 10262 THEN
            sigmoid_f := 13;
        ELSIF x =- 10261 THEN
            sigmoid_f := 13;
        ELSIF x =- 10260 THEN
            sigmoid_f := 13;
        ELSIF x =- 10259 THEN
            sigmoid_f := 13;
        ELSIF x =- 10258 THEN
            sigmoid_f := 13;
        ELSIF x =- 10257 THEN
            sigmoid_f := 13;
        ELSIF x =- 10256 THEN
            sigmoid_f := 13;
        ELSIF x =- 10255 THEN
            sigmoid_f := 13;
        ELSIF x =- 10254 THEN
            sigmoid_f := 13;
        ELSIF x =- 10253 THEN
            sigmoid_f := 13;
        ELSIF x =- 10252 THEN
            sigmoid_f := 13;
        ELSIF x =- 10251 THEN
            sigmoid_f := 13;
        ELSIF x =- 10250 THEN
            sigmoid_f := 13;
        ELSIF x =- 10249 THEN
            sigmoid_f := 13;
        ELSIF x =- 10248 THEN
            sigmoid_f := 13;
        ELSIF x =- 10247 THEN
            sigmoid_f := 13;
        ELSIF x =- 10246 THEN
            sigmoid_f := 13;
        ELSIF x =- 10245 THEN
            sigmoid_f := 13;
        ELSIF x =- 10244 THEN
            sigmoid_f := 13;
        ELSIF x =- 10243 THEN
            sigmoid_f := 13;
        ELSIF x =- 10242 THEN
            sigmoid_f := 13;
        ELSIF x =- 10241 THEN
            sigmoid_f := 13;
        ELSIF x =- 10240 THEN
            sigmoid_f := 14;
        ELSIF x =- 10239 THEN
            sigmoid_f := 14;
        ELSIF x =- 10238 THEN
            sigmoid_f := 14;
        ELSIF x =- 10237 THEN
            sigmoid_f := 14;
        ELSIF x =- 10236 THEN
            sigmoid_f := 14;
        ELSIF x =- 10235 THEN
            sigmoid_f := 14;
        ELSIF x =- 10234 THEN
            sigmoid_f := 14;
        ELSIF x =- 10233 THEN
            sigmoid_f := 14;
        ELSIF x =- 10232 THEN
            sigmoid_f := 14;
        ELSIF x =- 10231 THEN
            sigmoid_f := 14;
        ELSIF x =- 10230 THEN
            sigmoid_f := 14;
        ELSIF x =- 10229 THEN
            sigmoid_f := 14;
        ELSIF x =- 10228 THEN
            sigmoid_f := 14;
        ELSIF x =- 10227 THEN
            sigmoid_f := 14;
        ELSIF x =- 10226 THEN
            sigmoid_f := 14;
        ELSIF x =- 10225 THEN
            sigmoid_f := 14;
        ELSIF x =- 10224 THEN
            sigmoid_f := 14;
        ELSIF x =- 10223 THEN
            sigmoid_f := 14;
        ELSIF x =- 10222 THEN
            sigmoid_f := 14;
        ELSIF x =- 10221 THEN
            sigmoid_f := 14;
        ELSIF x =- 10220 THEN
            sigmoid_f := 14;
        ELSIF x =- 10219 THEN
            sigmoid_f := 14;
        ELSIF x =- 10218 THEN
            sigmoid_f := 14;
        ELSIF x =- 10217 THEN
            sigmoid_f := 14;
        ELSIF x =- 10216 THEN
            sigmoid_f := 14;
        ELSIF x =- 10215 THEN
            sigmoid_f := 14;
        ELSIF x =- 10214 THEN
            sigmoid_f := 14;
        ELSIF x =- 10213 THEN
            sigmoid_f := 14;
        ELSIF x =- 10212 THEN
            sigmoid_f := 14;
        ELSIF x =- 10211 THEN
            sigmoid_f := 14;
        ELSIF x =- 10210 THEN
            sigmoid_f := 14;
        ELSIF x =- 10209 THEN
            sigmoid_f := 14;
        ELSIF x =- 10208 THEN
            sigmoid_f := 14;
        ELSIF x =- 10207 THEN
            sigmoid_f := 14;
        ELSIF x =- 10206 THEN
            sigmoid_f := 14;
        ELSIF x =- 10205 THEN
            sigmoid_f := 14;
        ELSIF x =- 10204 THEN
            sigmoid_f := 14;
        ELSIF x =- 10203 THEN
            sigmoid_f := 14;
        ELSIF x =- 10202 THEN
            sigmoid_f := 14;
        ELSIF x =- 10201 THEN
            sigmoid_f := 14;
        ELSIF x =- 10200 THEN
            sigmoid_f := 14;
        ELSIF x =- 10199 THEN
            sigmoid_f := 14;
        ELSIF x =- 10198 THEN
            sigmoid_f := 14;
        ELSIF x =- 10197 THEN
            sigmoid_f := 14;
        ELSIF x =- 10196 THEN
            sigmoid_f := 14;
        ELSIF x =- 10195 THEN
            sigmoid_f := 14;
        ELSIF x =- 10194 THEN
            sigmoid_f := 14;
        ELSIF x =- 10193 THEN
            sigmoid_f := 14;
        ELSIF x =- 10192 THEN
            sigmoid_f := 14;
        ELSIF x =- 10191 THEN
            sigmoid_f := 14;
        ELSIF x =- 10190 THEN
            sigmoid_f := 14;
        ELSIF x =- 10189 THEN
            sigmoid_f := 14;
        ELSIF x =- 10188 THEN
            sigmoid_f := 14;
        ELSIF x =- 10187 THEN
            sigmoid_f := 14;
        ELSIF x =- 10186 THEN
            sigmoid_f := 14;
        ELSIF x =- 10185 THEN
            sigmoid_f := 14;
        ELSIF x =- 10184 THEN
            sigmoid_f := 14;
        ELSIF x =- 10183 THEN
            sigmoid_f := 14;
        ELSIF x =- 10182 THEN
            sigmoid_f := 14;
        ELSIF x =- 10181 THEN
            sigmoid_f := 14;
        ELSIF x =- 10180 THEN
            sigmoid_f := 14;
        ELSIF x =- 10179 THEN
            sigmoid_f := 14;
        ELSIF x =- 10178 THEN
            sigmoid_f := 14;
        ELSIF x =- 10177 THEN
            sigmoid_f := 14;
        ELSIF x =- 10176 THEN
            sigmoid_f := 14;
        ELSIF x =- 10175 THEN
            sigmoid_f := 14;
        ELSIF x =- 10174 THEN
            sigmoid_f := 14;
        ELSIF x =- 10173 THEN
            sigmoid_f := 14;
        ELSIF x =- 10172 THEN
            sigmoid_f := 14;
        ELSIF x =- 10171 THEN
            sigmoid_f := 14;
        ELSIF x =- 10170 THEN
            sigmoid_f := 14;
        ELSIF x =- 10169 THEN
            sigmoid_f := 14;
        ELSIF x =- 10168 THEN
            sigmoid_f := 14;
        ELSIF x =- 10167 THEN
            sigmoid_f := 14;
        ELSIF x =- 10166 THEN
            sigmoid_f := 14;
        ELSIF x =- 10165 THEN
            sigmoid_f := 14;
        ELSIF x =- 10164 THEN
            sigmoid_f := 14;
        ELSIF x =- 10163 THEN
            sigmoid_f := 14;
        ELSIF x =- 10162 THEN
            sigmoid_f := 14;
        ELSIF x =- 10161 THEN
            sigmoid_f := 14;
        ELSIF x =- 10160 THEN
            sigmoid_f := 14;
        ELSIF x =- 10159 THEN
            sigmoid_f := 14;
        ELSIF x =- 10158 THEN
            sigmoid_f := 14;
        ELSIF x =- 10157 THEN
            sigmoid_f := 14;
        ELSIF x =- 10156 THEN
            sigmoid_f := 14;
        ELSIF x =- 10155 THEN
            sigmoid_f := 14;
        ELSIF x =- 10154 THEN
            sigmoid_f := 14;
        ELSIF x =- 10153 THEN
            sigmoid_f := 14;
        ELSIF x =- 10152 THEN
            sigmoid_f := 14;
        ELSIF x =- 10151 THEN
            sigmoid_f := 14;
        ELSIF x =- 10150 THEN
            sigmoid_f := 14;
        ELSIF x =- 10149 THEN
            sigmoid_f := 14;
        ELSIF x =- 10148 THEN
            sigmoid_f := 14;
        ELSIF x =- 10147 THEN
            sigmoid_f := 14;
        ELSIF x =- 10146 THEN
            sigmoid_f := 14;
        ELSIF x =- 10145 THEN
            sigmoid_f := 14;
        ELSIF x =- 10144 THEN
            sigmoid_f := 14;
        ELSIF x =- 10143 THEN
            sigmoid_f := 14;
        ELSIF x =- 10142 THEN
            sigmoid_f := 14;
        ELSIF x =- 10141 THEN
            sigmoid_f := 14;
        ELSIF x =- 10140 THEN
            sigmoid_f := 14;
        ELSIF x =- 10139 THEN
            sigmoid_f := 14;
        ELSIF x =- 10138 THEN
            sigmoid_f := 14;
        ELSIF x =- 10137 THEN
            sigmoid_f := 14;
        ELSIF x =- 10136 THEN
            sigmoid_f := 14;
        ELSIF x =- 10135 THEN
            sigmoid_f := 14;
        ELSIF x =- 10134 THEN
            sigmoid_f := 14;
        ELSIF x =- 10133 THEN
            sigmoid_f := 14;
        ELSIF x =- 10132 THEN
            sigmoid_f := 14;
        ELSIF x =- 10131 THEN
            sigmoid_f := 14;
        ELSIF x =- 10130 THEN
            sigmoid_f := 14;
        ELSIF x =- 10129 THEN
            sigmoid_f := 14;
        ELSIF x =- 10128 THEN
            sigmoid_f := 14;
        ELSIF x =- 10127 THEN
            sigmoid_f := 14;
        ELSIF x =- 10126 THEN
            sigmoid_f := 14;
        ELSIF x =- 10125 THEN
            sigmoid_f := 14;
        ELSIF x =- 10124 THEN
            sigmoid_f := 14;
        ELSIF x =- 10123 THEN
            sigmoid_f := 14;
        ELSIF x =- 10122 THEN
            sigmoid_f := 14;
        ELSIF x =- 10121 THEN
            sigmoid_f := 14;
        ELSIF x =- 10120 THEN
            sigmoid_f := 14;
        ELSIF x =- 10119 THEN
            sigmoid_f := 14;
        ELSIF x =- 10118 THEN
            sigmoid_f := 14;
        ELSIF x =- 10117 THEN
            sigmoid_f := 14;
        ELSIF x =- 10116 THEN
            sigmoid_f := 14;
        ELSIF x =- 10115 THEN
            sigmoid_f := 14;
        ELSIF x =- 10114 THEN
            sigmoid_f := 14;
        ELSIF x =- 10113 THEN
            sigmoid_f := 14;
        ELSIF x =- 10112 THEN
            sigmoid_f := 14;
        ELSIF x =- 10111 THEN
            sigmoid_f := 14;
        ELSIF x =- 10110 THEN
            sigmoid_f := 14;
        ELSIF x =- 10109 THEN
            sigmoid_f := 14;
        ELSIF x =- 10108 THEN
            sigmoid_f := 14;
        ELSIF x =- 10107 THEN
            sigmoid_f := 14;
        ELSIF x =- 10106 THEN
            sigmoid_f := 14;
        ELSIF x =- 10105 THEN
            sigmoid_f := 14;
        ELSIF x =- 10104 THEN
            sigmoid_f := 14;
        ELSIF x =- 10103 THEN
            sigmoid_f := 14;
        ELSIF x =- 10102 THEN
            sigmoid_f := 14;
        ELSIF x =- 10101 THEN
            sigmoid_f := 14;
        ELSIF x =- 10100 THEN
            sigmoid_f := 14;
        ELSIF x =- 10099 THEN
            sigmoid_f := 14;
        ELSIF x =- 10098 THEN
            sigmoid_f := 14;
        ELSIF x =- 10097 THEN
            sigmoid_f := 14;
        ELSIF x =- 10096 THEN
            sigmoid_f := 14;
        ELSIF x =- 10095 THEN
            sigmoid_f := 14;
        ELSIF x =- 10094 THEN
            sigmoid_f := 14;
        ELSIF x =- 10093 THEN
            sigmoid_f := 14;
        ELSIF x =- 10092 THEN
            sigmoid_f := 14;
        ELSIF x =- 10091 THEN
            sigmoid_f := 14;
        ELSIF x =- 10090 THEN
            sigmoid_f := 14;
        ELSIF x =- 10089 THEN
            sigmoid_f := 14;
        ELSIF x =- 10088 THEN
            sigmoid_f := 14;
        ELSIF x =- 10087 THEN
            sigmoid_f := 14;
        ELSIF x =- 10086 THEN
            sigmoid_f := 14;
        ELSIF x =- 10085 THEN
            sigmoid_f := 14;
        ELSIF x =- 10084 THEN
            sigmoid_f := 14;
        ELSIF x =- 10083 THEN
            sigmoid_f := 14;
        ELSIF x =- 10082 THEN
            sigmoid_f := 15;
        ELSIF x =- 10081 THEN
            sigmoid_f := 15;
        ELSIF x =- 10080 THEN
            sigmoid_f := 15;
        ELSIF x =- 10079 THEN
            sigmoid_f := 15;
        ELSIF x =- 10078 THEN
            sigmoid_f := 15;
        ELSIF x =- 10077 THEN
            sigmoid_f := 15;
        ELSIF x =- 10076 THEN
            sigmoid_f := 15;
        ELSIF x =- 10075 THEN
            sigmoid_f := 15;
        ELSIF x =- 10074 THEN
            sigmoid_f := 15;
        ELSIF x =- 10073 THEN
            sigmoid_f := 15;
        ELSIF x =- 10072 THEN
            sigmoid_f := 15;
        ELSIF x =- 10071 THEN
            sigmoid_f := 15;
        ELSIF x =- 10070 THEN
            sigmoid_f := 15;
        ELSIF x =- 10069 THEN
            sigmoid_f := 15;
        ELSIF x =- 10068 THEN
            sigmoid_f := 15;
        ELSIF x =- 10067 THEN
            sigmoid_f := 15;
        ELSIF x =- 10066 THEN
            sigmoid_f := 15;
        ELSIF x =- 10065 THEN
            sigmoid_f := 15;
        ELSIF x =- 10064 THEN
            sigmoid_f := 15;
        ELSIF x =- 10063 THEN
            sigmoid_f := 15;
        ELSIF x =- 10062 THEN
            sigmoid_f := 15;
        ELSIF x =- 10061 THEN
            sigmoid_f := 15;
        ELSIF x =- 10060 THEN
            sigmoid_f := 15;
        ELSIF x =- 10059 THEN
            sigmoid_f := 15;
        ELSIF x =- 10058 THEN
            sigmoid_f := 15;
        ELSIF x =- 10057 THEN
            sigmoid_f := 15;
        ELSIF x =- 10056 THEN
            sigmoid_f := 15;
        ELSIF x =- 10055 THEN
            sigmoid_f := 15;
        ELSIF x =- 10054 THEN
            sigmoid_f := 15;
        ELSIF x =- 10053 THEN
            sigmoid_f := 15;
        ELSIF x =- 10052 THEN
            sigmoid_f := 15;
        ELSIF x =- 10051 THEN
            sigmoid_f := 15;
        ELSIF x =- 10050 THEN
            sigmoid_f := 15;
        ELSIF x =- 10049 THEN
            sigmoid_f := 15;
        ELSIF x =- 10048 THEN
            sigmoid_f := 15;
        ELSIF x =- 10047 THEN
            sigmoid_f := 15;
        ELSIF x =- 10046 THEN
            sigmoid_f := 15;
        ELSIF x =- 10045 THEN
            sigmoid_f := 15;
        ELSIF x =- 10044 THEN
            sigmoid_f := 15;
        ELSIF x =- 10043 THEN
            sigmoid_f := 15;
        ELSIF x =- 10042 THEN
            sigmoid_f := 15;
        ELSIF x =- 10041 THEN
            sigmoid_f := 15;
        ELSIF x =- 10040 THEN
            sigmoid_f := 15;
        ELSIF x =- 10039 THEN
            sigmoid_f := 15;
        ELSIF x =- 10038 THEN
            sigmoid_f := 15;
        ELSIF x =- 10037 THEN
            sigmoid_f := 15;
        ELSIF x =- 10036 THEN
            sigmoid_f := 15;
        ELSIF x =- 10035 THEN
            sigmoid_f := 15;
        ELSIF x =- 10034 THEN
            sigmoid_f := 15;
        ELSIF x =- 10033 THEN
            sigmoid_f := 15;
        ELSIF x =- 10032 THEN
            sigmoid_f := 15;
        ELSIF x =- 10031 THEN
            sigmoid_f := 15;
        ELSIF x =- 10030 THEN
            sigmoid_f := 15;
        ELSIF x =- 10029 THEN
            sigmoid_f := 15;
        ELSIF x =- 10028 THEN
            sigmoid_f := 15;
        ELSIF x =- 10027 THEN
            sigmoid_f := 15;
        ELSIF x =- 10026 THEN
            sigmoid_f := 15;
        ELSIF x =- 10025 THEN
            sigmoid_f := 15;
        ELSIF x =- 10024 THEN
            sigmoid_f := 15;
        ELSIF x =- 10023 THEN
            sigmoid_f := 15;
        ELSIF x =- 10022 THEN
            sigmoid_f := 15;
        ELSIF x =- 10021 THEN
            sigmoid_f := 15;
        ELSIF x =- 10020 THEN
            sigmoid_f := 15;
        ELSIF x =- 10019 THEN
            sigmoid_f := 15;
        ELSIF x =- 10018 THEN
            sigmoid_f := 15;
        ELSIF x =- 10017 THEN
            sigmoid_f := 15;
        ELSIF x =- 10016 THEN
            sigmoid_f := 15;
        ELSIF x =- 10015 THEN
            sigmoid_f := 15;
        ELSIF x =- 10014 THEN
            sigmoid_f := 15;
        ELSIF x =- 10013 THEN
            sigmoid_f := 15;
        ELSIF x =- 10012 THEN
            sigmoid_f := 15;
        ELSIF x =- 10011 THEN
            sigmoid_f := 15;
        ELSIF x =- 10010 THEN
            sigmoid_f := 15;
        ELSIF x =- 10009 THEN
            sigmoid_f := 15;
        ELSIF x =- 10008 THEN
            sigmoid_f := 15;
        ELSIF x =- 10007 THEN
            sigmoid_f := 15;
        ELSIF x =- 10006 THEN
            sigmoid_f := 15;
        ELSIF x =- 10005 THEN
            sigmoid_f := 15;
        ELSIF x =- 10004 THEN
            sigmoid_f := 15;
        ELSIF x =- 10003 THEN
            sigmoid_f := 15;
        ELSIF x =- 10002 THEN
            sigmoid_f := 15;
        ELSIF x =- 10001 THEN
            sigmoid_f := 15;
        ELSIF x =- 10000 THEN
            sigmoid_f := 15;
        ELSIF x =- 9999 THEN
            sigmoid_f := 15;
        ELSIF x =- 9998 THEN
            sigmoid_f := 15;
        ELSIF x =- 9997 THEN
            sigmoid_f := 15;
        ELSIF x =- 9996 THEN
            sigmoid_f := 15;
        ELSIF x =- 9995 THEN
            sigmoid_f := 15;
        ELSIF x =- 9994 THEN
            sigmoid_f := 15;
        ELSIF x =- 9993 THEN
            sigmoid_f := 15;
        ELSIF x =- 9992 THEN
            sigmoid_f := 15;
        ELSIF x =- 9991 THEN
            sigmoid_f := 15;
        ELSIF x =- 9990 THEN
            sigmoid_f := 15;
        ELSIF x =- 9989 THEN
            sigmoid_f := 15;
        ELSIF x =- 9988 THEN
            sigmoid_f := 15;
        ELSIF x =- 9987 THEN
            sigmoid_f := 15;
        ELSIF x =- 9986 THEN
            sigmoid_f := 15;
        ELSIF x =- 9985 THEN
            sigmoid_f := 15;
        ELSIF x =- 9984 THEN
            sigmoid_f := 15;
        ELSIF x =- 9983 THEN
            sigmoid_f := 15;
        ELSIF x =- 9982 THEN
            sigmoid_f := 15;
        ELSIF x =- 9981 THEN
            sigmoid_f := 15;
        ELSIF x =- 9980 THEN
            sigmoid_f := 15;
        ELSIF x =- 9979 THEN
            sigmoid_f := 15;
        ELSIF x =- 9978 THEN
            sigmoid_f := 15;
        ELSIF x =- 9977 THEN
            sigmoid_f := 15;
        ELSIF x =- 9976 THEN
            sigmoid_f := 15;
        ELSIF x =- 9975 THEN
            sigmoid_f := 15;
        ELSIF x =- 9974 THEN
            sigmoid_f := 15;
        ELSIF x =- 9973 THEN
            sigmoid_f := 15;
        ELSIF x =- 9972 THEN
            sigmoid_f := 15;
        ELSIF x =- 9971 THEN
            sigmoid_f := 15;
        ELSIF x =- 9970 THEN
            sigmoid_f := 15;
        ELSIF x =- 9969 THEN
            sigmoid_f := 15;
        ELSIF x =- 9968 THEN
            sigmoid_f := 15;
        ELSIF x =- 9967 THEN
            sigmoid_f := 15;
        ELSIF x =- 9966 THEN
            sigmoid_f := 15;
        ELSIF x =- 9965 THEN
            sigmoid_f := 15;
        ELSIF x =- 9964 THEN
            sigmoid_f := 15;
        ELSIF x =- 9963 THEN
            sigmoid_f := 15;
        ELSIF x =- 9962 THEN
            sigmoid_f := 15;
        ELSIF x =- 9961 THEN
            sigmoid_f := 15;
        ELSIF x =- 9960 THEN
            sigmoid_f := 15;
        ELSIF x =- 9959 THEN
            sigmoid_f := 15;
        ELSIF x =- 9958 THEN
            sigmoid_f := 15;
        ELSIF x =- 9957 THEN
            sigmoid_f := 15;
        ELSIF x =- 9956 THEN
            sigmoid_f := 15;
        ELSIF x =- 9955 THEN
            sigmoid_f := 15;
        ELSIF x =- 9954 THEN
            sigmoid_f := 15;
        ELSIF x =- 9953 THEN
            sigmoid_f := 15;
        ELSIF x =- 9952 THEN
            sigmoid_f := 15;
        ELSIF x =- 9951 THEN
            sigmoid_f := 15;
        ELSIF x =- 9950 THEN
            sigmoid_f := 15;
        ELSIF x =- 9949 THEN
            sigmoid_f := 15;
        ELSIF x =- 9948 THEN
            sigmoid_f := 15;
        ELSIF x =- 9947 THEN
            sigmoid_f := 15;
        ELSIF x =- 9946 THEN
            sigmoid_f := 15;
        ELSIF x =- 9945 THEN
            sigmoid_f := 15;
        ELSIF x =- 9944 THEN
            sigmoid_f := 15;
        ELSIF x =- 9943 THEN
            sigmoid_f := 15;
        ELSIF x =- 9942 THEN
            sigmoid_f := 15;
        ELSIF x =- 9941 THEN
            sigmoid_f := 15;
        ELSIF x =- 9940 THEN
            sigmoid_f := 15;
        ELSIF x =- 9939 THEN
            sigmoid_f := 15;
        ELSIF x =- 9938 THEN
            sigmoid_f := 15;
        ELSIF x =- 9937 THEN
            sigmoid_f := 15;
        ELSIF x =- 9936 THEN
            sigmoid_f := 15;
        ELSIF x =- 9935 THEN
            sigmoid_f := 15;
        ELSIF x =- 9934 THEN
            sigmoid_f := 15;
        ELSIF x =- 9933 THEN
            sigmoid_f := 15;
        ELSIF x =- 9932 THEN
            sigmoid_f := 15;
        ELSIF x =- 9931 THEN
            sigmoid_f := 15;
        ELSIF x =- 9930 THEN
            sigmoid_f := 15;
        ELSIF x =- 9929 THEN
            sigmoid_f := 15;
        ELSIF x =- 9928 THEN
            sigmoid_f := 15;
        ELSIF x =- 9927 THEN
            sigmoid_f := 15;
        ELSIF x =- 9926 THEN
            sigmoid_f := 15;
        ELSIF x =- 9925 THEN
            sigmoid_f := 15;
        ELSIF x =- 9924 THEN
            sigmoid_f := 16;
        ELSIF x =- 9923 THEN
            sigmoid_f := 16;
        ELSIF x =- 9922 THEN
            sigmoid_f := 16;
        ELSIF x =- 9921 THEN
            sigmoid_f := 16;
        ELSIF x =- 9920 THEN
            sigmoid_f := 16;
        ELSIF x =- 9919 THEN
            sigmoid_f := 16;
        ELSIF x =- 9918 THEN
            sigmoid_f := 16;
        ELSIF x =- 9917 THEN
            sigmoid_f := 16;
        ELSIF x =- 9916 THEN
            sigmoid_f := 16;
        ELSIF x =- 9915 THEN
            sigmoid_f := 16;
        ELSIF x =- 9914 THEN
            sigmoid_f := 16;
        ELSIF x =- 9913 THEN
            sigmoid_f := 16;
        ELSIF x =- 9912 THEN
            sigmoid_f := 16;
        ELSIF x =- 9911 THEN
            sigmoid_f := 16;
        ELSIF x =- 9910 THEN
            sigmoid_f := 16;
        ELSIF x =- 9909 THEN
            sigmoid_f := 16;
        ELSIF x =- 9908 THEN
            sigmoid_f := 16;
        ELSIF x =- 9907 THEN
            sigmoid_f := 16;
        ELSIF x =- 9906 THEN
            sigmoid_f := 16;
        ELSIF x =- 9905 THEN
            sigmoid_f := 16;
        ELSIF x =- 9904 THEN
            sigmoid_f := 16;
        ELSIF x =- 9903 THEN
            sigmoid_f := 16;
        ELSIF x =- 9902 THEN
            sigmoid_f := 16;
        ELSIF x =- 9901 THEN
            sigmoid_f := 16;
        ELSIF x =- 9900 THEN
            sigmoid_f := 16;
        ELSIF x =- 9899 THEN
            sigmoid_f := 16;
        ELSIF x =- 9898 THEN
            sigmoid_f := 16;
        ELSIF x =- 9897 THEN
            sigmoid_f := 16;
        ELSIF x =- 9896 THEN
            sigmoid_f := 16;
        ELSIF x =- 9895 THEN
            sigmoid_f := 16;
        ELSIF x =- 9894 THEN
            sigmoid_f := 16;
        ELSIF x =- 9893 THEN
            sigmoid_f := 16;
        ELSIF x =- 9892 THEN
            sigmoid_f := 16;
        ELSIF x =- 9891 THEN
            sigmoid_f := 16;
        ELSIF x =- 9890 THEN
            sigmoid_f := 16;
        ELSIF x =- 9889 THEN
            sigmoid_f := 16;
        ELSIF x =- 9888 THEN
            sigmoid_f := 16;
        ELSIF x =- 9887 THEN
            sigmoid_f := 16;
        ELSIF x =- 9886 THEN
            sigmoid_f := 16;
        ELSIF x =- 9885 THEN
            sigmoid_f := 16;
        ELSIF x =- 9884 THEN
            sigmoid_f := 16;
        ELSIF x =- 9883 THEN
            sigmoid_f := 16;
        ELSIF x =- 9882 THEN
            sigmoid_f := 16;
        ELSIF x =- 9881 THEN
            sigmoid_f := 16;
        ELSIF x =- 9880 THEN
            sigmoid_f := 16;
        ELSIF x =- 9879 THEN
            sigmoid_f := 16;
        ELSIF x =- 9878 THEN
            sigmoid_f := 16;
        ELSIF x =- 9877 THEN
            sigmoid_f := 16;
        ELSIF x =- 9876 THEN
            sigmoid_f := 16;
        ELSIF x =- 9875 THEN
            sigmoid_f := 16;
        ELSIF x =- 9874 THEN
            sigmoid_f := 16;
        ELSIF x =- 9873 THEN
            sigmoid_f := 16;
        ELSIF x =- 9872 THEN
            sigmoid_f := 16;
        ELSIF x =- 9871 THEN
            sigmoid_f := 16;
        ELSIF x =- 9870 THEN
            sigmoid_f := 16;
        ELSIF x =- 9869 THEN
            sigmoid_f := 16;
        ELSIF x =- 9868 THEN
            sigmoid_f := 16;
        ELSIF x =- 9867 THEN
            sigmoid_f := 16;
        ELSIF x =- 9866 THEN
            sigmoid_f := 16;
        ELSIF x =- 9865 THEN
            sigmoid_f := 16;
        ELSIF x =- 9864 THEN
            sigmoid_f := 16;
        ELSIF x =- 9863 THEN
            sigmoid_f := 16;
        ELSIF x =- 9862 THEN
            sigmoid_f := 16;
        ELSIF x =- 9861 THEN
            sigmoid_f := 16;
        ELSIF x =- 9860 THEN
            sigmoid_f := 16;
        ELSIF x =- 9859 THEN
            sigmoid_f := 16;
        ELSIF x =- 9858 THEN
            sigmoid_f := 16;
        ELSIF x =- 9857 THEN
            sigmoid_f := 16;
        ELSIF x =- 9856 THEN
            sigmoid_f := 16;
        ELSIF x =- 9855 THEN
            sigmoid_f := 16;
        ELSIF x =- 9854 THEN
            sigmoid_f := 16;
        ELSIF x =- 9853 THEN
            sigmoid_f := 16;
        ELSIF x =- 9852 THEN
            sigmoid_f := 16;
        ELSIF x =- 9851 THEN
            sigmoid_f := 16;
        ELSIF x =- 9850 THEN
            sigmoid_f := 16;
        ELSIF x =- 9849 THEN
            sigmoid_f := 16;
        ELSIF x =- 9848 THEN
            sigmoid_f := 16;
        ELSIF x =- 9847 THEN
            sigmoid_f := 16;
        ELSIF x =- 9846 THEN
            sigmoid_f := 16;
        ELSIF x =- 9845 THEN
            sigmoid_f := 16;
        ELSIF x =- 9844 THEN
            sigmoid_f := 16;
        ELSIF x =- 9843 THEN
            sigmoid_f := 16;
        ELSIF x =- 9842 THEN
            sigmoid_f := 16;
        ELSIF x =- 9841 THEN
            sigmoid_f := 16;
        ELSIF x =- 9840 THEN
            sigmoid_f := 16;
        ELSIF x =- 9839 THEN
            sigmoid_f := 16;
        ELSIF x =- 9838 THEN
            sigmoid_f := 16;
        ELSIF x =- 9837 THEN
            sigmoid_f := 16;
        ELSIF x =- 9836 THEN
            sigmoid_f := 16;
        ELSIF x =- 9835 THEN
            sigmoid_f := 16;
        ELSIF x =- 9834 THEN
            sigmoid_f := 16;
        ELSIF x =- 9833 THEN
            sigmoid_f := 16;
        ELSIF x =- 9832 THEN
            sigmoid_f := 16;
        ELSIF x =- 9831 THEN
            sigmoid_f := 16;
        ELSIF x =- 9830 THEN
            sigmoid_f := 16;
        ELSIF x =- 9829 THEN
            sigmoid_f := 16;
        ELSIF x =- 9828 THEN
            sigmoid_f := 16;
        ELSIF x =- 9827 THEN
            sigmoid_f := 16;
        ELSIF x =- 9826 THEN
            sigmoid_f := 16;
        ELSIF x =- 9825 THEN
            sigmoid_f := 16;
        ELSIF x =- 9824 THEN
            sigmoid_f := 16;
        ELSIF x =- 9823 THEN
            sigmoid_f := 16;
        ELSIF x =- 9822 THEN
            sigmoid_f := 16;
        ELSIF x =- 9821 THEN
            sigmoid_f := 16;
        ELSIF x =- 9820 THEN
            sigmoid_f := 16;
        ELSIF x =- 9819 THEN
            sigmoid_f := 16;
        ELSIF x =- 9818 THEN
            sigmoid_f := 16;
        ELSIF x =- 9817 THEN
            sigmoid_f := 16;
        ELSIF x =- 9816 THEN
            sigmoid_f := 16;
        ELSIF x =- 9815 THEN
            sigmoid_f := 16;
        ELSIF x =- 9814 THEN
            sigmoid_f := 16;
        ELSIF x =- 9813 THEN
            sigmoid_f := 16;
        ELSIF x =- 9812 THEN
            sigmoid_f := 16;
        ELSIF x =- 9811 THEN
            sigmoid_f := 16;
        ELSIF x =- 9810 THEN
            sigmoid_f := 16;
        ELSIF x =- 9809 THEN
            sigmoid_f := 16;
        ELSIF x =- 9808 THEN
            sigmoid_f := 16;
        ELSIF x =- 9807 THEN
            sigmoid_f := 16;
        ELSIF x =- 9806 THEN
            sigmoid_f := 16;
        ELSIF x =- 9805 THEN
            sigmoid_f := 16;
        ELSIF x =- 9804 THEN
            sigmoid_f := 16;
        ELSIF x =- 9803 THEN
            sigmoid_f := 16;
        ELSIF x =- 9802 THEN
            sigmoid_f := 16;
        ELSIF x =- 9801 THEN
            sigmoid_f := 16;
        ELSIF x =- 9800 THEN
            sigmoid_f := 16;
        ELSIF x =- 9799 THEN
            sigmoid_f := 16;
        ELSIF x =- 9798 THEN
            sigmoid_f := 16;
        ELSIF x =- 9797 THEN
            sigmoid_f := 16;
        ELSIF x =- 9796 THEN
            sigmoid_f := 16;
        ELSIF x =- 9795 THEN
            sigmoid_f := 16;
        ELSIF x =- 9794 THEN
            sigmoid_f := 16;
        ELSIF x =- 9793 THEN
            sigmoid_f := 16;
        ELSIF x =- 9792 THEN
            sigmoid_f := 16;
        ELSIF x =- 9791 THEN
            sigmoid_f := 16;
        ELSIF x =- 9790 THEN
            sigmoid_f := 16;
        ELSIF x =- 9789 THEN
            sigmoid_f := 16;
        ELSIF x =- 9788 THEN
            sigmoid_f := 16;
        ELSIF x =- 9787 THEN
            sigmoid_f := 16;
        ELSIF x =- 9786 THEN
            sigmoid_f := 16;
        ELSIF x =- 9785 THEN
            sigmoid_f := 16;
        ELSIF x =- 9784 THEN
            sigmoid_f := 16;
        ELSIF x =- 9783 THEN
            sigmoid_f := 16;
        ELSIF x =- 9782 THEN
            sigmoid_f := 16;
        ELSIF x =- 9781 THEN
            sigmoid_f := 16;
        ELSIF x =- 9780 THEN
            sigmoid_f := 16;
        ELSIF x =- 9779 THEN
            sigmoid_f := 16;
        ELSIF x =- 9778 THEN
            sigmoid_f := 16;
        ELSIF x =- 9777 THEN
            sigmoid_f := 16;
        ELSIF x =- 9776 THEN
            sigmoid_f := 16;
        ELSIF x =- 9775 THEN
            sigmoid_f := 16;
        ELSIF x =- 9774 THEN
            sigmoid_f := 16;
        ELSIF x =- 9773 THEN
            sigmoid_f := 16;
        ELSIF x =- 9772 THEN
            sigmoid_f := 16;
        ELSIF x =- 9771 THEN
            sigmoid_f := 16;
        ELSIF x =- 9770 THEN
            sigmoid_f := 16;
        ELSIF x =- 9769 THEN
            sigmoid_f := 16;
        ELSIF x =- 9768 THEN
            sigmoid_f := 16;
        ELSIF x =- 9767 THEN
            sigmoid_f := 17;
        ELSIF x =- 9766 THEN
            sigmoid_f := 17;
        ELSIF x =- 9765 THEN
            sigmoid_f := 17;
        ELSIF x =- 9764 THEN
            sigmoid_f := 17;
        ELSIF x =- 9763 THEN
            sigmoid_f := 17;
        ELSIF x =- 9762 THEN
            sigmoid_f := 17;
        ELSIF x =- 9761 THEN
            sigmoid_f := 17;
        ELSIF x =- 9760 THEN
            sigmoid_f := 17;
        ELSIF x =- 9759 THEN
            sigmoid_f := 17;
        ELSIF x =- 9758 THEN
            sigmoid_f := 17;
        ELSIF x =- 9757 THEN
            sigmoid_f := 17;
        ELSIF x =- 9756 THEN
            sigmoid_f := 17;
        ELSIF x =- 9755 THEN
            sigmoid_f := 17;
        ELSIF x =- 9754 THEN
            sigmoid_f := 17;
        ELSIF x =- 9753 THEN
            sigmoid_f := 17;
        ELSIF x =- 9752 THEN
            sigmoid_f := 17;
        ELSIF x =- 9751 THEN
            sigmoid_f := 17;
        ELSIF x =- 9750 THEN
            sigmoid_f := 17;
        ELSIF x =- 9749 THEN
            sigmoid_f := 17;
        ELSIF x =- 9748 THEN
            sigmoid_f := 17;
        ELSIF x =- 9747 THEN
            sigmoid_f := 17;
        ELSIF x =- 9746 THEN
            sigmoid_f := 17;
        ELSIF x =- 9745 THEN
            sigmoid_f := 17;
        ELSIF x =- 9744 THEN
            sigmoid_f := 17;
        ELSIF x =- 9743 THEN
            sigmoid_f := 17;
        ELSIF x =- 9742 THEN
            sigmoid_f := 17;
        ELSIF x =- 9741 THEN
            sigmoid_f := 17;
        ELSIF x =- 9740 THEN
            sigmoid_f := 17;
        ELSIF x =- 9739 THEN
            sigmoid_f := 17;
        ELSIF x =- 9738 THEN
            sigmoid_f := 17;
        ELSIF x =- 9737 THEN
            sigmoid_f := 17;
        ELSIF x =- 9736 THEN
            sigmoid_f := 17;
        ELSIF x =- 9735 THEN
            sigmoid_f := 17;
        ELSIF x =- 9734 THEN
            sigmoid_f := 17;
        ELSIF x =- 9733 THEN
            sigmoid_f := 17;
        ELSIF x =- 9732 THEN
            sigmoid_f := 17;
        ELSIF x =- 9731 THEN
            sigmoid_f := 17;
        ELSIF x =- 9730 THEN
            sigmoid_f := 17;
        ELSIF x =- 9729 THEN
            sigmoid_f := 17;
        ELSIF x =- 9728 THEN
            sigmoid_f := 17;
        ELSIF x =- 9727 THEN
            sigmoid_f := 17;
        ELSIF x =- 9726 THEN
            sigmoid_f := 17;
        ELSIF x =- 9725 THEN
            sigmoid_f := 17;
        ELSIF x =- 9724 THEN
            sigmoid_f := 17;
        ELSIF x =- 9723 THEN
            sigmoid_f := 17;
        ELSIF x =- 9722 THEN
            sigmoid_f := 17;
        ELSIF x =- 9721 THEN
            sigmoid_f := 17;
        ELSIF x =- 9720 THEN
            sigmoid_f := 17;
        ELSIF x =- 9719 THEN
            sigmoid_f := 17;
        ELSIF x =- 9718 THEN
            sigmoid_f := 17;
        ELSIF x =- 9717 THEN
            sigmoid_f := 17;
        ELSIF x =- 9716 THEN
            sigmoid_f := 17;
        ELSIF x =- 9715 THEN
            sigmoid_f := 17;
        ELSIF x =- 9714 THEN
            sigmoid_f := 17;
        ELSIF x =- 9713 THEN
            sigmoid_f := 17;
        ELSIF x =- 9712 THEN
            sigmoid_f := 17;
        ELSIF x =- 9711 THEN
            sigmoid_f := 17;
        ELSIF x =- 9710 THEN
            sigmoid_f := 17;
        ELSIF x =- 9709 THEN
            sigmoid_f := 17;
        ELSIF x =- 9708 THEN
            sigmoid_f := 17;
        ELSIF x =- 9707 THEN
            sigmoid_f := 17;
        ELSIF x =- 9706 THEN
            sigmoid_f := 17;
        ELSIF x =- 9705 THEN
            sigmoid_f := 17;
        ELSIF x =- 9704 THEN
            sigmoid_f := 17;
        ELSIF x =- 9703 THEN
            sigmoid_f := 17;
        ELSIF x =- 9702 THEN
            sigmoid_f := 17;
        ELSIF x =- 9701 THEN
            sigmoid_f := 17;
        ELSIF x =- 9700 THEN
            sigmoid_f := 17;
        ELSIF x =- 9699 THEN
            sigmoid_f := 17;
        ELSIF x =- 9698 THEN
            sigmoid_f := 17;
        ELSIF x =- 9697 THEN
            sigmoid_f := 17;
        ELSIF x =- 9696 THEN
            sigmoid_f := 17;
        ELSIF x =- 9695 THEN
            sigmoid_f := 17;
        ELSIF x =- 9694 THEN
            sigmoid_f := 17;
        ELSIF x =- 9693 THEN
            sigmoid_f := 17;
        ELSIF x =- 9692 THEN
            sigmoid_f := 17;
        ELSIF x =- 9691 THEN
            sigmoid_f := 17;
        ELSIF x =- 9690 THEN
            sigmoid_f := 17;
        ELSIF x =- 9689 THEN
            sigmoid_f := 17;
        ELSIF x =- 9688 THEN
            sigmoid_f := 17;
        ELSIF x =- 9687 THEN
            sigmoid_f := 17;
        ELSIF x =- 9686 THEN
            sigmoid_f := 17;
        ELSIF x =- 9685 THEN
            sigmoid_f := 17;
        ELSIF x =- 9684 THEN
            sigmoid_f := 17;
        ELSIF x =- 9683 THEN
            sigmoid_f := 17;
        ELSIF x =- 9682 THEN
            sigmoid_f := 17;
        ELSIF x =- 9681 THEN
            sigmoid_f := 17;
        ELSIF x =- 9680 THEN
            sigmoid_f := 17;
        ELSIF x =- 9679 THEN
            sigmoid_f := 17;
        ELSIF x =- 9678 THEN
            sigmoid_f := 17;
        ELSIF x =- 9677 THEN
            sigmoid_f := 17;
        ELSIF x =- 9676 THEN
            sigmoid_f := 17;
        ELSIF x =- 9675 THEN
            sigmoid_f := 17;
        ELSIF x =- 9674 THEN
            sigmoid_f := 17;
        ELSIF x =- 9673 THEN
            sigmoid_f := 17;
        ELSIF x =- 9672 THEN
            sigmoid_f := 17;
        ELSIF x =- 9671 THEN
            sigmoid_f := 17;
        ELSIF x =- 9670 THEN
            sigmoid_f := 17;
        ELSIF x =- 9669 THEN
            sigmoid_f := 17;
        ELSIF x =- 9668 THEN
            sigmoid_f := 17;
        ELSIF x =- 9667 THEN
            sigmoid_f := 17;
        ELSIF x =- 9666 THEN
            sigmoid_f := 17;
        ELSIF x =- 9665 THEN
            sigmoid_f := 17;
        ELSIF x =- 9664 THEN
            sigmoid_f := 17;
        ELSIF x =- 9663 THEN
            sigmoid_f := 17;
        ELSIF x =- 9662 THEN
            sigmoid_f := 17;
        ELSIF x =- 9661 THEN
            sigmoid_f := 17;
        ELSIF x =- 9660 THEN
            sigmoid_f := 17;
        ELSIF x =- 9659 THEN
            sigmoid_f := 17;
        ELSIF x =- 9658 THEN
            sigmoid_f := 17;
        ELSIF x =- 9657 THEN
            sigmoid_f := 17;
        ELSIF x =- 9656 THEN
            sigmoid_f := 17;
        ELSIF x =- 9655 THEN
            sigmoid_f := 17;
        ELSIF x =- 9654 THEN
            sigmoid_f := 18;
        ELSIF x =- 9653 THEN
            sigmoid_f := 18;
        ELSIF x =- 9652 THEN
            sigmoid_f := 18;
        ELSIF x =- 9651 THEN
            sigmoid_f := 18;
        ELSIF x =- 9650 THEN
            sigmoid_f := 18;
        ELSIF x =- 9649 THEN
            sigmoid_f := 18;
        ELSIF x =- 9648 THEN
            sigmoid_f := 18;
        ELSIF x =- 9647 THEN
            sigmoid_f := 18;
        ELSIF x =- 9646 THEN
            sigmoid_f := 18;
        ELSIF x =- 9645 THEN
            sigmoid_f := 18;
        ELSIF x =- 9644 THEN
            sigmoid_f := 18;
        ELSIF x =- 9643 THEN
            sigmoid_f := 18;
        ELSIF x =- 9642 THEN
            sigmoid_f := 18;
        ELSIF x =- 9641 THEN
            sigmoid_f := 18;
        ELSIF x =- 9640 THEN
            sigmoid_f := 18;
        ELSIF x =- 9639 THEN
            sigmoid_f := 18;
        ELSIF x =- 9638 THEN
            sigmoid_f := 18;
        ELSIF x =- 9637 THEN
            sigmoid_f := 18;
        ELSIF x =- 9636 THEN
            sigmoid_f := 18;
        ELSIF x =- 9635 THEN
            sigmoid_f := 18;
        ELSIF x =- 9634 THEN
            sigmoid_f := 18;
        ELSIF x =- 9633 THEN
            sigmoid_f := 18;
        ELSIF x =- 9632 THEN
            sigmoid_f := 18;
        ELSIF x =- 9631 THEN
            sigmoid_f := 18;
        ELSIF x =- 9630 THEN
            sigmoid_f := 18;
        ELSIF x =- 9629 THEN
            sigmoid_f := 18;
        ELSIF x =- 9628 THEN
            sigmoid_f := 18;
        ELSIF x =- 9627 THEN
            sigmoid_f := 18;
        ELSIF x =- 9626 THEN
            sigmoid_f := 18;
        ELSIF x =- 9625 THEN
            sigmoid_f := 18;
        ELSIF x =- 9624 THEN
            sigmoid_f := 18;
        ELSIF x =- 9623 THEN
            sigmoid_f := 18;
        ELSIF x =- 9622 THEN
            sigmoid_f := 18;
        ELSIF x =- 9621 THEN
            sigmoid_f := 18;
        ELSIF x =- 9620 THEN
            sigmoid_f := 18;
        ELSIF x =- 9619 THEN
            sigmoid_f := 18;
        ELSIF x =- 9618 THEN
            sigmoid_f := 18;
        ELSIF x =- 9617 THEN
            sigmoid_f := 18;
        ELSIF x =- 9616 THEN
            sigmoid_f := 18;
        ELSIF x =- 9615 THEN
            sigmoid_f := 18;
        ELSIF x =- 9614 THEN
            sigmoid_f := 18;
        ELSIF x =- 9613 THEN
            sigmoid_f := 18;
        ELSIF x =- 9612 THEN
            sigmoid_f := 18;
        ELSIF x =- 9611 THEN
            sigmoid_f := 18;
        ELSIF x =- 9610 THEN
            sigmoid_f := 18;
        ELSIF x =- 9609 THEN
            sigmoid_f := 18;
        ELSIF x =- 9608 THEN
            sigmoid_f := 18;
        ELSIF x =- 9607 THEN
            sigmoid_f := 18;
        ELSIF x =- 9606 THEN
            sigmoid_f := 18;
        ELSIF x =- 9605 THEN
            sigmoid_f := 18;
        ELSIF x =- 9604 THEN
            sigmoid_f := 18;
        ELSIF x =- 9603 THEN
            sigmoid_f := 18;
        ELSIF x =- 9602 THEN
            sigmoid_f := 18;
        ELSIF x =- 9601 THEN
            sigmoid_f := 18;
        ELSIF x =- 9600 THEN
            sigmoid_f := 18;
        ELSIF x =- 9599 THEN
            sigmoid_f := 18;
        ELSIF x =- 9598 THEN
            sigmoid_f := 18;
        ELSIF x =- 9597 THEN
            sigmoid_f := 18;
        ELSIF x =- 9596 THEN
            sigmoid_f := 18;
        ELSIF x =- 9595 THEN
            sigmoid_f := 18;
        ELSIF x =- 9594 THEN
            sigmoid_f := 18;
        ELSIF x =- 9593 THEN
            sigmoid_f := 18;
        ELSIF x =- 9592 THEN
            sigmoid_f := 18;
        ELSIF x =- 9591 THEN
            sigmoid_f := 18;
        ELSIF x =- 9590 THEN
            sigmoid_f := 18;
        ELSIF x =- 9589 THEN
            sigmoid_f := 18;
        ELSIF x =- 9588 THEN
            sigmoid_f := 18;
        ELSIF x =- 9587 THEN
            sigmoid_f := 18;
        ELSIF x =- 9586 THEN
            sigmoid_f := 18;
        ELSIF x =- 9585 THEN
            sigmoid_f := 18;
        ELSIF x =- 9584 THEN
            sigmoid_f := 18;
        ELSIF x =- 9583 THEN
            sigmoid_f := 18;
        ELSIF x =- 9582 THEN
            sigmoid_f := 18;
        ELSIF x =- 9581 THEN
            sigmoid_f := 18;
        ELSIF x =- 9580 THEN
            sigmoid_f := 18;
        ELSIF x =- 9579 THEN
            sigmoid_f := 18;
        ELSIF x =- 9578 THEN
            sigmoid_f := 18;
        ELSIF x =- 9577 THEN
            sigmoid_f := 18;
        ELSIF x =- 9576 THEN
            sigmoid_f := 18;
        ELSIF x =- 9575 THEN
            sigmoid_f := 18;
        ELSIF x =- 9574 THEN
            sigmoid_f := 18;
        ELSIF x =- 9573 THEN
            sigmoid_f := 18;
        ELSIF x =- 9572 THEN
            sigmoid_f := 18;
        ELSIF x =- 9571 THEN
            sigmoid_f := 18;
        ELSIF x =- 9570 THEN
            sigmoid_f := 18;
        ELSIF x =- 9569 THEN
            sigmoid_f := 18;
        ELSIF x =- 9568 THEN
            sigmoid_f := 18;
        ELSIF x =- 9567 THEN
            sigmoid_f := 18;
        ELSIF x =- 9566 THEN
            sigmoid_f := 18;
        ELSIF x =- 9565 THEN
            sigmoid_f := 18;
        ELSIF x =- 9564 THEN
            sigmoid_f := 18;
        ELSIF x =- 9563 THEN
            sigmoid_f := 18;
        ELSIF x =- 9562 THEN
            sigmoid_f := 18;
        ELSIF x =- 9561 THEN
            sigmoid_f := 18;
        ELSIF x =- 9560 THEN
            sigmoid_f := 18;
        ELSIF x =- 9559 THEN
            sigmoid_f := 18;
        ELSIF x =- 9558 THEN
            sigmoid_f := 18;
        ELSIF x =- 9557 THEN
            sigmoid_f := 19;
        ELSIF x =- 9556 THEN
            sigmoid_f := 19;
        ELSIF x =- 9555 THEN
            sigmoid_f := 19;
        ELSIF x =- 9554 THEN
            sigmoid_f := 19;
        ELSIF x =- 9553 THEN
            sigmoid_f := 19;
        ELSIF x =- 9552 THEN
            sigmoid_f := 19;
        ELSIF x =- 9551 THEN
            sigmoid_f := 19;
        ELSIF x =- 9550 THEN
            sigmoid_f := 19;
        ELSIF x =- 9549 THEN
            sigmoid_f := 19;
        ELSIF x =- 9548 THEN
            sigmoid_f := 19;
        ELSIF x =- 9547 THEN
            sigmoid_f := 19;
        ELSIF x =- 9546 THEN
            sigmoid_f := 19;
        ELSIF x =- 9545 THEN
            sigmoid_f := 19;
        ELSIF x =- 9544 THEN
            sigmoid_f := 19;
        ELSIF x =- 9543 THEN
            sigmoid_f := 19;
        ELSIF x =- 9542 THEN
            sigmoid_f := 19;
        ELSIF x =- 9541 THEN
            sigmoid_f := 19;
        ELSIF x =- 9540 THEN
            sigmoid_f := 19;
        ELSIF x =- 9539 THEN
            sigmoid_f := 19;
        ELSIF x =- 9538 THEN
            sigmoid_f := 19;
        ELSIF x =- 9537 THEN
            sigmoid_f := 19;
        ELSIF x =- 9536 THEN
            sigmoid_f := 19;
        ELSIF x =- 9535 THEN
            sigmoid_f := 19;
        ELSIF x =- 9534 THEN
            sigmoid_f := 19;
        ELSIF x =- 9533 THEN
            sigmoid_f := 19;
        ELSIF x =- 9532 THEN
            sigmoid_f := 19;
        ELSIF x =- 9531 THEN
            sigmoid_f := 19;
        ELSIF x =- 9530 THEN
            sigmoid_f := 19;
        ELSIF x =- 9529 THEN
            sigmoid_f := 19;
        ELSIF x =- 9528 THEN
            sigmoid_f := 19;
        ELSIF x =- 9527 THEN
            sigmoid_f := 19;
        ELSIF x =- 9526 THEN
            sigmoid_f := 19;
        ELSIF x =- 9525 THEN
            sigmoid_f := 19;
        ELSIF x =- 9524 THEN
            sigmoid_f := 19;
        ELSIF x =- 9523 THEN
            sigmoid_f := 19;
        ELSIF x =- 9522 THEN
            sigmoid_f := 19;
        ELSIF x =- 9521 THEN
            sigmoid_f := 19;
        ELSIF x =- 9520 THEN
            sigmoid_f := 19;
        ELSIF x =- 9519 THEN
            sigmoid_f := 19;
        ELSIF x =- 9518 THEN
            sigmoid_f := 19;
        ELSIF x =- 9517 THEN
            sigmoid_f := 19;
        ELSIF x =- 9516 THEN
            sigmoid_f := 19;
        ELSIF x =- 9515 THEN
            sigmoid_f := 19;
        ELSIF x =- 9514 THEN
            sigmoid_f := 19;
        ELSIF x =- 9513 THEN
            sigmoid_f := 19;
        ELSIF x =- 9512 THEN
            sigmoid_f := 19;
        ELSIF x =- 9511 THEN
            sigmoid_f := 19;
        ELSIF x =- 9510 THEN
            sigmoid_f := 19;
        ELSIF x =- 9509 THEN
            sigmoid_f := 19;
        ELSIF x =- 9508 THEN
            sigmoid_f := 19;
        ELSIF x =- 9507 THEN
            sigmoid_f := 19;
        ELSIF x =- 9506 THEN
            sigmoid_f := 19;
        ELSIF x =- 9505 THEN
            sigmoid_f := 19;
        ELSIF x =- 9504 THEN
            sigmoid_f := 19;
        ELSIF x =- 9503 THEN
            sigmoid_f := 19;
        ELSIF x =- 9502 THEN
            sigmoid_f := 19;
        ELSIF x =- 9501 THEN
            sigmoid_f := 19;
        ELSIF x =- 9500 THEN
            sigmoid_f := 19;
        ELSIF x =- 9499 THEN
            sigmoid_f := 19;
        ELSIF x =- 9498 THEN
            sigmoid_f := 19;
        ELSIF x =- 9497 THEN
            sigmoid_f := 19;
        ELSIF x =- 9496 THEN
            sigmoid_f := 19;
        ELSIF x =- 9495 THEN
            sigmoid_f := 19;
        ELSIF x =- 9494 THEN
            sigmoid_f := 19;
        ELSIF x =- 9493 THEN
            sigmoid_f := 19;
        ELSIF x =- 9492 THEN
            sigmoid_f := 19;
        ELSIF x =- 9491 THEN
            sigmoid_f := 19;
        ELSIF x =- 9490 THEN
            sigmoid_f := 19;
        ELSIF x =- 9489 THEN
            sigmoid_f := 19;
        ELSIF x =- 9488 THEN
            sigmoid_f := 19;
        ELSIF x =- 9487 THEN
            sigmoid_f := 19;
        ELSIF x =- 9486 THEN
            sigmoid_f := 19;
        ELSIF x =- 9485 THEN
            sigmoid_f := 19;
        ELSIF x =- 9484 THEN
            sigmoid_f := 19;
        ELSIF x =- 9483 THEN
            sigmoid_f := 19;
        ELSIF x =- 9482 THEN
            sigmoid_f := 19;
        ELSIF x =- 9481 THEN
            sigmoid_f := 19;
        ELSIF x =- 9480 THEN
            sigmoid_f := 19;
        ELSIF x =- 9479 THEN
            sigmoid_f := 19;
        ELSIF x =- 9478 THEN
            sigmoid_f := 19;
        ELSIF x =- 9477 THEN
            sigmoid_f := 19;
        ELSIF x =- 9476 THEN
            sigmoid_f := 19;
        ELSIF x =- 9475 THEN
            sigmoid_f := 19;
        ELSIF x =- 9474 THEN
            sigmoid_f := 19;
        ELSIF x =- 9473 THEN
            sigmoid_f := 19;
        ELSIF x =- 9472 THEN
            sigmoid_f := 19;
        ELSIF x =- 9471 THEN
            sigmoid_f := 19;
        ELSIF x =- 9470 THEN
            sigmoid_f := 19;
        ELSIF x =- 9469 THEN
            sigmoid_f := 19;
        ELSIF x =- 9468 THEN
            sigmoid_f := 19;
        ELSIF x =- 9467 THEN
            sigmoid_f := 19;
        ELSIF x =- 9466 THEN
            sigmoid_f := 19;
        ELSIF x =- 9465 THEN
            sigmoid_f := 19;
        ELSIF x =- 9464 THEN
            sigmoid_f := 19;
        ELSIF x =- 9463 THEN
            sigmoid_f := 19;
        ELSIF x =- 9462 THEN
            sigmoid_f := 19;
        ELSIF x =- 9461 THEN
            sigmoid_f := 19;
        ELSIF x =- 9460 THEN
            sigmoid_f := 19;
        ELSIF x =- 9459 THEN
            sigmoid_f := 20;
        ELSIF x =- 9458 THEN
            sigmoid_f := 20;
        ELSIF x =- 9457 THEN
            sigmoid_f := 20;
        ELSIF x =- 9456 THEN
            sigmoid_f := 20;
        ELSIF x =- 9455 THEN
            sigmoid_f := 20;
        ELSIF x =- 9454 THEN
            sigmoid_f := 20;
        ELSIF x =- 9453 THEN
            sigmoid_f := 20;
        ELSIF x =- 9452 THEN
            sigmoid_f := 20;
        ELSIF x =- 9451 THEN
            sigmoid_f := 20;
        ELSIF x =- 9450 THEN
            sigmoid_f := 20;
        ELSIF x =- 9449 THEN
            sigmoid_f := 20;
        ELSIF x =- 9448 THEN
            sigmoid_f := 20;
        ELSIF x =- 9447 THEN
            sigmoid_f := 20;
        ELSIF x =- 9446 THEN
            sigmoid_f := 20;
        ELSIF x =- 9445 THEN
            sigmoid_f := 20;
        ELSIF x =- 9444 THEN
            sigmoid_f := 20;
        ELSIF x =- 9443 THEN
            sigmoid_f := 20;
        ELSIF x =- 9442 THEN
            sigmoid_f := 20;
        ELSIF x =- 9441 THEN
            sigmoid_f := 20;
        ELSIF x =- 9440 THEN
            sigmoid_f := 20;
        ELSIF x =- 9439 THEN
            sigmoid_f := 20;
        ELSIF x =- 9438 THEN
            sigmoid_f := 20;
        ELSIF x =- 9437 THEN
            sigmoid_f := 20;
        ELSIF x =- 9436 THEN
            sigmoid_f := 20;
        ELSIF x =- 9435 THEN
            sigmoid_f := 20;
        ELSIF x =- 9434 THEN
            sigmoid_f := 20;
        ELSIF x =- 9433 THEN
            sigmoid_f := 20;
        ELSIF x =- 9432 THEN
            sigmoid_f := 20;
        ELSIF x =- 9431 THEN
            sigmoid_f := 20;
        ELSIF x =- 9430 THEN
            sigmoid_f := 20;
        ELSIF x =- 9429 THEN
            sigmoid_f := 20;
        ELSIF x =- 9428 THEN
            sigmoid_f := 20;
        ELSIF x =- 9427 THEN
            sigmoid_f := 20;
        ELSIF x =- 9426 THEN
            sigmoid_f := 20;
        ELSIF x =- 9425 THEN
            sigmoid_f := 20;
        ELSIF x =- 9424 THEN
            sigmoid_f := 20;
        ELSIF x =- 9423 THEN
            sigmoid_f := 20;
        ELSIF x =- 9422 THEN
            sigmoid_f := 20;
        ELSIF x =- 9421 THEN
            sigmoid_f := 20;
        ELSIF x =- 9420 THEN
            sigmoid_f := 20;
        ELSIF x =- 9419 THEN
            sigmoid_f := 20;
        ELSIF x =- 9418 THEN
            sigmoid_f := 20;
        ELSIF x =- 9417 THEN
            sigmoid_f := 20;
        ELSIF x =- 9416 THEN
            sigmoid_f := 20;
        ELSIF x =- 9415 THEN
            sigmoid_f := 20;
        ELSIF x =- 9414 THEN
            sigmoid_f := 20;
        ELSIF x =- 9413 THEN
            sigmoid_f := 20;
        ELSIF x =- 9412 THEN
            sigmoid_f := 20;
        ELSIF x =- 9411 THEN
            sigmoid_f := 20;
        ELSIF x =- 9410 THEN
            sigmoid_f := 20;
        ELSIF x =- 9409 THEN
            sigmoid_f := 20;
        ELSIF x =- 9408 THEN
            sigmoid_f := 20;
        ELSIF x =- 9407 THEN
            sigmoid_f := 20;
        ELSIF x =- 9406 THEN
            sigmoid_f := 20;
        ELSIF x =- 9405 THEN
            sigmoid_f := 20;
        ELSIF x =- 9404 THEN
            sigmoid_f := 20;
        ELSIF x =- 9403 THEN
            sigmoid_f := 20;
        ELSIF x =- 9402 THEN
            sigmoid_f := 20;
        ELSIF x =- 9401 THEN
            sigmoid_f := 20;
        ELSIF x =- 9400 THEN
            sigmoid_f := 20;
        ELSIF x =- 9399 THEN
            sigmoid_f := 20;
        ELSIF x =- 9398 THEN
            sigmoid_f := 20;
        ELSIF x =- 9397 THEN
            sigmoid_f := 20;
        ELSIF x =- 9396 THEN
            sigmoid_f := 20;
        ELSIF x =- 9395 THEN
            sigmoid_f := 20;
        ELSIF x =- 9394 THEN
            sigmoid_f := 20;
        ELSIF x =- 9393 THEN
            sigmoid_f := 20;
        ELSIF x =- 9392 THEN
            sigmoid_f := 20;
        ELSIF x =- 9391 THEN
            sigmoid_f := 20;
        ELSIF x =- 9390 THEN
            sigmoid_f := 20;
        ELSIF x =- 9389 THEN
            sigmoid_f := 20;
        ELSIF x =- 9388 THEN
            sigmoid_f := 20;
        ELSIF x =- 9387 THEN
            sigmoid_f := 20;
        ELSIF x =- 9386 THEN
            sigmoid_f := 20;
        ELSIF x =- 9385 THEN
            sigmoid_f := 20;
        ELSIF x =- 9384 THEN
            sigmoid_f := 20;
        ELSIF x =- 9383 THEN
            sigmoid_f := 20;
        ELSIF x =- 9382 THEN
            sigmoid_f := 20;
        ELSIF x =- 9381 THEN
            sigmoid_f := 20;
        ELSIF x =- 9380 THEN
            sigmoid_f := 20;
        ELSIF x =- 9379 THEN
            sigmoid_f := 20;
        ELSIF x =- 9378 THEN
            sigmoid_f := 20;
        ELSIF x =- 9377 THEN
            sigmoid_f := 20;
        ELSIF x =- 9376 THEN
            sigmoid_f := 20;
        ELSIF x =- 9375 THEN
            sigmoid_f := 20;
        ELSIF x =- 9374 THEN
            sigmoid_f := 20;
        ELSIF x =- 9373 THEN
            sigmoid_f := 20;
        ELSIF x =- 9372 THEN
            sigmoid_f := 20;
        ELSIF x =- 9371 THEN
            sigmoid_f := 20;
        ELSIF x =- 9370 THEN
            sigmoid_f := 20;
        ELSIF x =- 9369 THEN
            sigmoid_f := 20;
        ELSIF x =- 9368 THEN
            sigmoid_f := 20;
        ELSIF x =- 9367 THEN
            sigmoid_f := 20;
        ELSIF x =- 9366 THEN
            sigmoid_f := 20;
        ELSIF x =- 9365 THEN
            sigmoid_f := 20;
        ELSIF x =- 9364 THEN
            sigmoid_f := 20;
        ELSIF x =- 9363 THEN
            sigmoid_f := 20;
        ELSIF x =- 9362 THEN
            sigmoid_f := 21;
        ELSIF x =- 9361 THEN
            sigmoid_f := 21;
        ELSIF x =- 9360 THEN
            sigmoid_f := 21;
        ELSIF x =- 9359 THEN
            sigmoid_f := 21;
        ELSIF x =- 9358 THEN
            sigmoid_f := 21;
        ELSIF x =- 9357 THEN
            sigmoid_f := 21;
        ELSIF x =- 9356 THEN
            sigmoid_f := 21;
        ELSIF x =- 9355 THEN
            sigmoid_f := 21;
        ELSIF x =- 9354 THEN
            sigmoid_f := 21;
        ELSIF x =- 9353 THEN
            sigmoid_f := 21;
        ELSIF x =- 9352 THEN
            sigmoid_f := 21;
        ELSIF x =- 9351 THEN
            sigmoid_f := 21;
        ELSIF x =- 9350 THEN
            sigmoid_f := 21;
        ELSIF x =- 9349 THEN
            sigmoid_f := 21;
        ELSIF x =- 9348 THEN
            sigmoid_f := 21;
        ELSIF x =- 9347 THEN
            sigmoid_f := 21;
        ELSIF x =- 9346 THEN
            sigmoid_f := 21;
        ELSIF x =- 9345 THEN
            sigmoid_f := 21;
        ELSIF x =- 9344 THEN
            sigmoid_f := 21;
        ELSIF x =- 9343 THEN
            sigmoid_f := 21;
        ELSIF x =- 9342 THEN
            sigmoid_f := 21;
        ELSIF x =- 9341 THEN
            sigmoid_f := 21;
        ELSIF x =- 9340 THEN
            sigmoid_f := 21;
        ELSIF x =- 9339 THEN
            sigmoid_f := 21;
        ELSIF x =- 9338 THEN
            sigmoid_f := 21;
        ELSIF x =- 9337 THEN
            sigmoid_f := 21;
        ELSIF x =- 9336 THEN
            sigmoid_f := 21;
        ELSIF x =- 9335 THEN
            sigmoid_f := 21;
        ELSIF x =- 9334 THEN
            sigmoid_f := 21;
        ELSIF x =- 9333 THEN
            sigmoid_f := 21;
        ELSIF x =- 9332 THEN
            sigmoid_f := 21;
        ELSIF x =- 9331 THEN
            sigmoid_f := 21;
        ELSIF x =- 9330 THEN
            sigmoid_f := 21;
        ELSIF x =- 9329 THEN
            sigmoid_f := 21;
        ELSIF x =- 9328 THEN
            sigmoid_f := 21;
        ELSIF x =- 9327 THEN
            sigmoid_f := 21;
        ELSIF x =- 9326 THEN
            sigmoid_f := 21;
        ELSIF x =- 9325 THEN
            sigmoid_f := 21;
        ELSIF x =- 9324 THEN
            sigmoid_f := 21;
        ELSIF x =- 9323 THEN
            sigmoid_f := 21;
        ELSIF x =- 9322 THEN
            sigmoid_f := 21;
        ELSIF x =- 9321 THEN
            sigmoid_f := 21;
        ELSIF x =- 9320 THEN
            sigmoid_f := 21;
        ELSIF x =- 9319 THEN
            sigmoid_f := 21;
        ELSIF x =- 9318 THEN
            sigmoid_f := 21;
        ELSIF x =- 9317 THEN
            sigmoid_f := 21;
        ELSIF x =- 9316 THEN
            sigmoid_f := 21;
        ELSIF x =- 9315 THEN
            sigmoid_f := 21;
        ELSIF x =- 9314 THEN
            sigmoid_f := 21;
        ELSIF x =- 9313 THEN
            sigmoid_f := 21;
        ELSIF x =- 9312 THEN
            sigmoid_f := 21;
        ELSIF x =- 9311 THEN
            sigmoid_f := 21;
        ELSIF x =- 9310 THEN
            sigmoid_f := 21;
        ELSIF x =- 9309 THEN
            sigmoid_f := 21;
        ELSIF x =- 9308 THEN
            sigmoid_f := 21;
        ELSIF x =- 9307 THEN
            sigmoid_f := 21;
        ELSIF x =- 9306 THEN
            sigmoid_f := 21;
        ELSIF x =- 9305 THEN
            sigmoid_f := 21;
        ELSIF x =- 9304 THEN
            sigmoid_f := 21;
        ELSIF x =- 9303 THEN
            sigmoid_f := 21;
        ELSIF x =- 9302 THEN
            sigmoid_f := 21;
        ELSIF x =- 9301 THEN
            sigmoid_f := 21;
        ELSIF x =- 9300 THEN
            sigmoid_f := 21;
        ELSIF x =- 9299 THEN
            sigmoid_f := 21;
        ELSIF x =- 9298 THEN
            sigmoid_f := 21;
        ELSIF x =- 9297 THEN
            sigmoid_f := 21;
        ELSIF x =- 9296 THEN
            sigmoid_f := 21;
        ELSIF x =- 9295 THEN
            sigmoid_f := 21;
        ELSIF x =- 9294 THEN
            sigmoid_f := 21;
        ELSIF x =- 9293 THEN
            sigmoid_f := 21;
        ELSIF x =- 9292 THEN
            sigmoid_f := 21;
        ELSIF x =- 9291 THEN
            sigmoid_f := 21;
        ELSIF x =- 9290 THEN
            sigmoid_f := 21;
        ELSIF x =- 9289 THEN
            sigmoid_f := 21;
        ELSIF x =- 9288 THEN
            sigmoid_f := 21;
        ELSIF x =- 9287 THEN
            sigmoid_f := 21;
        ELSIF x =- 9286 THEN
            sigmoid_f := 21;
        ELSIF x =- 9285 THEN
            sigmoid_f := 21;
        ELSIF x =- 9284 THEN
            sigmoid_f := 21;
        ELSIF x =- 9283 THEN
            sigmoid_f := 21;
        ELSIF x =- 9282 THEN
            sigmoid_f := 21;
        ELSIF x =- 9281 THEN
            sigmoid_f := 21;
        ELSIF x =- 9280 THEN
            sigmoid_f := 21;
        ELSIF x =- 9279 THEN
            sigmoid_f := 21;
        ELSIF x =- 9278 THEN
            sigmoid_f := 21;
        ELSIF x =- 9277 THEN
            sigmoid_f := 21;
        ELSIF x =- 9276 THEN
            sigmoid_f := 21;
        ELSIF x =- 9275 THEN
            sigmoid_f := 21;
        ELSIF x =- 9274 THEN
            sigmoid_f := 21;
        ELSIF x =- 9273 THEN
            sigmoid_f := 21;
        ELSIF x =- 9272 THEN
            sigmoid_f := 21;
        ELSIF x =- 9271 THEN
            sigmoid_f := 21;
        ELSIF x =- 9270 THEN
            sigmoid_f := 21;
        ELSIF x =- 9269 THEN
            sigmoid_f := 21;
        ELSIF x =- 9268 THEN
            sigmoid_f := 21;
        ELSIF x =- 9267 THEN
            sigmoid_f := 21;
        ELSIF x =- 9266 THEN
            sigmoid_f := 21;
        ELSIF x =- 9265 THEN
            sigmoid_f := 21;
        ELSIF x =- 9264 THEN
            sigmoid_f := 22;
        ELSIF x =- 9263 THEN
            sigmoid_f := 22;
        ELSIF x =- 9262 THEN
            sigmoid_f := 22;
        ELSIF x =- 9261 THEN
            sigmoid_f := 22;
        ELSIF x =- 9260 THEN
            sigmoid_f := 22;
        ELSIF x =- 9259 THEN
            sigmoid_f := 22;
        ELSIF x =- 9258 THEN
            sigmoid_f := 22;
        ELSIF x =- 9257 THEN
            sigmoid_f := 22;
        ELSIF x =- 9256 THEN
            sigmoid_f := 22;
        ELSIF x =- 9255 THEN
            sigmoid_f := 22;
        ELSIF x =- 9254 THEN
            sigmoid_f := 22;
        ELSIF x =- 9253 THEN
            sigmoid_f := 22;
        ELSIF x =- 9252 THEN
            sigmoid_f := 22;
        ELSIF x =- 9251 THEN
            sigmoid_f := 22;
        ELSIF x =- 9250 THEN
            sigmoid_f := 22;
        ELSIF x =- 9249 THEN
            sigmoid_f := 22;
        ELSIF x =- 9248 THEN
            sigmoid_f := 22;
        ELSIF x =- 9247 THEN
            sigmoid_f := 22;
        ELSIF x =- 9246 THEN
            sigmoid_f := 22;
        ELSIF x =- 9245 THEN
            sigmoid_f := 22;
        ELSIF x =- 9244 THEN
            sigmoid_f := 22;
        ELSIF x =- 9243 THEN
            sigmoid_f := 22;
        ELSIF x =- 9242 THEN
            sigmoid_f := 22;
        ELSIF x =- 9241 THEN
            sigmoid_f := 22;
        ELSIF x =- 9240 THEN
            sigmoid_f := 22;
        ELSIF x =- 9239 THEN
            sigmoid_f := 22;
        ELSIF x =- 9238 THEN
            sigmoid_f := 22;
        ELSIF x =- 9237 THEN
            sigmoid_f := 22;
        ELSIF x =- 9236 THEN
            sigmoid_f := 22;
        ELSIF x =- 9235 THEN
            sigmoid_f := 22;
        ELSIF x =- 9234 THEN
            sigmoid_f := 22;
        ELSIF x =- 9233 THEN
            sigmoid_f := 22;
        ELSIF x =- 9232 THEN
            sigmoid_f := 22;
        ELSIF x =- 9231 THEN
            sigmoid_f := 22;
        ELSIF x =- 9230 THEN
            sigmoid_f := 22;
        ELSIF x =- 9229 THEN
            sigmoid_f := 22;
        ELSIF x =- 9228 THEN
            sigmoid_f := 22;
        ELSIF x =- 9227 THEN
            sigmoid_f := 22;
        ELSIF x =- 9226 THEN
            sigmoid_f := 22;
        ELSIF x =- 9225 THEN
            sigmoid_f := 22;
        ELSIF x =- 9224 THEN
            sigmoid_f := 22;
        ELSIF x =- 9223 THEN
            sigmoid_f := 22;
        ELSIF x =- 9222 THEN
            sigmoid_f := 22;
        ELSIF x =- 9221 THEN
            sigmoid_f := 22;
        ELSIF x =- 9220 THEN
            sigmoid_f := 22;
        ELSIF x =- 9219 THEN
            sigmoid_f := 22;
        ELSIF x =- 9218 THEN
            sigmoid_f := 22;
        ELSIF x =- 9217 THEN
            sigmoid_f := 22;
        ELSIF x =- 9216 THEN
            sigmoid_f := 22;
        ELSIF x =- 9215 THEN
            sigmoid_f := 22;
        ELSIF x =- 9214 THEN
            sigmoid_f := 22;
        ELSIF x =- 9213 THEN
            sigmoid_f := 22;
        ELSIF x =- 9212 THEN
            sigmoid_f := 22;
        ELSIF x =- 9211 THEN
            sigmoid_f := 22;
        ELSIF x =- 9210 THEN
            sigmoid_f := 22;
        ELSIF x =- 9209 THEN
            sigmoid_f := 22;
        ELSIF x =- 9208 THEN
            sigmoid_f := 22;
        ELSIF x =- 9207 THEN
            sigmoid_f := 22;
        ELSIF x =- 9206 THEN
            sigmoid_f := 22;
        ELSIF x =- 9205 THEN
            sigmoid_f := 22;
        ELSIF x =- 9204 THEN
            sigmoid_f := 22;
        ELSIF x =- 9203 THEN
            sigmoid_f := 22;
        ELSIF x =- 9202 THEN
            sigmoid_f := 22;
        ELSIF x =- 9201 THEN
            sigmoid_f := 22;
        ELSIF x =- 9200 THEN
            sigmoid_f := 22;
        ELSIF x =- 9199 THEN
            sigmoid_f := 22;
        ELSIF x =- 9198 THEN
            sigmoid_f := 22;
        ELSIF x =- 9197 THEN
            sigmoid_f := 22;
        ELSIF x =- 9196 THEN
            sigmoid_f := 22;
        ELSIF x =- 9195 THEN
            sigmoid_f := 22;
        ELSIF x =- 9194 THEN
            sigmoid_f := 22;
        ELSIF x =- 9193 THEN
            sigmoid_f := 22;
        ELSIF x =- 9192 THEN
            sigmoid_f := 22;
        ELSIF x =- 9191 THEN
            sigmoid_f := 22;
        ELSIF x =- 9190 THEN
            sigmoid_f := 22;
        ELSIF x =- 9189 THEN
            sigmoid_f := 22;
        ELSIF x =- 9188 THEN
            sigmoid_f := 22;
        ELSIF x =- 9187 THEN
            sigmoid_f := 22;
        ELSIF x =- 9186 THEN
            sigmoid_f := 22;
        ELSIF x =- 9185 THEN
            sigmoid_f := 22;
        ELSIF x =- 9184 THEN
            sigmoid_f := 22;
        ELSIF x =- 9183 THEN
            sigmoid_f := 22;
        ELSIF x =- 9182 THEN
            sigmoid_f := 22;
        ELSIF x =- 9181 THEN
            sigmoid_f := 22;
        ELSIF x =- 9180 THEN
            sigmoid_f := 22;
        ELSIF x =- 9179 THEN
            sigmoid_f := 22;
        ELSIF x =- 9178 THEN
            sigmoid_f := 22;
        ELSIF x =- 9177 THEN
            sigmoid_f := 22;
        ELSIF x =- 9176 THEN
            sigmoid_f := 22;
        ELSIF x =- 9175 THEN
            sigmoid_f := 23;
        ELSIF x =- 9174 THEN
            sigmoid_f := 23;
        ELSIF x =- 9173 THEN
            sigmoid_f := 23;
        ELSIF x =- 9172 THEN
            sigmoid_f := 23;
        ELSIF x =- 9171 THEN
            sigmoid_f := 23;
        ELSIF x =- 9170 THEN
            sigmoid_f := 23;
        ELSIF x =- 9169 THEN
            sigmoid_f := 23;
        ELSIF x =- 9168 THEN
            sigmoid_f := 23;
        ELSIF x =- 9167 THEN
            sigmoid_f := 23;
        ELSIF x =- 9166 THEN
            sigmoid_f := 23;
        ELSIF x =- 9165 THEN
            sigmoid_f := 23;
        ELSIF x =- 9164 THEN
            sigmoid_f := 23;
        ELSIF x =- 9163 THEN
            sigmoid_f := 23;
        ELSIF x =- 9162 THEN
            sigmoid_f := 23;
        ELSIF x =- 9161 THEN
            sigmoid_f := 23;
        ELSIF x =- 9160 THEN
            sigmoid_f := 23;
        ELSIF x =- 9159 THEN
            sigmoid_f := 23;
        ELSIF x =- 9158 THEN
            sigmoid_f := 23;
        ELSIF x =- 9157 THEN
            sigmoid_f := 23;
        ELSIF x =- 9156 THEN
            sigmoid_f := 23;
        ELSIF x =- 9155 THEN
            sigmoid_f := 23;
        ELSIF x =- 9154 THEN
            sigmoid_f := 23;
        ELSIF x =- 9153 THEN
            sigmoid_f := 23;
        ELSIF x =- 9152 THEN
            sigmoid_f := 23;
        ELSIF x =- 9151 THEN
            sigmoid_f := 23;
        ELSIF x =- 9150 THEN
            sigmoid_f := 23;
        ELSIF x =- 9149 THEN
            sigmoid_f := 23;
        ELSIF x =- 9148 THEN
            sigmoid_f := 23;
        ELSIF x =- 9147 THEN
            sigmoid_f := 23;
        ELSIF x =- 9146 THEN
            sigmoid_f := 23;
        ELSIF x =- 9145 THEN
            sigmoid_f := 23;
        ELSIF x =- 9144 THEN
            sigmoid_f := 23;
        ELSIF x =- 9143 THEN
            sigmoid_f := 23;
        ELSIF x =- 9142 THEN
            sigmoid_f := 23;
        ELSIF x =- 9141 THEN
            sigmoid_f := 23;
        ELSIF x =- 9140 THEN
            sigmoid_f := 23;
        ELSIF x =- 9139 THEN
            sigmoid_f := 23;
        ELSIF x =- 9138 THEN
            sigmoid_f := 23;
        ELSIF x =- 9137 THEN
            sigmoid_f := 23;
        ELSIF x =- 9136 THEN
            sigmoid_f := 23;
        ELSIF x =- 9135 THEN
            sigmoid_f := 23;
        ELSIF x =- 9134 THEN
            sigmoid_f := 23;
        ELSIF x =- 9133 THEN
            sigmoid_f := 23;
        ELSIF x =- 9132 THEN
            sigmoid_f := 23;
        ELSIF x =- 9131 THEN
            sigmoid_f := 23;
        ELSIF x =- 9130 THEN
            sigmoid_f := 23;
        ELSIF x =- 9129 THEN
            sigmoid_f := 23;
        ELSIF x =- 9128 THEN
            sigmoid_f := 23;
        ELSIF x =- 9127 THEN
            sigmoid_f := 23;
        ELSIF x =- 9126 THEN
            sigmoid_f := 23;
        ELSIF x =- 9125 THEN
            sigmoid_f := 23;
        ELSIF x =- 9124 THEN
            sigmoid_f := 23;
        ELSIF x =- 9123 THEN
            sigmoid_f := 23;
        ELSIF x =- 9122 THEN
            sigmoid_f := 23;
        ELSIF x =- 9121 THEN
            sigmoid_f := 23;
        ELSIF x =- 9120 THEN
            sigmoid_f := 23;
        ELSIF x =- 9119 THEN
            sigmoid_f := 23;
        ELSIF x =- 9118 THEN
            sigmoid_f := 23;
        ELSIF x =- 9117 THEN
            sigmoid_f := 23;
        ELSIF x =- 9116 THEN
            sigmoid_f := 23;
        ELSIF x =- 9115 THEN
            sigmoid_f := 23;
        ELSIF x =- 9114 THEN
            sigmoid_f := 23;
        ELSIF x =- 9113 THEN
            sigmoid_f := 23;
        ELSIF x =- 9112 THEN
            sigmoid_f := 23;
        ELSIF x =- 9111 THEN
            sigmoid_f := 23;
        ELSIF x =- 9110 THEN
            sigmoid_f := 23;
        ELSIF x =- 9109 THEN
            sigmoid_f := 23;
        ELSIF x =- 9108 THEN
            sigmoid_f := 23;
        ELSIF x =- 9107 THEN
            sigmoid_f := 23;
        ELSIF x =- 9106 THEN
            sigmoid_f := 23;
        ELSIF x =- 9105 THEN
            sigmoid_f := 23;
        ELSIF x =- 9104 THEN
            sigmoid_f := 23;
        ELSIF x =- 9103 THEN
            sigmoid_f := 23;
        ELSIF x =- 9102 THEN
            sigmoid_f := 23;
        ELSIF x =- 9101 THEN
            sigmoid_f := 23;
        ELSIF x =- 9100 THEN
            sigmoid_f := 23;
        ELSIF x =- 9099 THEN
            sigmoid_f := 23;
        ELSIF x =- 9098 THEN
            sigmoid_f := 23;
        ELSIF x =- 9097 THEN
            sigmoid_f := 23;
        ELSIF x =- 9096 THEN
            sigmoid_f := 23;
        ELSIF x =- 9095 THEN
            sigmoid_f := 23;
        ELSIF x =- 9094 THEN
            sigmoid_f := 23;
        ELSIF x =- 9093 THEN
            sigmoid_f := 24;
        ELSIF x =- 9092 THEN
            sigmoid_f := 24;
        ELSIF x =- 9091 THEN
            sigmoid_f := 24;
        ELSIF x =- 9090 THEN
            sigmoid_f := 24;
        ELSIF x =- 9089 THEN
            sigmoid_f := 24;
        ELSIF x =- 9088 THEN
            sigmoid_f := 24;
        ELSIF x =- 9087 THEN
            sigmoid_f := 24;
        ELSIF x =- 9086 THEN
            sigmoid_f := 24;
        ELSIF x =- 9085 THEN
            sigmoid_f := 24;
        ELSIF x =- 9084 THEN
            sigmoid_f := 24;
        ELSIF x =- 9083 THEN
            sigmoid_f := 24;
        ELSIF x =- 9082 THEN
            sigmoid_f := 24;
        ELSIF x =- 9081 THEN
            sigmoid_f := 24;
        ELSIF x =- 9080 THEN
            sigmoid_f := 24;
        ELSIF x =- 9079 THEN
            sigmoid_f := 24;
        ELSIF x =- 9078 THEN
            sigmoid_f := 24;
        ELSIF x =- 9077 THEN
            sigmoid_f := 24;
        ELSIF x =- 9076 THEN
            sigmoid_f := 24;
        ELSIF x =- 9075 THEN
            sigmoid_f := 24;
        ELSIF x =- 9074 THEN
            sigmoid_f := 24;
        ELSIF x =- 9073 THEN
            sigmoid_f := 24;
        ELSIF x =- 9072 THEN
            sigmoid_f := 24;
        ELSIF x =- 9071 THEN
            sigmoid_f := 24;
        ELSIF x =- 9070 THEN
            sigmoid_f := 24;
        ELSIF x =- 9069 THEN
            sigmoid_f := 24;
        ELSIF x =- 9068 THEN
            sigmoid_f := 24;
        ELSIF x =- 9067 THEN
            sigmoid_f := 24;
        ELSIF x =- 9066 THEN
            sigmoid_f := 24;
        ELSIF x =- 9065 THEN
            sigmoid_f := 24;
        ELSIF x =- 9064 THEN
            sigmoid_f := 24;
        ELSIF x =- 9063 THEN
            sigmoid_f := 24;
        ELSIF x =- 9062 THEN
            sigmoid_f := 24;
        ELSIF x =- 9061 THEN
            sigmoid_f := 24;
        ELSIF x =- 9060 THEN
            sigmoid_f := 24;
        ELSIF x =- 9059 THEN
            sigmoid_f := 24;
        ELSIF x =- 9058 THEN
            sigmoid_f := 24;
        ELSIF x =- 9057 THEN
            sigmoid_f := 24;
        ELSIF x =- 9056 THEN
            sigmoid_f := 24;
        ELSIF x =- 9055 THEN
            sigmoid_f := 24;
        ELSIF x =- 9054 THEN
            sigmoid_f := 24;
        ELSIF x =- 9053 THEN
            sigmoid_f := 24;
        ELSIF x =- 9052 THEN
            sigmoid_f := 24;
        ELSIF x =- 9051 THEN
            sigmoid_f := 24;
        ELSIF x =- 9050 THEN
            sigmoid_f := 24;
        ELSIF x =- 9049 THEN
            sigmoid_f := 24;
        ELSIF x =- 9048 THEN
            sigmoid_f := 24;
        ELSIF x =- 9047 THEN
            sigmoid_f := 24;
        ELSIF x =- 9046 THEN
            sigmoid_f := 24;
        ELSIF x =- 9045 THEN
            sigmoid_f := 24;
        ELSIF x =- 9044 THEN
            sigmoid_f := 24;
        ELSIF x =- 9043 THEN
            sigmoid_f := 24;
        ELSIF x =- 9042 THEN
            sigmoid_f := 24;
        ELSIF x =- 9041 THEN
            sigmoid_f := 24;
        ELSIF x =- 9040 THEN
            sigmoid_f := 24;
        ELSIF x =- 9039 THEN
            sigmoid_f := 24;
        ELSIF x =- 9038 THEN
            sigmoid_f := 24;
        ELSIF x =- 9037 THEN
            sigmoid_f := 24;
        ELSIF x =- 9036 THEN
            sigmoid_f := 24;
        ELSIF x =- 9035 THEN
            sigmoid_f := 24;
        ELSIF x =- 9034 THEN
            sigmoid_f := 24;
        ELSIF x =- 9033 THEN
            sigmoid_f := 24;
        ELSIF x =- 9032 THEN
            sigmoid_f := 24;
        ELSIF x =- 9031 THEN
            sigmoid_f := 24;
        ELSIF x =- 9030 THEN
            sigmoid_f := 24;
        ELSIF x =- 9029 THEN
            sigmoid_f := 24;
        ELSIF x =- 9028 THEN
            sigmoid_f := 24;
        ELSIF x =- 9027 THEN
            sigmoid_f := 24;
        ELSIF x =- 9026 THEN
            sigmoid_f := 24;
        ELSIF x =- 9025 THEN
            sigmoid_f := 24;
        ELSIF x =- 9024 THEN
            sigmoid_f := 24;
        ELSIF x =- 9023 THEN
            sigmoid_f := 24;
        ELSIF x =- 9022 THEN
            sigmoid_f := 24;
        ELSIF x =- 9021 THEN
            sigmoid_f := 24;
        ELSIF x =- 9020 THEN
            sigmoid_f := 24;
        ELSIF x =- 9019 THEN
            sigmoid_f := 24;
        ELSIF x =- 9018 THEN
            sigmoid_f := 24;
        ELSIF x =- 9017 THEN
            sigmoid_f := 24;
        ELSIF x =- 9016 THEN
            sigmoid_f := 24;
        ELSIF x =- 9015 THEN
            sigmoid_f := 24;
        ELSIF x =- 9014 THEN
            sigmoid_f := 24;
        ELSIF x =- 9013 THEN
            sigmoid_f := 24;
        ELSIF x =- 9012 THEN
            sigmoid_f := 24;
        ELSIF x =- 9011 THEN
            sigmoid_f := 25;
        ELSIF x =- 9010 THEN
            sigmoid_f := 25;
        ELSIF x =- 9009 THEN
            sigmoid_f := 25;
        ELSIF x =- 9008 THEN
            sigmoid_f := 25;
        ELSIF x =- 9007 THEN
            sigmoid_f := 25;
        ELSIF x =- 9006 THEN
            sigmoid_f := 25;
        ELSIF x =- 9005 THEN
            sigmoid_f := 25;
        ELSIF x =- 9004 THEN
            sigmoid_f := 25;
        ELSIF x =- 9003 THEN
            sigmoid_f := 25;
        ELSIF x =- 9002 THEN
            sigmoid_f := 25;
        ELSIF x =- 9001 THEN
            sigmoid_f := 25;
        ELSIF x =- 9000 THEN
            sigmoid_f := 25;
        ELSIF x =- 8999 THEN
            sigmoid_f := 25;
        ELSIF x =- 8998 THEN
            sigmoid_f := 25;
        ELSIF x =- 8997 THEN
            sigmoid_f := 25;
        ELSIF x =- 8996 THEN
            sigmoid_f := 25;
        ELSIF x =- 8995 THEN
            sigmoid_f := 25;
        ELSIF x =- 8994 THEN
            sigmoid_f := 25;
        ELSIF x =- 8993 THEN
            sigmoid_f := 25;
        ELSIF x =- 8992 THEN
            sigmoid_f := 25;
        ELSIF x =- 8991 THEN
            sigmoid_f := 25;
        ELSIF x =- 8990 THEN
            sigmoid_f := 25;
        ELSIF x =- 8989 THEN
            sigmoid_f := 25;
        ELSIF x =- 8988 THEN
            sigmoid_f := 25;
        ELSIF x =- 8987 THEN
            sigmoid_f := 25;
        ELSIF x =- 8986 THEN
            sigmoid_f := 25;
        ELSIF x =- 8985 THEN
            sigmoid_f := 25;
        ELSIF x =- 8984 THEN
            sigmoid_f := 25;
        ELSIF x =- 8983 THEN
            sigmoid_f := 25;
        ELSIF x =- 8982 THEN
            sigmoid_f := 25;
        ELSIF x =- 8981 THEN
            sigmoid_f := 25;
        ELSIF x =- 8980 THEN
            sigmoid_f := 25;
        ELSIF x =- 8979 THEN
            sigmoid_f := 25;
        ELSIF x =- 8978 THEN
            sigmoid_f := 25;
        ELSIF x =- 8977 THEN
            sigmoid_f := 25;
        ELSIF x =- 8976 THEN
            sigmoid_f := 25;
        ELSIF x =- 8975 THEN
            sigmoid_f := 25;
        ELSIF x =- 8974 THEN
            sigmoid_f := 25;
        ELSIF x =- 8973 THEN
            sigmoid_f := 25;
        ELSIF x =- 8972 THEN
            sigmoid_f := 25;
        ELSIF x =- 8971 THEN
            sigmoid_f := 25;
        ELSIF x =- 8970 THEN
            sigmoid_f := 25;
        ELSIF x =- 8969 THEN
            sigmoid_f := 25;
        ELSIF x =- 8968 THEN
            sigmoid_f := 25;
        ELSIF x =- 8967 THEN
            sigmoid_f := 25;
        ELSIF x =- 8966 THEN
            sigmoid_f := 25;
        ELSIF x =- 8965 THEN
            sigmoid_f := 25;
        ELSIF x =- 8964 THEN
            sigmoid_f := 25;
        ELSIF x =- 8963 THEN
            sigmoid_f := 25;
        ELSIF x =- 8962 THEN
            sigmoid_f := 25;
        ELSIF x =- 8961 THEN
            sigmoid_f := 25;
        ELSIF x =- 8960 THEN
            sigmoid_f := 25;
        ELSIF x =- 8959 THEN
            sigmoid_f := 25;
        ELSIF x =- 8958 THEN
            sigmoid_f := 25;
        ELSIF x =- 8957 THEN
            sigmoid_f := 25;
        ELSIF x =- 8956 THEN
            sigmoid_f := 25;
        ELSIF x =- 8955 THEN
            sigmoid_f := 25;
        ELSIF x =- 8954 THEN
            sigmoid_f := 25;
        ELSIF x =- 8953 THEN
            sigmoid_f := 25;
        ELSIF x =- 8952 THEN
            sigmoid_f := 25;
        ELSIF x =- 8951 THEN
            sigmoid_f := 25;
        ELSIF x =- 8950 THEN
            sigmoid_f := 25;
        ELSIF x =- 8949 THEN
            sigmoid_f := 25;
        ELSIF x =- 8948 THEN
            sigmoid_f := 25;
        ELSIF x =- 8947 THEN
            sigmoid_f := 25;
        ELSIF x =- 8946 THEN
            sigmoid_f := 25;
        ELSIF x =- 8945 THEN
            sigmoid_f := 25;
        ELSIF x =- 8944 THEN
            sigmoid_f := 25;
        ELSIF x =- 8943 THEN
            sigmoid_f := 25;
        ELSIF x =- 8942 THEN
            sigmoid_f := 25;
        ELSIF x =- 8941 THEN
            sigmoid_f := 25;
        ELSIF x =- 8940 THEN
            sigmoid_f := 25;
        ELSIF x =- 8939 THEN
            sigmoid_f := 25;
        ELSIF x =- 8938 THEN
            sigmoid_f := 25;
        ELSIF x =- 8937 THEN
            sigmoid_f := 25;
        ELSIF x =- 8936 THEN
            sigmoid_f := 25;
        ELSIF x =- 8935 THEN
            sigmoid_f := 25;
        ELSIF x =- 8934 THEN
            sigmoid_f := 25;
        ELSIF x =- 8933 THEN
            sigmoid_f := 25;
        ELSIF x =- 8932 THEN
            sigmoid_f := 25;
        ELSIF x =- 8931 THEN
            sigmoid_f := 25;
        ELSIF x =- 8930 THEN
            sigmoid_f := 25;
        ELSIF x =- 8929 THEN
            sigmoid_f := 26;
        ELSIF x =- 8928 THEN
            sigmoid_f := 26;
        ELSIF x =- 8927 THEN
            sigmoid_f := 26;
        ELSIF x =- 8926 THEN
            sigmoid_f := 26;
        ELSIF x =- 8925 THEN
            sigmoid_f := 26;
        ELSIF x =- 8924 THEN
            sigmoid_f := 26;
        ELSIF x =- 8923 THEN
            sigmoid_f := 26;
        ELSIF x =- 8922 THEN
            sigmoid_f := 26;
        ELSIF x =- 8921 THEN
            sigmoid_f := 26;
        ELSIF x =- 8920 THEN
            sigmoid_f := 26;
        ELSIF x =- 8919 THEN
            sigmoid_f := 26;
        ELSIF x =- 8918 THEN
            sigmoid_f := 26;
        ELSIF x =- 8917 THEN
            sigmoid_f := 26;
        ELSIF x =- 8916 THEN
            sigmoid_f := 26;
        ELSIF x =- 8915 THEN
            sigmoid_f := 26;
        ELSIF x =- 8914 THEN
            sigmoid_f := 26;
        ELSIF x =- 8913 THEN
            sigmoid_f := 26;
        ELSIF x =- 8912 THEN
            sigmoid_f := 26;
        ELSIF x =- 8911 THEN
            sigmoid_f := 26;
        ELSIF x =- 8910 THEN
            sigmoid_f := 26;
        ELSIF x =- 8909 THEN
            sigmoid_f := 26;
        ELSIF x =- 8908 THEN
            sigmoid_f := 26;
        ELSIF x =- 8907 THEN
            sigmoid_f := 26;
        ELSIF x =- 8906 THEN
            sigmoid_f := 26;
        ELSIF x =- 8905 THEN
            sigmoid_f := 26;
        ELSIF x =- 8904 THEN
            sigmoid_f := 26;
        ELSIF x =- 8903 THEN
            sigmoid_f := 26;
        ELSIF x =- 8902 THEN
            sigmoid_f := 26;
        ELSIF x =- 8901 THEN
            sigmoid_f := 26;
        ELSIF x =- 8900 THEN
            sigmoid_f := 26;
        ELSIF x =- 8899 THEN
            sigmoid_f := 26;
        ELSIF x =- 8898 THEN
            sigmoid_f := 26;
        ELSIF x =- 8897 THEN
            sigmoid_f := 26;
        ELSIF x =- 8896 THEN
            sigmoid_f := 26;
        ELSIF x =- 8895 THEN
            sigmoid_f := 26;
        ELSIF x =- 8894 THEN
            sigmoid_f := 26;
        ELSIF x =- 8893 THEN
            sigmoid_f := 26;
        ELSIF x =- 8892 THEN
            sigmoid_f := 26;
        ELSIF x =- 8891 THEN
            sigmoid_f := 26;
        ELSIF x =- 8890 THEN
            sigmoid_f := 26;
        ELSIF x =- 8889 THEN
            sigmoid_f := 26;
        ELSIF x =- 8888 THEN
            sigmoid_f := 26;
        ELSIF x =- 8887 THEN
            sigmoid_f := 26;
        ELSIF x =- 8886 THEN
            sigmoid_f := 26;
        ELSIF x =- 8885 THEN
            sigmoid_f := 26;
        ELSIF x =- 8884 THEN
            sigmoid_f := 26;
        ELSIF x =- 8883 THEN
            sigmoid_f := 26;
        ELSIF x =- 8882 THEN
            sigmoid_f := 26;
        ELSIF x =- 8881 THEN
            sigmoid_f := 26;
        ELSIF x =- 8880 THEN
            sigmoid_f := 26;
        ELSIF x =- 8879 THEN
            sigmoid_f := 26;
        ELSIF x =- 8878 THEN
            sigmoid_f := 26;
        ELSIF x =- 8877 THEN
            sigmoid_f := 26;
        ELSIF x =- 8876 THEN
            sigmoid_f := 26;
        ELSIF x =- 8875 THEN
            sigmoid_f := 26;
        ELSIF x =- 8874 THEN
            sigmoid_f := 26;
        ELSIF x =- 8873 THEN
            sigmoid_f := 26;
        ELSIF x =- 8872 THEN
            sigmoid_f := 26;
        ELSIF x =- 8871 THEN
            sigmoid_f := 26;
        ELSIF x =- 8870 THEN
            sigmoid_f := 26;
        ELSIF x =- 8869 THEN
            sigmoid_f := 26;
        ELSIF x =- 8868 THEN
            sigmoid_f := 26;
        ELSIF x =- 8867 THEN
            sigmoid_f := 26;
        ELSIF x =- 8866 THEN
            sigmoid_f := 26;
        ELSIF x =- 8865 THEN
            sigmoid_f := 26;
        ELSIF x =- 8864 THEN
            sigmoid_f := 26;
        ELSIF x =- 8863 THEN
            sigmoid_f := 26;
        ELSIF x =- 8862 THEN
            sigmoid_f := 26;
        ELSIF x =- 8861 THEN
            sigmoid_f := 26;
        ELSIF x =- 8860 THEN
            sigmoid_f := 26;
        ELSIF x =- 8859 THEN
            sigmoid_f := 26;
        ELSIF x =- 8858 THEN
            sigmoid_f := 26;
        ELSIF x =- 8857 THEN
            sigmoid_f := 26;
        ELSIF x =- 8856 THEN
            sigmoid_f := 26;
        ELSIF x =- 8855 THEN
            sigmoid_f := 26;
        ELSIF x =- 8854 THEN
            sigmoid_f := 26;
        ELSIF x =- 8853 THEN
            sigmoid_f := 26;
        ELSIF x =- 8852 THEN
            sigmoid_f := 26;
        ELSIF x =- 8851 THEN
            sigmoid_f := 26;
        ELSIF x =- 8850 THEN
            sigmoid_f := 26;
        ELSIF x =- 8849 THEN
            sigmoid_f := 26;
        ELSIF x =- 8848 THEN
            sigmoid_f := 26;
        ELSIF x =- 8847 THEN
            sigmoid_f := 27;
        ELSIF x =- 8846 THEN
            sigmoid_f := 27;
        ELSIF x =- 8845 THEN
            sigmoid_f := 27;
        ELSIF x =- 8844 THEN
            sigmoid_f := 27;
        ELSIF x =- 8843 THEN
            sigmoid_f := 27;
        ELSIF x =- 8842 THEN
            sigmoid_f := 27;
        ELSIF x =- 8841 THEN
            sigmoid_f := 27;
        ELSIF x =- 8840 THEN
            sigmoid_f := 27;
        ELSIF x =- 8839 THEN
            sigmoid_f := 27;
        ELSIF x =- 8838 THEN
            sigmoid_f := 27;
        ELSIF x =- 8837 THEN
            sigmoid_f := 27;
        ELSIF x =- 8836 THEN
            sigmoid_f := 27;
        ELSIF x =- 8835 THEN
            sigmoid_f := 27;
        ELSIF x =- 8834 THEN
            sigmoid_f := 27;
        ELSIF x =- 8833 THEN
            sigmoid_f := 27;
        ELSIF x =- 8832 THEN
            sigmoid_f := 27;
        ELSIF x =- 8831 THEN
            sigmoid_f := 27;
        ELSIF x =- 8830 THEN
            sigmoid_f := 27;
        ELSIF x =- 8829 THEN
            sigmoid_f := 27;
        ELSIF x =- 8828 THEN
            sigmoid_f := 27;
        ELSIF x =- 8827 THEN
            sigmoid_f := 27;
        ELSIF x =- 8826 THEN
            sigmoid_f := 27;
        ELSIF x =- 8825 THEN
            sigmoid_f := 27;
        ELSIF x =- 8824 THEN
            sigmoid_f := 27;
        ELSIF x =- 8823 THEN
            sigmoid_f := 27;
        ELSIF x =- 8822 THEN
            sigmoid_f := 27;
        ELSIF x =- 8821 THEN
            sigmoid_f := 27;
        ELSIF x =- 8820 THEN
            sigmoid_f := 27;
        ELSIF x =- 8819 THEN
            sigmoid_f := 27;
        ELSIF x =- 8818 THEN
            sigmoid_f := 27;
        ELSIF x =- 8817 THEN
            sigmoid_f := 27;
        ELSIF x =- 8816 THEN
            sigmoid_f := 27;
        ELSIF x =- 8815 THEN
            sigmoid_f := 27;
        ELSIF x =- 8814 THEN
            sigmoid_f := 27;
        ELSIF x =- 8813 THEN
            sigmoid_f := 27;
        ELSIF x =- 8812 THEN
            sigmoid_f := 27;
        ELSIF x =- 8811 THEN
            sigmoid_f := 27;
        ELSIF x =- 8810 THEN
            sigmoid_f := 27;
        ELSIF x =- 8809 THEN
            sigmoid_f := 27;
        ELSIF x =- 8808 THEN
            sigmoid_f := 27;
        ELSIF x =- 8807 THEN
            sigmoid_f := 27;
        ELSIF x =- 8806 THEN
            sigmoid_f := 27;
        ELSIF x =- 8805 THEN
            sigmoid_f := 27;
        ELSIF x =- 8804 THEN
            sigmoid_f := 27;
        ELSIF x =- 8803 THEN
            sigmoid_f := 27;
        ELSIF x =- 8802 THEN
            sigmoid_f := 27;
        ELSIF x =- 8801 THEN
            sigmoid_f := 27;
        ELSIF x =- 8800 THEN
            sigmoid_f := 27;
        ELSIF x =- 8799 THEN
            sigmoid_f := 27;
        ELSIF x =- 8798 THEN
            sigmoid_f := 27;
        ELSIF x =- 8797 THEN
            sigmoid_f := 27;
        ELSIF x =- 8796 THEN
            sigmoid_f := 27;
        ELSIF x =- 8795 THEN
            sigmoid_f := 27;
        ELSIF x =- 8794 THEN
            sigmoid_f := 27;
        ELSIF x =- 8793 THEN
            sigmoid_f := 27;
        ELSIF x =- 8792 THEN
            sigmoid_f := 27;
        ELSIF x =- 8791 THEN
            sigmoid_f := 27;
        ELSIF x =- 8790 THEN
            sigmoid_f := 27;
        ELSIF x =- 8789 THEN
            sigmoid_f := 27;
        ELSIF x =- 8788 THEN
            sigmoid_f := 27;
        ELSIF x =- 8787 THEN
            sigmoid_f := 27;
        ELSIF x =- 8786 THEN
            sigmoid_f := 27;
        ELSIF x =- 8785 THEN
            sigmoid_f := 27;
        ELSIF x =- 8784 THEN
            sigmoid_f := 27;
        ELSIF x =- 8783 THEN
            sigmoid_f := 27;
        ELSIF x =- 8782 THEN
            sigmoid_f := 27;
        ELSIF x =- 8781 THEN
            sigmoid_f := 27;
        ELSIF x =- 8780 THEN
            sigmoid_f := 27;
        ELSIF x =- 8779 THEN
            sigmoid_f := 27;
        ELSIF x =- 8778 THEN
            sigmoid_f := 27;
        ELSIF x =- 8777 THEN
            sigmoid_f := 27;
        ELSIF x =- 8776 THEN
            sigmoid_f := 27;
        ELSIF x =- 8775 THEN
            sigmoid_f := 27;
        ELSIF x =- 8774 THEN
            sigmoid_f := 27;
        ELSIF x =- 8773 THEN
            sigmoid_f := 27;
        ELSIF x =- 8772 THEN
            sigmoid_f := 27;
        ELSIF x =- 8771 THEN
            sigmoid_f := 27;
        ELSIF x =- 8770 THEN
            sigmoid_f := 27;
        ELSIF x =- 8769 THEN
            sigmoid_f := 27;
        ELSIF x =- 8768 THEN
            sigmoid_f := 27;
        ELSIF x =- 8767 THEN
            sigmoid_f := 27;
        ELSIF x =- 8766 THEN
            sigmoid_f := 27;
        ELSIF x =- 8765 THEN
            sigmoid_f := 28;
        ELSIF x =- 8764 THEN
            sigmoid_f := 28;
        ELSIF x =- 8763 THEN
            sigmoid_f := 28;
        ELSIF x =- 8762 THEN
            sigmoid_f := 28;
        ELSIF x =- 8761 THEN
            sigmoid_f := 28;
        ELSIF x =- 8760 THEN
            sigmoid_f := 28;
        ELSIF x =- 8759 THEN
            sigmoid_f := 28;
        ELSIF x =- 8758 THEN
            sigmoid_f := 28;
        ELSIF x =- 8757 THEN
            sigmoid_f := 28;
        ELSIF x =- 8756 THEN
            sigmoid_f := 28;
        ELSIF x =- 8755 THEN
            sigmoid_f := 28;
        ELSIF x =- 8754 THEN
            sigmoid_f := 28;
        ELSIF x =- 8753 THEN
            sigmoid_f := 28;
        ELSIF x =- 8752 THEN
            sigmoid_f := 28;
        ELSIF x =- 8751 THEN
            sigmoid_f := 28;
        ELSIF x =- 8750 THEN
            sigmoid_f := 28;
        ELSIF x =- 8749 THEN
            sigmoid_f := 28;
        ELSIF x =- 8748 THEN
            sigmoid_f := 28;
        ELSIF x =- 8747 THEN
            sigmoid_f := 28;
        ELSIF x =- 8746 THEN
            sigmoid_f := 28;
        ELSIF x =- 8745 THEN
            sigmoid_f := 28;
        ELSIF x =- 8744 THEN
            sigmoid_f := 28;
        ELSIF x =- 8743 THEN
            sigmoid_f := 28;
        ELSIF x =- 8742 THEN
            sigmoid_f := 28;
        ELSIF x =- 8741 THEN
            sigmoid_f := 28;
        ELSIF x =- 8740 THEN
            sigmoid_f := 28;
        ELSIF x =- 8739 THEN
            sigmoid_f := 28;
        ELSIF x =- 8738 THEN
            sigmoid_f := 28;
        ELSIF x =- 8737 THEN
            sigmoid_f := 28;
        ELSIF x =- 8736 THEN
            sigmoid_f := 28;
        ELSIF x =- 8735 THEN
            sigmoid_f := 28;
        ELSIF x =- 8734 THEN
            sigmoid_f := 28;
        ELSIF x =- 8733 THEN
            sigmoid_f := 28;
        ELSIF x =- 8732 THEN
            sigmoid_f := 28;
        ELSIF x =- 8731 THEN
            sigmoid_f := 28;
        ELSIF x =- 8730 THEN
            sigmoid_f := 28;
        ELSIF x =- 8729 THEN
            sigmoid_f := 28;
        ELSIF x =- 8728 THEN
            sigmoid_f := 28;
        ELSIF x =- 8727 THEN
            sigmoid_f := 28;
        ELSIF x =- 8726 THEN
            sigmoid_f := 28;
        ELSIF x =- 8725 THEN
            sigmoid_f := 28;
        ELSIF x =- 8724 THEN
            sigmoid_f := 28;
        ELSIF x =- 8723 THEN
            sigmoid_f := 28;
        ELSIF x =- 8722 THEN
            sigmoid_f := 28;
        ELSIF x =- 8721 THEN
            sigmoid_f := 28;
        ELSIF x =- 8720 THEN
            sigmoid_f := 28;
        ELSIF x =- 8719 THEN
            sigmoid_f := 28;
        ELSIF x =- 8718 THEN
            sigmoid_f := 28;
        ELSIF x =- 8717 THEN
            sigmoid_f := 28;
        ELSIF x =- 8716 THEN
            sigmoid_f := 28;
        ELSIF x =- 8715 THEN
            sigmoid_f := 28;
        ELSIF x =- 8714 THEN
            sigmoid_f := 28;
        ELSIF x =- 8713 THEN
            sigmoid_f := 28;
        ELSIF x =- 8712 THEN
            sigmoid_f := 28;
        ELSIF x =- 8711 THEN
            sigmoid_f := 28;
        ELSIF x =- 8710 THEN
            sigmoid_f := 28;
        ELSIF x =- 8709 THEN
            sigmoid_f := 28;
        ELSIF x =- 8708 THEN
            sigmoid_f := 28;
        ELSIF x =- 8707 THEN
            sigmoid_f := 28;
        ELSIF x =- 8706 THEN
            sigmoid_f := 28;
        ELSIF x =- 8705 THEN
            sigmoid_f := 28;
        ELSIF x =- 8704 THEN
            sigmoid_f := 28;
        ELSIF x =- 8703 THEN
            sigmoid_f := 28;
        ELSIF x =- 8702 THEN
            sigmoid_f := 28;
        ELSIF x =- 8701 THEN
            sigmoid_f := 28;
        ELSIF x =- 8700 THEN
            sigmoid_f := 28;
        ELSIF x =- 8699 THEN
            sigmoid_f := 28;
        ELSIF x =- 8698 THEN
            sigmoid_f := 28;
        ELSIF x =- 8697 THEN
            sigmoid_f := 28;
        ELSIF x =- 8696 THEN
            sigmoid_f := 28;
        ELSIF x =- 8695 THEN
            sigmoid_f := 28;
        ELSIF x =- 8694 THEN
            sigmoid_f := 28;
        ELSIF x =- 8693 THEN
            sigmoid_f := 28;
        ELSIF x =- 8692 THEN
            sigmoid_f := 28;
        ELSIF x =- 8691 THEN
            sigmoid_f := 28;
        ELSIF x =- 8690 THEN
            sigmoid_f := 28;
        ELSIF x =- 8689 THEN
            sigmoid_f := 28;
        ELSIF x =- 8688 THEN
            sigmoid_f := 28;
        ELSIF x =- 8687 THEN
            sigmoid_f := 28;
        ELSIF x =- 8686 THEN
            sigmoid_f := 28;
        ELSIF x =- 8685 THEN
            sigmoid_f := 28;
        ELSIF x =- 8684 THEN
            sigmoid_f := 28;
        ELSIF x =- 8683 THEN
            sigmoid_f := 28;
        ELSIF x =- 8682 THEN
            sigmoid_f := 28;
        ELSIF x =- 8681 THEN
            sigmoid_f := 28;
        ELSIF x =- 8680 THEN
            sigmoid_f := 28;
        ELSIF x =- 8679 THEN
            sigmoid_f := 28;
        ELSIF x =- 8678 THEN
            sigmoid_f := 28;
        ELSIF x =- 8677 THEN
            sigmoid_f := 28;
        ELSIF x =- 8676 THEN
            sigmoid_f := 28;
        ELSIF x =- 8675 THEN
            sigmoid_f := 28;
        ELSIF x =- 8674 THEN
            sigmoid_f := 28;
        ELSIF x =- 8673 THEN
            sigmoid_f := 29;
        ELSIF x =- 8672 THEN
            sigmoid_f := 29;
        ELSIF x =- 8671 THEN
            sigmoid_f := 29;
        ELSIF x =- 8670 THEN
            sigmoid_f := 29;
        ELSIF x =- 8669 THEN
            sigmoid_f := 29;
        ELSIF x =- 8668 THEN
            sigmoid_f := 29;
        ELSIF x =- 8667 THEN
            sigmoid_f := 29;
        ELSIF x =- 8666 THEN
            sigmoid_f := 29;
        ELSIF x =- 8665 THEN
            sigmoid_f := 29;
        ELSIF x =- 8664 THEN
            sigmoid_f := 29;
        ELSIF x =- 8663 THEN
            sigmoid_f := 29;
        ELSIF x =- 8662 THEN
            sigmoid_f := 29;
        ELSIF x =- 8661 THEN
            sigmoid_f := 29;
        ELSIF x =- 8660 THEN
            sigmoid_f := 29;
        ELSIF x =- 8659 THEN
            sigmoid_f := 29;
        ELSIF x =- 8658 THEN
            sigmoid_f := 29;
        ELSIF x =- 8657 THEN
            sigmoid_f := 29;
        ELSIF x =- 8656 THEN
            sigmoid_f := 29;
        ELSIF x =- 8655 THEN
            sigmoid_f := 29;
        ELSIF x =- 8654 THEN
            sigmoid_f := 29;
        ELSIF x =- 8653 THEN
            sigmoid_f := 29;
        ELSIF x =- 8652 THEN
            sigmoid_f := 29;
        ELSIF x =- 8651 THEN
            sigmoid_f := 29;
        ELSIF x =- 8650 THEN
            sigmoid_f := 29;
        ELSIF x =- 8649 THEN
            sigmoid_f := 29;
        ELSIF x =- 8648 THEN
            sigmoid_f := 29;
        ELSIF x =- 8647 THEN
            sigmoid_f := 29;
        ELSIF x =- 8646 THEN
            sigmoid_f := 29;
        ELSIF x =- 8645 THEN
            sigmoid_f := 29;
        ELSIF x =- 8644 THEN
            sigmoid_f := 29;
        ELSIF x =- 8643 THEN
            sigmoid_f := 29;
        ELSIF x =- 8642 THEN
            sigmoid_f := 29;
        ELSIF x =- 8641 THEN
            sigmoid_f := 29;
        ELSIF x =- 8640 THEN
            sigmoid_f := 29;
        ELSIF x =- 8639 THEN
            sigmoid_f := 29;
        ELSIF x =- 8638 THEN
            sigmoid_f := 29;
        ELSIF x =- 8637 THEN
            sigmoid_f := 29;
        ELSIF x =- 8636 THEN
            sigmoid_f := 29;
        ELSIF x =- 8635 THEN
            sigmoid_f := 29;
        ELSIF x =- 8634 THEN
            sigmoid_f := 29;
        ELSIF x =- 8633 THEN
            sigmoid_f := 29;
        ELSIF x =- 8632 THEN
            sigmoid_f := 29;
        ELSIF x =- 8631 THEN
            sigmoid_f := 29;
        ELSIF x =- 8630 THEN
            sigmoid_f := 29;
        ELSIF x =- 8629 THEN
            sigmoid_f := 29;
        ELSIF x =- 8628 THEN
            sigmoid_f := 29;
        ELSIF x =- 8627 THEN
            sigmoid_f := 29;
        ELSIF x =- 8626 THEN
            sigmoid_f := 29;
        ELSIF x =- 8625 THEN
            sigmoid_f := 29;
        ELSIF x =- 8624 THEN
            sigmoid_f := 29;
        ELSIF x =- 8623 THEN
            sigmoid_f := 29;
        ELSIF x =- 8622 THEN
            sigmoid_f := 29;
        ELSIF x =- 8621 THEN
            sigmoid_f := 29;
        ELSIF x =- 8620 THEN
            sigmoid_f := 29;
        ELSIF x =- 8619 THEN
            sigmoid_f := 29;
        ELSIF x =- 8618 THEN
            sigmoid_f := 29;
        ELSIF x =- 8617 THEN
            sigmoid_f := 29;
        ELSIF x =- 8616 THEN
            sigmoid_f := 29;
        ELSIF x =- 8615 THEN
            sigmoid_f := 29;
        ELSIF x =- 8614 THEN
            sigmoid_f := 29;
        ELSIF x =- 8613 THEN
            sigmoid_f := 30;
        ELSIF x =- 8612 THEN
            sigmoid_f := 30;
        ELSIF x =- 8611 THEN
            sigmoid_f := 30;
        ELSIF x =- 8610 THEN
            sigmoid_f := 30;
        ELSIF x =- 8609 THEN
            sigmoid_f := 30;
        ELSIF x =- 8608 THEN
            sigmoid_f := 30;
        ELSIF x =- 8607 THEN
            sigmoid_f := 30;
        ELSIF x =- 8606 THEN
            sigmoid_f := 30;
        ELSIF x =- 8605 THEN
            sigmoid_f := 30;
        ELSIF x =- 8604 THEN
            sigmoid_f := 30;
        ELSIF x =- 8603 THEN
            sigmoid_f := 30;
        ELSIF x =- 8602 THEN
            sigmoid_f := 30;
        ELSIF x =- 8601 THEN
            sigmoid_f := 30;
        ELSIF x =- 8600 THEN
            sigmoid_f := 30;
        ELSIF x =- 8599 THEN
            sigmoid_f := 30;
        ELSIF x =- 8598 THEN
            sigmoid_f := 30;
        ELSIF x =- 8597 THEN
            sigmoid_f := 30;
        ELSIF x =- 8596 THEN
            sigmoid_f := 30;
        ELSIF x =- 8595 THEN
            sigmoid_f := 30;
        ELSIF x =- 8594 THEN
            sigmoid_f := 30;
        ELSIF x =- 8593 THEN
            sigmoid_f := 30;
        ELSIF x =- 8592 THEN
            sigmoid_f := 30;
        ELSIF x =- 8591 THEN
            sigmoid_f := 30;
        ELSIF x =- 8590 THEN
            sigmoid_f := 30;
        ELSIF x =- 8589 THEN
            sigmoid_f := 30;
        ELSIF x =- 8588 THEN
            sigmoid_f := 30;
        ELSIF x =- 8587 THEN
            sigmoid_f := 30;
        ELSIF x =- 8586 THEN
            sigmoid_f := 30;
        ELSIF x =- 8585 THEN
            sigmoid_f := 30;
        ELSIF x =- 8584 THEN
            sigmoid_f := 30;
        ELSIF x =- 8583 THEN
            sigmoid_f := 30;
        ELSIF x =- 8582 THEN
            sigmoid_f := 30;
        ELSIF x =- 8581 THEN
            sigmoid_f := 30;
        ELSIF x =- 8580 THEN
            sigmoid_f := 30;
        ELSIF x =- 8579 THEN
            sigmoid_f := 30;
        ELSIF x =- 8578 THEN
            sigmoid_f := 30;
        ELSIF x =- 8577 THEN
            sigmoid_f := 30;
        ELSIF x =- 8576 THEN
            sigmoid_f := 30;
        ELSIF x =- 8575 THEN
            sigmoid_f := 30;
        ELSIF x =- 8574 THEN
            sigmoid_f := 30;
        ELSIF x =- 8573 THEN
            sigmoid_f := 30;
        ELSIF x =- 8572 THEN
            sigmoid_f := 30;
        ELSIF x =- 8571 THEN
            sigmoid_f := 30;
        ELSIF x =- 8570 THEN
            sigmoid_f := 30;
        ELSIF x =- 8569 THEN
            sigmoid_f := 30;
        ELSIF x =- 8568 THEN
            sigmoid_f := 30;
        ELSIF x =- 8567 THEN
            sigmoid_f := 30;
        ELSIF x =- 8566 THEN
            sigmoid_f := 30;
        ELSIF x =- 8565 THEN
            sigmoid_f := 30;
        ELSIF x =- 8564 THEN
            sigmoid_f := 30;
        ELSIF x =- 8563 THEN
            sigmoid_f := 30;
        ELSIF x =- 8562 THEN
            sigmoid_f := 30;
        ELSIF x =- 8561 THEN
            sigmoid_f := 30;
        ELSIF x =- 8560 THEN
            sigmoid_f := 30;
        ELSIF x =- 8559 THEN
            sigmoid_f := 30;
        ELSIF x =- 8558 THEN
            sigmoid_f := 30;
        ELSIF x =- 8557 THEN
            sigmoid_f := 30;
        ELSIF x =- 8556 THEN
            sigmoid_f := 30;
        ELSIF x =- 8555 THEN
            sigmoid_f := 30;
        ELSIF x =- 8554 THEN
            sigmoid_f := 30;
        ELSIF x =- 8553 THEN
            sigmoid_f := 31;
        ELSIF x =- 8552 THEN
            sigmoid_f := 31;
        ELSIF x =- 8551 THEN
            sigmoid_f := 31;
        ELSIF x =- 8550 THEN
            sigmoid_f := 31;
        ELSIF x =- 8549 THEN
            sigmoid_f := 31;
        ELSIF x =- 8548 THEN
            sigmoid_f := 31;
        ELSIF x =- 8547 THEN
            sigmoid_f := 31;
        ELSIF x =- 8546 THEN
            sigmoid_f := 31;
        ELSIF x =- 8545 THEN
            sigmoid_f := 31;
        ELSIF x =- 8544 THEN
            sigmoid_f := 31;
        ELSIF x =- 8543 THEN
            sigmoid_f := 31;
        ELSIF x =- 8542 THEN
            sigmoid_f := 31;
        ELSIF x =- 8541 THEN
            sigmoid_f := 31;
        ELSIF x =- 8540 THEN
            sigmoid_f := 31;
        ELSIF x =- 8539 THEN
            sigmoid_f := 31;
        ELSIF x =- 8538 THEN
            sigmoid_f := 31;
        ELSIF x =- 8537 THEN
            sigmoid_f := 31;
        ELSIF x =- 8536 THEN
            sigmoid_f := 31;
        ELSIF x =- 8535 THEN
            sigmoid_f := 31;
        ELSIF x =- 8534 THEN
            sigmoid_f := 31;
        ELSIF x =- 8533 THEN
            sigmoid_f := 31;
        ELSIF x =- 8532 THEN
            sigmoid_f := 31;
        ELSIF x =- 8531 THEN
            sigmoid_f := 31;
        ELSIF x =- 8530 THEN
            sigmoid_f := 31;
        ELSIF x =- 8529 THEN
            sigmoid_f := 31;
        ELSIF x =- 8528 THEN
            sigmoid_f := 31;
        ELSIF x =- 8527 THEN
            sigmoid_f := 31;
        ELSIF x =- 8526 THEN
            sigmoid_f := 31;
        ELSIF x =- 8525 THEN
            sigmoid_f := 31;
        ELSIF x =- 8524 THEN
            sigmoid_f := 31;
        ELSIF x =- 8523 THEN
            sigmoid_f := 31;
        ELSIF x =- 8522 THEN
            sigmoid_f := 31;
        ELSIF x =- 8521 THEN
            sigmoid_f := 31;
        ELSIF x =- 8520 THEN
            sigmoid_f := 31;
        ELSIF x =- 8519 THEN
            sigmoid_f := 31;
        ELSIF x =- 8518 THEN
            sigmoid_f := 31;
        ELSIF x =- 8517 THEN
            sigmoid_f := 31;
        ELSIF x =- 8516 THEN
            sigmoid_f := 31;
        ELSIF x =- 8515 THEN
            sigmoid_f := 31;
        ELSIF x =- 8514 THEN
            sigmoid_f := 31;
        ELSIF x =- 8513 THEN
            sigmoid_f := 31;
        ELSIF x =- 8512 THEN
            sigmoid_f := 31;
        ELSIF x =- 8511 THEN
            sigmoid_f := 31;
        ELSIF x =- 8510 THEN
            sigmoid_f := 31;
        ELSIF x =- 8509 THEN
            sigmoid_f := 31;
        ELSIF x =- 8508 THEN
            sigmoid_f := 31;
        ELSIF x =- 8507 THEN
            sigmoid_f := 31;
        ELSIF x =- 8506 THEN
            sigmoid_f := 31;
        ELSIF x =- 8505 THEN
            sigmoid_f := 31;
        ELSIF x =- 8504 THEN
            sigmoid_f := 31;
        ELSIF x =- 8503 THEN
            sigmoid_f := 31;
        ELSIF x =- 8502 THEN
            sigmoid_f := 31;
        ELSIF x =- 8501 THEN
            sigmoid_f := 31;
        ELSIF x =- 8500 THEN
            sigmoid_f := 31;
        ELSIF x =- 8499 THEN
            sigmoid_f := 31;
        ELSIF x =- 8498 THEN
            sigmoid_f := 31;
        ELSIF x =- 8497 THEN
            sigmoid_f := 31;
        ELSIF x =- 8496 THEN
            sigmoid_f := 31;
        ELSIF x =- 8495 THEN
            sigmoid_f := 31;
        ELSIF x =- 8494 THEN
            sigmoid_f := 31;
        ELSIF x =- 8493 THEN
            sigmoid_f := 32;
        ELSIF x =- 8492 THEN
            sigmoid_f := 32;
        ELSIF x =- 8491 THEN
            sigmoid_f := 32;
        ELSIF x =- 8490 THEN
            sigmoid_f := 32;
        ELSIF x =- 8489 THEN
            sigmoid_f := 32;
        ELSIF x =- 8488 THEN
            sigmoid_f := 32;
        ELSIF x =- 8487 THEN
            sigmoid_f := 32;
        ELSIF x =- 8486 THEN
            sigmoid_f := 32;
        ELSIF x =- 8485 THEN
            sigmoid_f := 32;
        ELSIF x =- 8484 THEN
            sigmoid_f := 32;
        ELSIF x =- 8483 THEN
            sigmoid_f := 32;
        ELSIF x =- 8482 THEN
            sigmoid_f := 32;
        ELSIF x =- 8481 THEN
            sigmoid_f := 32;
        ELSIF x =- 8480 THEN
            sigmoid_f := 32;
        ELSIF x =- 8479 THEN
            sigmoid_f := 32;
        ELSIF x =- 8478 THEN
            sigmoid_f := 32;
        ELSIF x =- 8477 THEN
            sigmoid_f := 32;
        ELSIF x =- 8476 THEN
            sigmoid_f := 32;
        ELSIF x =- 8475 THEN
            sigmoid_f := 32;
        ELSIF x =- 8474 THEN
            sigmoid_f := 32;
        ELSIF x =- 8473 THEN
            sigmoid_f := 32;
        ELSIF x =- 8472 THEN
            sigmoid_f := 32;
        ELSIF x =- 8471 THEN
            sigmoid_f := 32;
        ELSIF x =- 8470 THEN
            sigmoid_f := 32;
        ELSIF x =- 8469 THEN
            sigmoid_f := 32;
        ELSIF x =- 8468 THEN
            sigmoid_f := 32;
        ELSIF x =- 8467 THEN
            sigmoid_f := 32;
        ELSIF x =- 8466 THEN
            sigmoid_f := 32;
        ELSIF x =- 8465 THEN
            sigmoid_f := 32;
        ELSIF x =- 8464 THEN
            sigmoid_f := 32;
        ELSIF x =- 8463 THEN
            sigmoid_f := 32;
        ELSIF x =- 8462 THEN
            sigmoid_f := 32;
        ELSIF x =- 8461 THEN
            sigmoid_f := 32;
        ELSIF x =- 8460 THEN
            sigmoid_f := 32;
        ELSIF x =- 8459 THEN
            sigmoid_f := 32;
        ELSIF x =- 8458 THEN
            sigmoid_f := 32;
        ELSIF x =- 8457 THEN
            sigmoid_f := 32;
        ELSIF x =- 8456 THEN
            sigmoid_f := 32;
        ELSIF x =- 8455 THEN
            sigmoid_f := 32;
        ELSIF x =- 8454 THEN
            sigmoid_f := 32;
        ELSIF x =- 8453 THEN
            sigmoid_f := 32;
        ELSIF x =- 8452 THEN
            sigmoid_f := 32;
        ELSIF x =- 8451 THEN
            sigmoid_f := 32;
        ELSIF x =- 8450 THEN
            sigmoid_f := 32;
        ELSIF x =- 8449 THEN
            sigmoid_f := 32;
        ELSIF x =- 8448 THEN
            sigmoid_f := 32;
        ELSIF x =- 8447 THEN
            sigmoid_f := 32;
        ELSIF x =- 8446 THEN
            sigmoid_f := 32;
        ELSIF x =- 8445 THEN
            sigmoid_f := 32;
        ELSIF x =- 8444 THEN
            sigmoid_f := 32;
        ELSIF x =- 8443 THEN
            sigmoid_f := 32;
        ELSIF x =- 8442 THEN
            sigmoid_f := 32;
        ELSIF x =- 8441 THEN
            sigmoid_f := 32;
        ELSIF x =- 8440 THEN
            sigmoid_f := 32;
        ELSIF x =- 8439 THEN
            sigmoid_f := 32;
        ELSIF x =- 8438 THEN
            sigmoid_f := 32;
        ELSIF x =- 8437 THEN
            sigmoid_f := 32;
        ELSIF x =- 8436 THEN
            sigmoid_f := 32;
        ELSIF x =- 8435 THEN
            sigmoid_f := 32;
        ELSIF x =- 8434 THEN
            sigmoid_f := 32;
        ELSIF x =- 8433 THEN
            sigmoid_f := 32;
        ELSIF x =- 8432 THEN
            sigmoid_f := 33;
        ELSIF x =- 8431 THEN
            sigmoid_f := 33;
        ELSIF x =- 8430 THEN
            sigmoid_f := 33;
        ELSIF x =- 8429 THEN
            sigmoid_f := 33;
        ELSIF x =- 8428 THEN
            sigmoid_f := 33;
        ELSIF x =- 8427 THEN
            sigmoid_f := 33;
        ELSIF x =- 8426 THEN
            sigmoid_f := 33;
        ELSIF x =- 8425 THEN
            sigmoid_f := 33;
        ELSIF x =- 8424 THEN
            sigmoid_f := 33;
        ELSIF x =- 8423 THEN
            sigmoid_f := 33;
        ELSIF x =- 8422 THEN
            sigmoid_f := 33;
        ELSIF x =- 8421 THEN
            sigmoid_f := 33;
        ELSIF x =- 8420 THEN
            sigmoid_f := 33;
        ELSIF x =- 8419 THEN
            sigmoid_f := 33;
        ELSIF x =- 8418 THEN
            sigmoid_f := 33;
        ELSIF x =- 8417 THEN
            sigmoid_f := 33;
        ELSIF x =- 8416 THEN
            sigmoid_f := 33;
        ELSIF x =- 8415 THEN
            sigmoid_f := 33;
        ELSIF x =- 8414 THEN
            sigmoid_f := 33;
        ELSIF x =- 8413 THEN
            sigmoid_f := 33;
        ELSIF x =- 8412 THEN
            sigmoid_f := 33;
        ELSIF x =- 8411 THEN
            sigmoid_f := 33;
        ELSIF x =- 8410 THEN
            sigmoid_f := 33;
        ELSIF x =- 8409 THEN
            sigmoid_f := 33;
        ELSIF x =- 8408 THEN
            sigmoid_f := 33;
        ELSIF x =- 8407 THEN
            sigmoid_f := 33;
        ELSIF x =- 8406 THEN
            sigmoid_f := 33;
        ELSIF x =- 8405 THEN
            sigmoid_f := 33;
        ELSIF x =- 8404 THEN
            sigmoid_f := 33;
        ELSIF x =- 8403 THEN
            sigmoid_f := 33;
        ELSIF x =- 8402 THEN
            sigmoid_f := 33;
        ELSIF x =- 8401 THEN
            sigmoid_f := 33;
        ELSIF x =- 8400 THEN
            sigmoid_f := 33;
        ELSIF x =- 8399 THEN
            sigmoid_f := 33;
        ELSIF x =- 8398 THEN
            sigmoid_f := 33;
        ELSIF x =- 8397 THEN
            sigmoid_f := 33;
        ELSIF x =- 8396 THEN
            sigmoid_f := 33;
        ELSIF x =- 8395 THEN
            sigmoid_f := 33;
        ELSIF x =- 8394 THEN
            sigmoid_f := 33;
        ELSIF x =- 8393 THEN
            sigmoid_f := 33;
        ELSIF x =- 8392 THEN
            sigmoid_f := 33;
        ELSIF x =- 8391 THEN
            sigmoid_f := 33;
        ELSIF x =- 8390 THEN
            sigmoid_f := 33;
        ELSIF x =- 8389 THEN
            sigmoid_f := 33;
        ELSIF x =- 8388 THEN
            sigmoid_f := 33;
        ELSIF x =- 8387 THEN
            sigmoid_f := 33;
        ELSIF x =- 8386 THEN
            sigmoid_f := 33;
        ELSIF x =- 8385 THEN
            sigmoid_f := 33;
        ELSIF x =- 8384 THEN
            sigmoid_f := 33;
        ELSIF x =- 8383 THEN
            sigmoid_f := 33;
        ELSIF x =- 8382 THEN
            sigmoid_f := 33;
        ELSIF x =- 8381 THEN
            sigmoid_f := 33;
        ELSIF x =- 8380 THEN
            sigmoid_f := 33;
        ELSIF x =- 8379 THEN
            sigmoid_f := 33;
        ELSIF x =- 8378 THEN
            sigmoid_f := 33;
        ELSIF x =- 8377 THEN
            sigmoid_f := 33;
        ELSIF x =- 8376 THEN
            sigmoid_f := 33;
        ELSIF x =- 8375 THEN
            sigmoid_f := 33;
        ELSIF x =- 8374 THEN
            sigmoid_f := 33;
        ELSIF x =- 8373 THEN
            sigmoid_f := 33;
        ELSIF x =- 8372 THEN
            sigmoid_f := 34;
        ELSIF x =- 8371 THEN
            sigmoid_f := 34;
        ELSIF x =- 8370 THEN
            sigmoid_f := 34;
        ELSIF x =- 8369 THEN
            sigmoid_f := 34;
        ELSIF x =- 8368 THEN
            sigmoid_f := 34;
        ELSIF x =- 8367 THEN
            sigmoid_f := 34;
        ELSIF x =- 8366 THEN
            sigmoid_f := 34;
        ELSIF x =- 8365 THEN
            sigmoid_f := 34;
        ELSIF x =- 8364 THEN
            sigmoid_f := 34;
        ELSIF x =- 8363 THEN
            sigmoid_f := 34;
        ELSIF x =- 8362 THEN
            sigmoid_f := 34;
        ELSIF x =- 8361 THEN
            sigmoid_f := 34;
        ELSIF x =- 8360 THEN
            sigmoid_f := 34;
        ELSIF x =- 8359 THEN
            sigmoid_f := 34;
        ELSIF x =- 8358 THEN
            sigmoid_f := 34;
        ELSIF x =- 8357 THEN
            sigmoid_f := 34;
        ELSIF x =- 8356 THEN
            sigmoid_f := 34;
        ELSIF x =- 8355 THEN
            sigmoid_f := 34;
        ELSIF x =- 8354 THEN
            sigmoid_f := 34;
        ELSIF x =- 8353 THEN
            sigmoid_f := 34;
        ELSIF x =- 8352 THEN
            sigmoid_f := 34;
        ELSIF x =- 8351 THEN
            sigmoid_f := 34;
        ELSIF x =- 8350 THEN
            sigmoid_f := 34;
        ELSIF x =- 8349 THEN
            sigmoid_f := 34;
        ELSIF x =- 8348 THEN
            sigmoid_f := 34;
        ELSIF x =- 8347 THEN
            sigmoid_f := 34;
        ELSIF x =- 8346 THEN
            sigmoid_f := 34;
        ELSIF x =- 8345 THEN
            sigmoid_f := 34;
        ELSIF x =- 8344 THEN
            sigmoid_f := 34;
        ELSIF x =- 8343 THEN
            sigmoid_f := 34;
        ELSIF x =- 8342 THEN
            sigmoid_f := 34;
        ELSIF x =- 8341 THEN
            sigmoid_f := 34;
        ELSIF x =- 8340 THEN
            sigmoid_f := 34;
        ELSIF x =- 8339 THEN
            sigmoid_f := 34;
        ELSIF x =- 8338 THEN
            sigmoid_f := 34;
        ELSIF x =- 8337 THEN
            sigmoid_f := 34;
        ELSIF x =- 8336 THEN
            sigmoid_f := 34;
        ELSIF x =- 8335 THEN
            sigmoid_f := 34;
        ELSIF x =- 8334 THEN
            sigmoid_f := 34;
        ELSIF x =- 8333 THEN
            sigmoid_f := 34;
        ELSIF x =- 8332 THEN
            sigmoid_f := 34;
        ELSIF x =- 8331 THEN
            sigmoid_f := 34;
        ELSIF x =- 8330 THEN
            sigmoid_f := 34;
        ELSIF x =- 8329 THEN
            sigmoid_f := 34;
        ELSIF x =- 8328 THEN
            sigmoid_f := 34;
        ELSIF x =- 8327 THEN
            sigmoid_f := 34;
        ELSIF x =- 8326 THEN
            sigmoid_f := 34;
        ELSIF x =- 8325 THEN
            sigmoid_f := 34;
        ELSIF x =- 8324 THEN
            sigmoid_f := 34;
        ELSIF x =- 8323 THEN
            sigmoid_f := 34;
        ELSIF x =- 8322 THEN
            sigmoid_f := 34;
        ELSIF x =- 8321 THEN
            sigmoid_f := 34;
        ELSIF x =- 8320 THEN
            sigmoid_f := 34;
        ELSIF x =- 8319 THEN
            sigmoid_f := 34;
        ELSIF x =- 8318 THEN
            sigmoid_f := 34;
        ELSIF x =- 8317 THEN
            sigmoid_f := 34;
        ELSIF x =- 8316 THEN
            sigmoid_f := 34;
        ELSIF x =- 8315 THEN
            sigmoid_f := 34;
        ELSIF x =- 8314 THEN
            sigmoid_f := 34;
        ELSIF x =- 8313 THEN
            sigmoid_f := 34;
        ELSIF x =- 8312 THEN
            sigmoid_f := 35;
        ELSIF x =- 8311 THEN
            sigmoid_f := 35;
        ELSIF x =- 8310 THEN
            sigmoid_f := 35;
        ELSIF x =- 8309 THEN
            sigmoid_f := 35;
        ELSIF x =- 8308 THEN
            sigmoid_f := 35;
        ELSIF x =- 8307 THEN
            sigmoid_f := 35;
        ELSIF x =- 8306 THEN
            sigmoid_f := 35;
        ELSIF x =- 8305 THEN
            sigmoid_f := 35;
        ELSIF x =- 8304 THEN
            sigmoid_f := 35;
        ELSIF x =- 8303 THEN
            sigmoid_f := 35;
        ELSIF x =- 8302 THEN
            sigmoid_f := 35;
        ELSIF x =- 8301 THEN
            sigmoid_f := 35;
        ELSIF x =- 8300 THEN
            sigmoid_f := 35;
        ELSIF x =- 8299 THEN
            sigmoid_f := 35;
        ELSIF x =- 8298 THEN
            sigmoid_f := 35;
        ELSIF x =- 8297 THEN
            sigmoid_f := 35;
        ELSIF x =- 8296 THEN
            sigmoid_f := 35;
        ELSIF x =- 8295 THEN
            sigmoid_f := 35;
        ELSIF x =- 8294 THEN
            sigmoid_f := 35;
        ELSIF x =- 8293 THEN
            sigmoid_f := 35;
        ELSIF x =- 8292 THEN
            sigmoid_f := 35;
        ELSIF x =- 8291 THEN
            sigmoid_f := 35;
        ELSIF x =- 8290 THEN
            sigmoid_f := 35;
        ELSIF x =- 8289 THEN
            sigmoid_f := 35;
        ELSIF x =- 8288 THEN
            sigmoid_f := 35;
        ELSIF x =- 8287 THEN
            sigmoid_f := 35;
        ELSIF x =- 8286 THEN
            sigmoid_f := 35;
        ELSIF x =- 8285 THEN
            sigmoid_f := 35;
        ELSIF x =- 8284 THEN
            sigmoid_f := 35;
        ELSIF x =- 8283 THEN
            sigmoid_f := 35;
        ELSIF x =- 8282 THEN
            sigmoid_f := 35;
        ELSIF x =- 8281 THEN
            sigmoid_f := 35;
        ELSIF x =- 8280 THEN
            sigmoid_f := 35;
        ELSIF x =- 8279 THEN
            sigmoid_f := 35;
        ELSIF x =- 8278 THEN
            sigmoid_f := 35;
        ELSIF x =- 8277 THEN
            sigmoid_f := 35;
        ELSIF x =- 8276 THEN
            sigmoid_f := 35;
        ELSIF x =- 8275 THEN
            sigmoid_f := 35;
        ELSIF x =- 8274 THEN
            sigmoid_f := 35;
        ELSIF x =- 8273 THEN
            sigmoid_f := 35;
        ELSIF x =- 8272 THEN
            sigmoid_f := 35;
        ELSIF x =- 8271 THEN
            sigmoid_f := 35;
        ELSIF x =- 8270 THEN
            sigmoid_f := 35;
        ELSIF x =- 8269 THEN
            sigmoid_f := 35;
        ELSIF x =- 8268 THEN
            sigmoid_f := 35;
        ELSIF x =- 8267 THEN
            sigmoid_f := 35;
        ELSIF x =- 8266 THEN
            sigmoid_f := 35;
        ELSIF x =- 8265 THEN
            sigmoid_f := 35;
        ELSIF x =- 8264 THEN
            sigmoid_f := 35;
        ELSIF x =- 8263 THEN
            sigmoid_f := 35;
        ELSIF x =- 8262 THEN
            sigmoid_f := 35;
        ELSIF x =- 8261 THEN
            sigmoid_f := 35;
        ELSIF x =- 8260 THEN
            sigmoid_f := 35;
        ELSIF x =- 8259 THEN
            sigmoid_f := 35;
        ELSIF x =- 8258 THEN
            sigmoid_f := 35;
        ELSIF x =- 8257 THEN
            sigmoid_f := 35;
        ELSIF x =- 8256 THEN
            sigmoid_f := 35;
        ELSIF x =- 8255 THEN
            sigmoid_f := 35;
        ELSIF x =- 8254 THEN
            sigmoid_f := 35;
        ELSIF x =- 8253 THEN
            sigmoid_f := 35;
        ELSIF x =- 8252 THEN
            sigmoid_f := 36;
        ELSIF x =- 8251 THEN
            sigmoid_f := 36;
        ELSIF x =- 8250 THEN
            sigmoid_f := 36;
        ELSIF x =- 8249 THEN
            sigmoid_f := 36;
        ELSIF x =- 8248 THEN
            sigmoid_f := 36;
        ELSIF x =- 8247 THEN
            sigmoid_f := 36;
        ELSIF x =- 8246 THEN
            sigmoid_f := 36;
        ELSIF x =- 8245 THEN
            sigmoid_f := 36;
        ELSIF x =- 8244 THEN
            sigmoid_f := 36;
        ELSIF x =- 8243 THEN
            sigmoid_f := 36;
        ELSIF x =- 8242 THEN
            sigmoid_f := 36;
        ELSIF x =- 8241 THEN
            sigmoid_f := 36;
        ELSIF x =- 8240 THEN
            sigmoid_f := 36;
        ELSIF x =- 8239 THEN
            sigmoid_f := 36;
        ELSIF x =- 8238 THEN
            sigmoid_f := 36;
        ELSIF x =- 8237 THEN
            sigmoid_f := 36;
        ELSIF x =- 8236 THEN
            sigmoid_f := 36;
        ELSIF x =- 8235 THEN
            sigmoid_f := 36;
        ELSIF x =- 8234 THEN
            sigmoid_f := 36;
        ELSIF x =- 8233 THEN
            sigmoid_f := 36;
        ELSIF x =- 8232 THEN
            sigmoid_f := 36;
        ELSIF x =- 8231 THEN
            sigmoid_f := 36;
        ELSIF x =- 8230 THEN
            sigmoid_f := 36;
        ELSIF x =- 8229 THEN
            sigmoid_f := 36;
        ELSIF x =- 8228 THEN
            sigmoid_f := 36;
        ELSIF x =- 8227 THEN
            sigmoid_f := 36;
        ELSIF x =- 8226 THEN
            sigmoid_f := 36;
        ELSIF x =- 8225 THEN
            sigmoid_f := 36;
        ELSIF x =- 8224 THEN
            sigmoid_f := 36;
        ELSIF x =- 8223 THEN
            sigmoid_f := 36;
        ELSIF x =- 8222 THEN
            sigmoid_f := 36;
        ELSIF x =- 8221 THEN
            sigmoid_f := 36;
        ELSIF x =- 8220 THEN
            sigmoid_f := 36;
        ELSIF x =- 8219 THEN
            sigmoid_f := 36;
        ELSIF x =- 8218 THEN
            sigmoid_f := 36;
        ELSIF x =- 8217 THEN
            sigmoid_f := 36;
        ELSIF x =- 8216 THEN
            sigmoid_f := 36;
        ELSIF x =- 8215 THEN
            sigmoid_f := 36;
        ELSIF x =- 8214 THEN
            sigmoid_f := 36;
        ELSIF x =- 8213 THEN
            sigmoid_f := 36;
        ELSIF x =- 8212 THEN
            sigmoid_f := 36;
        ELSIF x =- 8211 THEN
            sigmoid_f := 36;
        ELSIF x =- 8210 THEN
            sigmoid_f := 36;
        ELSIF x =- 8209 THEN
            sigmoid_f := 36;
        ELSIF x =- 8208 THEN
            sigmoid_f := 36;
        ELSIF x =- 8207 THEN
            sigmoid_f := 36;
        ELSIF x =- 8206 THEN
            sigmoid_f := 36;
        ELSIF x =- 8205 THEN
            sigmoid_f := 36;
        ELSIF x =- 8204 THEN
            sigmoid_f := 36;
        ELSIF x =- 8203 THEN
            sigmoid_f := 36;
        ELSIF x =- 8202 THEN
            sigmoid_f := 36;
        ELSIF x =- 8201 THEN
            sigmoid_f := 36;
        ELSIF x =- 8200 THEN
            sigmoid_f := 36;
        ELSIF x =- 8199 THEN
            sigmoid_f := 36;
        ELSIF x =- 8198 THEN
            sigmoid_f := 36;
        ELSIF x =- 8197 THEN
            sigmoid_f := 36;
        ELSIF x =- 8196 THEN
            sigmoid_f := 36;
        ELSIF x =- 8195 THEN
            sigmoid_f := 36;
        ELSIF x =- 8194 THEN
            sigmoid_f := 36;
        ELSIF x =- 8193 THEN
            sigmoid_f := 36;
        ELSIF x =- 8192 THEN
            sigmoid_f := 37;
        ELSIF x =- 8191 THEN
            sigmoid_f := 37;
        ELSIF x =- 8190 THEN
            sigmoid_f := 37;
        ELSIF x =- 8189 THEN
            sigmoid_f := 37;
        ELSIF x =- 8188 THEN
            sigmoid_f := 37;
        ELSIF x =- 8187 THEN
            sigmoid_f := 37;
        ELSIF x =- 8186 THEN
            sigmoid_f := 37;
        ELSIF x =- 8185 THEN
            sigmoid_f := 37;
        ELSIF x =- 8184 THEN
            sigmoid_f := 37;
        ELSIF x =- 8183 THEN
            sigmoid_f := 37;
        ELSIF x =- 8182 THEN
            sigmoid_f := 37;
        ELSIF x =- 8181 THEN
            sigmoid_f := 37;
        ELSIF x =- 8180 THEN
            sigmoid_f := 37;
        ELSIF x =- 8179 THEN
            sigmoid_f := 37;
        ELSIF x =- 8178 THEN
            sigmoid_f := 37;
        ELSIF x =- 8177 THEN
            sigmoid_f := 37;
        ELSIF x =- 8176 THEN
            sigmoid_f := 37;
        ELSIF x =- 8175 THEN
            sigmoid_f := 37;
        ELSIF x =- 8174 THEN
            sigmoid_f := 37;
        ELSIF x =- 8173 THEN
            sigmoid_f := 37;
        ELSIF x =- 8172 THEN
            sigmoid_f := 37;
        ELSIF x =- 8171 THEN
            sigmoid_f := 37;
        ELSIF x =- 8170 THEN
            sigmoid_f := 37;
        ELSIF x =- 8169 THEN
            sigmoid_f := 37;
        ELSIF x =- 8168 THEN
            sigmoid_f := 37;
        ELSIF x =- 8167 THEN
            sigmoid_f := 37;
        ELSIF x =- 8166 THEN
            sigmoid_f := 37;
        ELSIF x =- 8165 THEN
            sigmoid_f := 37;
        ELSIF x =- 8164 THEN
            sigmoid_f := 37;
        ELSIF x =- 8163 THEN
            sigmoid_f := 37;
        ELSIF x =- 8162 THEN
            sigmoid_f := 37;
        ELSIF x =- 8161 THEN
            sigmoid_f := 37;
        ELSIF x =- 8160 THEN
            sigmoid_f := 37;
        ELSIF x =- 8159 THEN
            sigmoid_f := 37;
        ELSIF x =- 8158 THEN
            sigmoid_f := 37;
        ELSIF x =- 8157 THEN
            sigmoid_f := 37;
        ELSIF x =- 8156 THEN
            sigmoid_f := 37;
        ELSIF x =- 8155 THEN
            sigmoid_f := 37;
        ELSIF x =- 8154 THEN
            sigmoid_f := 37;
        ELSIF x =- 8153 THEN
            sigmoid_f := 37;
        ELSIF x =- 8152 THEN
            sigmoid_f := 37;
        ELSIF x =- 8151 THEN
            sigmoid_f := 37;
        ELSIF x =- 8150 THEN
            sigmoid_f := 37;
        ELSIF x =- 8149 THEN
            sigmoid_f := 37;
        ELSIF x =- 8148 THEN
            sigmoid_f := 37;
        ELSIF x =- 8147 THEN
            sigmoid_f := 37;
        ELSIF x =- 8146 THEN
            sigmoid_f := 37;
        ELSIF x =- 8145 THEN
            sigmoid_f := 37;
        ELSIF x =- 8144 THEN
            sigmoid_f := 37;
        ELSIF x =- 8143 THEN
            sigmoid_f := 37;
        ELSIF x =- 8142 THEN
            sigmoid_f := 37;
        ELSIF x =- 8141 THEN
            sigmoid_f := 37;
        ELSIF x =- 8140 THEN
            sigmoid_f := 37;
        ELSIF x =- 8139 THEN
            sigmoid_f := 38;
        ELSIF x =- 8138 THEN
            sigmoid_f := 38;
        ELSIF x =- 8137 THEN
            sigmoid_f := 38;
        ELSIF x =- 8136 THEN
            sigmoid_f := 38;
        ELSIF x =- 8135 THEN
            sigmoid_f := 38;
        ELSIF x =- 8134 THEN
            sigmoid_f := 38;
        ELSIF x =- 8133 THEN
            sigmoid_f := 38;
        ELSIF x =- 8132 THEN
            sigmoid_f := 38;
        ELSIF x =- 8131 THEN
            sigmoid_f := 38;
        ELSIF x =- 8130 THEN
            sigmoid_f := 38;
        ELSIF x =- 8129 THEN
            sigmoid_f := 38;
        ELSIF x =- 8128 THEN
            sigmoid_f := 38;
        ELSIF x =- 8127 THEN
            sigmoid_f := 38;
        ELSIF x =- 8126 THEN
            sigmoid_f := 38;
        ELSIF x =- 8125 THEN
            sigmoid_f := 38;
        ELSIF x =- 8124 THEN
            sigmoid_f := 38;
        ELSIF x =- 8123 THEN
            sigmoid_f := 38;
        ELSIF x =- 8122 THEN
            sigmoid_f := 38;
        ELSIF x =- 8121 THEN
            sigmoid_f := 38;
        ELSIF x =- 8120 THEN
            sigmoid_f := 38;
        ELSIF x =- 8119 THEN
            sigmoid_f := 38;
        ELSIF x =- 8118 THEN
            sigmoid_f := 38;
        ELSIF x =- 8117 THEN
            sigmoid_f := 38;
        ELSIF x =- 8116 THEN
            sigmoid_f := 38;
        ELSIF x =- 8115 THEN
            sigmoid_f := 38;
        ELSIF x =- 8114 THEN
            sigmoid_f := 38;
        ELSIF x =- 8113 THEN
            sigmoid_f := 38;
        ELSIF x =- 8112 THEN
            sigmoid_f := 38;
        ELSIF x =- 8111 THEN
            sigmoid_f := 38;
        ELSIF x =- 8110 THEN
            sigmoid_f := 38;
        ELSIF x =- 8109 THEN
            sigmoid_f := 38;
        ELSIF x =- 8108 THEN
            sigmoid_f := 38;
        ELSIF x =- 8107 THEN
            sigmoid_f := 38;
        ELSIF x =- 8106 THEN
            sigmoid_f := 38;
        ELSIF x =- 8105 THEN
            sigmoid_f := 38;
        ELSIF x =- 8104 THEN
            sigmoid_f := 38;
        ELSIF x =- 8103 THEN
            sigmoid_f := 38;
        ELSIF x =- 8102 THEN
            sigmoid_f := 38;
        ELSIF x =- 8101 THEN
            sigmoid_f := 38;
        ELSIF x =- 8100 THEN
            sigmoid_f := 38;
        ELSIF x =- 8099 THEN
            sigmoid_f := 38;
        ELSIF x =- 8098 THEN
            sigmoid_f := 38;
        ELSIF x =- 8097 THEN
            sigmoid_f := 38;
        ELSIF x =- 8096 THEN
            sigmoid_f := 38;
        ELSIF x =- 8095 THEN
            sigmoid_f := 38;
        ELSIF x =- 8094 THEN
            sigmoid_f := 38;
        ELSIF x =- 8093 THEN
            sigmoid_f := 38;
        ELSIF x =- 8092 THEN
            sigmoid_f := 38;
        ELSIF x =- 8091 THEN
            sigmoid_f := 38;
        ELSIF x =- 8090 THEN
            sigmoid_f := 38;
        ELSIF x =- 8089 THEN
            sigmoid_f := 38;
        ELSIF x =- 8088 THEN
            sigmoid_f := 38;
        ELSIF x =- 8087 THEN
            sigmoid_f := 38;
        ELSIF x =- 8086 THEN
            sigmoid_f := 39;
        ELSIF x =- 8085 THEN
            sigmoid_f := 39;
        ELSIF x =- 8084 THEN
            sigmoid_f := 39;
        ELSIF x =- 8083 THEN
            sigmoid_f := 39;
        ELSIF x =- 8082 THEN
            sigmoid_f := 39;
        ELSIF x =- 8081 THEN
            sigmoid_f := 39;
        ELSIF x =- 8080 THEN
            sigmoid_f := 39;
        ELSIF x =- 8079 THEN
            sigmoid_f := 39;
        ELSIF x =- 8078 THEN
            sigmoid_f := 39;
        ELSIF x =- 8077 THEN
            sigmoid_f := 39;
        ELSIF x =- 8076 THEN
            sigmoid_f := 39;
        ELSIF x =- 8075 THEN
            sigmoid_f := 39;
        ELSIF x =- 8074 THEN
            sigmoid_f := 39;
        ELSIF x =- 8073 THEN
            sigmoid_f := 39;
        ELSIF x =- 8072 THEN
            sigmoid_f := 39;
        ELSIF x =- 8071 THEN
            sigmoid_f := 39;
        ELSIF x =- 8070 THEN
            sigmoid_f := 39;
        ELSIF x =- 8069 THEN
            sigmoid_f := 39;
        ELSIF x =- 8068 THEN
            sigmoid_f := 39;
        ELSIF x =- 8067 THEN
            sigmoid_f := 39;
        ELSIF x =- 8066 THEN
            sigmoid_f := 39;
        ELSIF x =- 8065 THEN
            sigmoid_f := 39;
        ELSIF x =- 8064 THEN
            sigmoid_f := 39;
        ELSIF x =- 8063 THEN
            sigmoid_f := 39;
        ELSIF x =- 8062 THEN
            sigmoid_f := 39;
        ELSIF x =- 8061 THEN
            sigmoid_f := 39;
        ELSIF x =- 8060 THEN
            sigmoid_f := 39;
        ELSIF x =- 8059 THEN
            sigmoid_f := 39;
        ELSIF x =- 8058 THEN
            sigmoid_f := 39;
        ELSIF x =- 8057 THEN
            sigmoid_f := 39;
        ELSIF x =- 8056 THEN
            sigmoid_f := 39;
        ELSIF x =- 8055 THEN
            sigmoid_f := 39;
        ELSIF x =- 8054 THEN
            sigmoid_f := 39;
        ELSIF x =- 8053 THEN
            sigmoid_f := 39;
        ELSIF x =- 8052 THEN
            sigmoid_f := 39;
        ELSIF x =- 8051 THEN
            sigmoid_f := 39;
        ELSIF x =- 8050 THEN
            sigmoid_f := 39;
        ELSIF x =- 8049 THEN
            sigmoid_f := 39;
        ELSIF x =- 8048 THEN
            sigmoid_f := 39;
        ELSIF x =- 8047 THEN
            sigmoid_f := 39;
        ELSIF x =- 8046 THEN
            sigmoid_f := 39;
        ELSIF x =- 8045 THEN
            sigmoid_f := 39;
        ELSIF x =- 8044 THEN
            sigmoid_f := 39;
        ELSIF x =- 8043 THEN
            sigmoid_f := 39;
        ELSIF x =- 8042 THEN
            sigmoid_f := 39;
        ELSIF x =- 8041 THEN
            sigmoid_f := 39;
        ELSIF x =- 8040 THEN
            sigmoid_f := 39;
        ELSIF x =- 8039 THEN
            sigmoid_f := 39;
        ELSIF x =- 8038 THEN
            sigmoid_f := 39;
        ELSIF x =- 8037 THEN
            sigmoid_f := 39;
        ELSIF x =- 8036 THEN
            sigmoid_f := 39;
        ELSIF x =- 8035 THEN
            sigmoid_f := 39;
        ELSIF x =- 8034 THEN
            sigmoid_f := 40;
        ELSIF x =- 8033 THEN
            sigmoid_f := 40;
        ELSIF x =- 8032 THEN
            sigmoid_f := 40;
        ELSIF x =- 8031 THEN
            sigmoid_f := 40;
        ELSIF x =- 8030 THEN
            sigmoid_f := 40;
        ELSIF x =- 8029 THEN
            sigmoid_f := 40;
        ELSIF x =- 8028 THEN
            sigmoid_f := 40;
        ELSIF x =- 8027 THEN
            sigmoid_f := 40;
        ELSIF x =- 8026 THEN
            sigmoid_f := 40;
        ELSIF x =- 8025 THEN
            sigmoid_f := 40;
        ELSIF x =- 8024 THEN
            sigmoid_f := 40;
        ELSIF x =- 8023 THEN
            sigmoid_f := 40;
        ELSIF x =- 8022 THEN
            sigmoid_f := 40;
        ELSIF x =- 8021 THEN
            sigmoid_f := 40;
        ELSIF x =- 8020 THEN
            sigmoid_f := 40;
        ELSIF x =- 8019 THEN
            sigmoid_f := 40;
        ELSIF x =- 8018 THEN
            sigmoid_f := 40;
        ELSIF x =- 8017 THEN
            sigmoid_f := 40;
        ELSIF x =- 8016 THEN
            sigmoid_f := 40;
        ELSIF x =- 8015 THEN
            sigmoid_f := 40;
        ELSIF x =- 8014 THEN
            sigmoid_f := 40;
        ELSIF x =- 8013 THEN
            sigmoid_f := 40;
        ELSIF x =- 8012 THEN
            sigmoid_f := 40;
        ELSIF x =- 8011 THEN
            sigmoid_f := 40;
        ELSIF x =- 8010 THEN
            sigmoid_f := 40;
        ELSIF x =- 8009 THEN
            sigmoid_f := 40;
        ELSIF x =- 8008 THEN
            sigmoid_f := 40;
        ELSIF x =- 8007 THEN
            sigmoid_f := 40;
        ELSIF x =- 8006 THEN
            sigmoid_f := 40;
        ELSIF x =- 8005 THEN
            sigmoid_f := 40;
        ELSIF x =- 8004 THEN
            sigmoid_f := 40;
        ELSIF x =- 8003 THEN
            sigmoid_f := 40;
        ELSIF x =- 8002 THEN
            sigmoid_f := 40;
        ELSIF x =- 8001 THEN
            sigmoid_f := 40;
        ELSIF x =- 8000 THEN
            sigmoid_f := 40;
        ELSIF x =- 7999 THEN
            sigmoid_f := 40;
        ELSIF x =- 7998 THEN
            sigmoid_f := 40;
        ELSIF x =- 7997 THEN
            sigmoid_f := 40;
        ELSIF x =- 7996 THEN
            sigmoid_f := 40;
        ELSIF x =- 7995 THEN
            sigmoid_f := 40;
        ELSIF x =- 7994 THEN
            sigmoid_f := 40;
        ELSIF x =- 7993 THEN
            sigmoid_f := 40;
        ELSIF x =- 7992 THEN
            sigmoid_f := 40;
        ELSIF x =- 7991 THEN
            sigmoid_f := 40;
        ELSIF x =- 7990 THEN
            sigmoid_f := 40;
        ELSIF x =- 7989 THEN
            sigmoid_f := 40;
        ELSIF x =- 7988 THEN
            sigmoid_f := 40;
        ELSIF x =- 7987 THEN
            sigmoid_f := 40;
        ELSIF x =- 7986 THEN
            sigmoid_f := 40;
        ELSIF x =- 7985 THEN
            sigmoid_f := 40;
        ELSIF x =- 7984 THEN
            sigmoid_f := 40;
        ELSIF x =- 7983 THEN
            sigmoid_f := 40;
        ELSIF x =- 7982 THEN
            sigmoid_f := 40;
        ELSIF x =- 7981 THEN
            sigmoid_f := 41;
        ELSIF x =- 7980 THEN
            sigmoid_f := 41;
        ELSIF x =- 7979 THEN
            sigmoid_f := 41;
        ELSIF x =- 7978 THEN
            sigmoid_f := 41;
        ELSIF x =- 7977 THEN
            sigmoid_f := 41;
        ELSIF x =- 7976 THEN
            sigmoid_f := 41;
        ELSIF x =- 7975 THEN
            sigmoid_f := 41;
        ELSIF x =- 7974 THEN
            sigmoid_f := 41;
        ELSIF x =- 7973 THEN
            sigmoid_f := 41;
        ELSIF x =- 7972 THEN
            sigmoid_f := 41;
        ELSIF x =- 7971 THEN
            sigmoid_f := 41;
        ELSIF x =- 7970 THEN
            sigmoid_f := 41;
        ELSIF x =- 7969 THEN
            sigmoid_f := 41;
        ELSIF x =- 7968 THEN
            sigmoid_f := 41;
        ELSIF x =- 7967 THEN
            sigmoid_f := 41;
        ELSIF x =- 7966 THEN
            sigmoid_f := 41;
        ELSIF x =- 7965 THEN
            sigmoid_f := 41;
        ELSIF x =- 7964 THEN
            sigmoid_f := 41;
        ELSIF x =- 7963 THEN
            sigmoid_f := 41;
        ELSIF x =- 7962 THEN
            sigmoid_f := 41;
        ELSIF x =- 7961 THEN
            sigmoid_f := 41;
        ELSIF x =- 7960 THEN
            sigmoid_f := 41;
        ELSIF x =- 7959 THEN
            sigmoid_f := 41;
        ELSIF x =- 7958 THEN
            sigmoid_f := 41;
        ELSIF x =- 7957 THEN
            sigmoid_f := 41;
        ELSIF x =- 7956 THEN
            sigmoid_f := 41;
        ELSIF x =- 7955 THEN
            sigmoid_f := 41;
        ELSIF x =- 7954 THEN
            sigmoid_f := 41;
        ELSIF x =- 7953 THEN
            sigmoid_f := 41;
        ELSIF x =- 7952 THEN
            sigmoid_f := 41;
        ELSIF x =- 7951 THEN
            sigmoid_f := 41;
        ELSIF x =- 7950 THEN
            sigmoid_f := 41;
        ELSIF x =- 7949 THEN
            sigmoid_f := 41;
        ELSIF x =- 7948 THEN
            sigmoid_f := 41;
        ELSIF x =- 7947 THEN
            sigmoid_f := 41;
        ELSIF x =- 7946 THEN
            sigmoid_f := 41;
        ELSIF x =- 7945 THEN
            sigmoid_f := 41;
        ELSIF x =- 7944 THEN
            sigmoid_f := 41;
        ELSIF x =- 7943 THEN
            sigmoid_f := 41;
        ELSIF x =- 7942 THEN
            sigmoid_f := 41;
        ELSIF x =- 7941 THEN
            sigmoid_f := 41;
        ELSIF x =- 7940 THEN
            sigmoid_f := 41;
        ELSIF x =- 7939 THEN
            sigmoid_f := 41;
        ELSIF x =- 7938 THEN
            sigmoid_f := 41;
        ELSIF x =- 7937 THEN
            sigmoid_f := 41;
        ELSIF x =- 7936 THEN
            sigmoid_f := 41;
        ELSIF x =- 7935 THEN
            sigmoid_f := 41;
        ELSIF x =- 7934 THEN
            sigmoid_f := 41;
        ELSIF x =- 7933 THEN
            sigmoid_f := 41;
        ELSIF x =- 7932 THEN
            sigmoid_f := 41;
        ELSIF x =- 7931 THEN
            sigmoid_f := 41;
        ELSIF x =- 7930 THEN
            sigmoid_f := 41;
        ELSIF x =- 7929 THEN
            sigmoid_f := 42;
        ELSIF x =- 7928 THEN
            sigmoid_f := 42;
        ELSIF x =- 7927 THEN
            sigmoid_f := 42;
        ELSIF x =- 7926 THEN
            sigmoid_f := 42;
        ELSIF x =- 7925 THEN
            sigmoid_f := 42;
        ELSIF x =- 7924 THEN
            sigmoid_f := 42;
        ELSIF x =- 7923 THEN
            sigmoid_f := 42;
        ELSIF x =- 7922 THEN
            sigmoid_f := 42;
        ELSIF x =- 7921 THEN
            sigmoid_f := 42;
        ELSIF x =- 7920 THEN
            sigmoid_f := 42;
        ELSIF x =- 7919 THEN
            sigmoid_f := 42;
        ELSIF x =- 7918 THEN
            sigmoid_f := 42;
        ELSIF x =- 7917 THEN
            sigmoid_f := 42;
        ELSIF x =- 7916 THEN
            sigmoid_f := 42;
        ELSIF x =- 7915 THEN
            sigmoid_f := 42;
        ELSIF x =- 7914 THEN
            sigmoid_f := 42;
        ELSIF x =- 7913 THEN
            sigmoid_f := 42;
        ELSIF x =- 7912 THEN
            sigmoid_f := 42;
        ELSIF x =- 7911 THEN
            sigmoid_f := 42;
        ELSIF x =- 7910 THEN
            sigmoid_f := 42;
        ELSIF x =- 7909 THEN
            sigmoid_f := 42;
        ELSIF x =- 7908 THEN
            sigmoid_f := 42;
        ELSIF x =- 7907 THEN
            sigmoid_f := 42;
        ELSIF x =- 7906 THEN
            sigmoid_f := 42;
        ELSIF x =- 7905 THEN
            sigmoid_f := 42;
        ELSIF x =- 7904 THEN
            sigmoid_f := 42;
        ELSIF x =- 7903 THEN
            sigmoid_f := 42;
        ELSIF x =- 7902 THEN
            sigmoid_f := 42;
        ELSIF x =- 7901 THEN
            sigmoid_f := 42;
        ELSIF x =- 7900 THEN
            sigmoid_f := 42;
        ELSIF x =- 7899 THEN
            sigmoid_f := 42;
        ELSIF x =- 7898 THEN
            sigmoid_f := 42;
        ELSIF x =- 7897 THEN
            sigmoid_f := 42;
        ELSIF x =- 7896 THEN
            sigmoid_f := 42;
        ELSIF x =- 7895 THEN
            sigmoid_f := 42;
        ELSIF x =- 7894 THEN
            sigmoid_f := 42;
        ELSIF x =- 7893 THEN
            sigmoid_f := 42;
        ELSIF x =- 7892 THEN
            sigmoid_f := 42;
        ELSIF x =- 7891 THEN
            sigmoid_f := 42;
        ELSIF x =- 7890 THEN
            sigmoid_f := 42;
        ELSIF x =- 7889 THEN
            sigmoid_f := 42;
        ELSIF x =- 7888 THEN
            sigmoid_f := 42;
        ELSIF x =- 7887 THEN
            sigmoid_f := 42;
        ELSIF x =- 7886 THEN
            sigmoid_f := 42;
        ELSIF x =- 7885 THEN
            sigmoid_f := 42;
        ELSIF x =- 7884 THEN
            sigmoid_f := 42;
        ELSIF x =- 7883 THEN
            sigmoid_f := 42;
        ELSIF x =- 7882 THEN
            sigmoid_f := 42;
        ELSIF x =- 7881 THEN
            sigmoid_f := 42;
        ELSIF x =- 7880 THEN
            sigmoid_f := 42;
        ELSIF x =- 7879 THEN
            sigmoid_f := 42;
        ELSIF x =- 7878 THEN
            sigmoid_f := 42;
        ELSIF x =- 7877 THEN
            sigmoid_f := 42;
        ELSIF x =- 7876 THEN
            sigmoid_f := 43;
        ELSIF x =- 7875 THEN
            sigmoid_f := 43;
        ELSIF x =- 7874 THEN
            sigmoid_f := 43;
        ELSIF x =- 7873 THEN
            sigmoid_f := 43;
        ELSIF x =- 7872 THEN
            sigmoid_f := 43;
        ELSIF x =- 7871 THEN
            sigmoid_f := 43;
        ELSIF x =- 7870 THEN
            sigmoid_f := 43;
        ELSIF x =- 7869 THEN
            sigmoid_f := 43;
        ELSIF x =- 7868 THEN
            sigmoid_f := 43;
        ELSIF x =- 7867 THEN
            sigmoid_f := 43;
        ELSIF x =- 7866 THEN
            sigmoid_f := 43;
        ELSIF x =- 7865 THEN
            sigmoid_f := 43;
        ELSIF x =- 7864 THEN
            sigmoid_f := 43;
        ELSIF x =- 7863 THEN
            sigmoid_f := 43;
        ELSIF x =- 7862 THEN
            sigmoid_f := 43;
        ELSIF x =- 7861 THEN
            sigmoid_f := 43;
        ELSIF x =- 7860 THEN
            sigmoid_f := 43;
        ELSIF x =- 7859 THEN
            sigmoid_f := 43;
        ELSIF x =- 7858 THEN
            sigmoid_f := 43;
        ELSIF x =- 7857 THEN
            sigmoid_f := 43;
        ELSIF x =- 7856 THEN
            sigmoid_f := 43;
        ELSIF x =- 7855 THEN
            sigmoid_f := 43;
        ELSIF x =- 7854 THEN
            sigmoid_f := 43;
        ELSIF x =- 7853 THEN
            sigmoid_f := 43;
        ELSIF x =- 7852 THEN
            sigmoid_f := 43;
        ELSIF x =- 7851 THEN
            sigmoid_f := 43;
        ELSIF x =- 7850 THEN
            sigmoid_f := 43;
        ELSIF x =- 7849 THEN
            sigmoid_f := 43;
        ELSIF x =- 7848 THEN
            sigmoid_f := 43;
        ELSIF x =- 7847 THEN
            sigmoid_f := 43;
        ELSIF x =- 7846 THEN
            sigmoid_f := 43;
        ELSIF x =- 7845 THEN
            sigmoid_f := 43;
        ELSIF x =- 7844 THEN
            sigmoid_f := 43;
        ELSIF x =- 7843 THEN
            sigmoid_f := 43;
        ELSIF x =- 7842 THEN
            sigmoid_f := 43;
        ELSIF x =- 7841 THEN
            sigmoid_f := 43;
        ELSIF x =- 7840 THEN
            sigmoid_f := 43;
        ELSIF x =- 7839 THEN
            sigmoid_f := 43;
        ELSIF x =- 7838 THEN
            sigmoid_f := 43;
        ELSIF x =- 7837 THEN
            sigmoid_f := 43;
        ELSIF x =- 7836 THEN
            sigmoid_f := 43;
        ELSIF x =- 7835 THEN
            sigmoid_f := 43;
        ELSIF x =- 7834 THEN
            sigmoid_f := 43;
        ELSIF x =- 7833 THEN
            sigmoid_f := 43;
        ELSIF x =- 7832 THEN
            sigmoid_f := 43;
        ELSIF x =- 7831 THEN
            sigmoid_f := 43;
        ELSIF x =- 7830 THEN
            sigmoid_f := 43;
        ELSIF x =- 7829 THEN
            sigmoid_f := 43;
        ELSIF x =- 7828 THEN
            sigmoid_f := 43;
        ELSIF x =- 7827 THEN
            sigmoid_f := 43;
        ELSIF x =- 7826 THEN
            sigmoid_f := 43;
        ELSIF x =- 7825 THEN
            sigmoid_f := 43;
        ELSIF x =- 7824 THEN
            sigmoid_f := 44;
        ELSIF x =- 7823 THEN
            sigmoid_f := 44;
        ELSIF x =- 7822 THEN
            sigmoid_f := 44;
        ELSIF x =- 7821 THEN
            sigmoid_f := 44;
        ELSIF x =- 7820 THEN
            sigmoid_f := 44;
        ELSIF x =- 7819 THEN
            sigmoid_f := 44;
        ELSIF x =- 7818 THEN
            sigmoid_f := 44;
        ELSIF x =- 7817 THEN
            sigmoid_f := 44;
        ELSIF x =- 7816 THEN
            sigmoid_f := 44;
        ELSIF x =- 7815 THEN
            sigmoid_f := 44;
        ELSIF x =- 7814 THEN
            sigmoid_f := 44;
        ELSIF x =- 7813 THEN
            sigmoid_f := 44;
        ELSIF x =- 7812 THEN
            sigmoid_f := 44;
        ELSIF x =- 7811 THEN
            sigmoid_f := 44;
        ELSIF x =- 7810 THEN
            sigmoid_f := 44;
        ELSIF x =- 7809 THEN
            sigmoid_f := 44;
        ELSIF x =- 7808 THEN
            sigmoid_f := 44;
        ELSIF x =- 7807 THEN
            sigmoid_f := 44;
        ELSIF x =- 7806 THEN
            sigmoid_f := 44;
        ELSIF x =- 7805 THEN
            sigmoid_f := 44;
        ELSIF x =- 7804 THEN
            sigmoid_f := 44;
        ELSIF x =- 7803 THEN
            sigmoid_f := 44;
        ELSIF x =- 7802 THEN
            sigmoid_f := 44;
        ELSIF x =- 7801 THEN
            sigmoid_f := 44;
        ELSIF x =- 7800 THEN
            sigmoid_f := 44;
        ELSIF x =- 7799 THEN
            sigmoid_f := 44;
        ELSIF x =- 7798 THEN
            sigmoid_f := 44;
        ELSIF x =- 7797 THEN
            sigmoid_f := 44;
        ELSIF x =- 7796 THEN
            sigmoid_f := 44;
        ELSIF x =- 7795 THEN
            sigmoid_f := 44;
        ELSIF x =- 7794 THEN
            sigmoid_f := 44;
        ELSIF x =- 7793 THEN
            sigmoid_f := 44;
        ELSIF x =- 7792 THEN
            sigmoid_f := 44;
        ELSIF x =- 7791 THEN
            sigmoid_f := 44;
        ELSIF x =- 7790 THEN
            sigmoid_f := 44;
        ELSIF x =- 7789 THEN
            sigmoid_f := 44;
        ELSIF x =- 7788 THEN
            sigmoid_f := 44;
        ELSIF x =- 7787 THEN
            sigmoid_f := 44;
        ELSIF x =- 7786 THEN
            sigmoid_f := 44;
        ELSIF x =- 7785 THEN
            sigmoid_f := 44;
        ELSIF x =- 7784 THEN
            sigmoid_f := 44;
        ELSIF x =- 7783 THEN
            sigmoid_f := 44;
        ELSIF x =- 7782 THEN
            sigmoid_f := 44;
        ELSIF x =- 7781 THEN
            sigmoid_f := 44;
        ELSIF x =- 7780 THEN
            sigmoid_f := 44;
        ELSIF x =- 7779 THEN
            sigmoid_f := 44;
        ELSIF x =- 7778 THEN
            sigmoid_f := 44;
        ELSIF x =- 7777 THEN
            sigmoid_f := 44;
        ELSIF x =- 7776 THEN
            sigmoid_f := 44;
        ELSIF x =- 7775 THEN
            sigmoid_f := 44;
        ELSIF x =- 7774 THEN
            sigmoid_f := 44;
        ELSIF x =- 7773 THEN
            sigmoid_f := 44;
        ELSIF x =- 7772 THEN
            sigmoid_f := 44;
        ELSIF x =- 7771 THEN
            sigmoid_f := 45;
        ELSIF x =- 7770 THEN
            sigmoid_f := 45;
        ELSIF x =- 7769 THEN
            sigmoid_f := 45;
        ELSIF x =- 7768 THEN
            sigmoid_f := 45;
        ELSIF x =- 7767 THEN
            sigmoid_f := 45;
        ELSIF x =- 7766 THEN
            sigmoid_f := 45;
        ELSIF x =- 7765 THEN
            sigmoid_f := 45;
        ELSIF x =- 7764 THEN
            sigmoid_f := 45;
        ELSIF x =- 7763 THEN
            sigmoid_f := 45;
        ELSIF x =- 7762 THEN
            sigmoid_f := 45;
        ELSIF x =- 7761 THEN
            sigmoid_f := 45;
        ELSIF x =- 7760 THEN
            sigmoid_f := 45;
        ELSIF x =- 7759 THEN
            sigmoid_f := 45;
        ELSIF x =- 7758 THEN
            sigmoid_f := 45;
        ELSIF x =- 7757 THEN
            sigmoid_f := 45;
        ELSIF x =- 7756 THEN
            sigmoid_f := 45;
        ELSIF x =- 7755 THEN
            sigmoid_f := 45;
        ELSIF x =- 7754 THEN
            sigmoid_f := 45;
        ELSIF x =- 7753 THEN
            sigmoid_f := 45;
        ELSIF x =- 7752 THEN
            sigmoid_f := 45;
        ELSIF x =- 7751 THEN
            sigmoid_f := 45;
        ELSIF x =- 7750 THEN
            sigmoid_f := 45;
        ELSIF x =- 7749 THEN
            sigmoid_f := 45;
        ELSIF x =- 7748 THEN
            sigmoid_f := 45;
        ELSIF x =- 7747 THEN
            sigmoid_f := 45;
        ELSIF x =- 7746 THEN
            sigmoid_f := 45;
        ELSIF x =- 7745 THEN
            sigmoid_f := 45;
        ELSIF x =- 7744 THEN
            sigmoid_f := 45;
        ELSIF x =- 7743 THEN
            sigmoid_f := 45;
        ELSIF x =- 7742 THEN
            sigmoid_f := 45;
        ELSIF x =- 7741 THEN
            sigmoid_f := 45;
        ELSIF x =- 7740 THEN
            sigmoid_f := 45;
        ELSIF x =- 7739 THEN
            sigmoid_f := 45;
        ELSIF x =- 7738 THEN
            sigmoid_f := 45;
        ELSIF x =- 7737 THEN
            sigmoid_f := 45;
        ELSIF x =- 7736 THEN
            sigmoid_f := 45;
        ELSIF x =- 7735 THEN
            sigmoid_f := 45;
        ELSIF x =- 7734 THEN
            sigmoid_f := 45;
        ELSIF x =- 7733 THEN
            sigmoid_f := 45;
        ELSIF x =- 7732 THEN
            sigmoid_f := 45;
        ELSIF x =- 7731 THEN
            sigmoid_f := 45;
        ELSIF x =- 7730 THEN
            sigmoid_f := 45;
        ELSIF x =- 7729 THEN
            sigmoid_f := 45;
        ELSIF x =- 7728 THEN
            sigmoid_f := 45;
        ELSIF x =- 7727 THEN
            sigmoid_f := 45;
        ELSIF x =- 7726 THEN
            sigmoid_f := 45;
        ELSIF x =- 7725 THEN
            sigmoid_f := 45;
        ELSIF x =- 7724 THEN
            sigmoid_f := 45;
        ELSIF x =- 7723 THEN
            sigmoid_f := 45;
        ELSIF x =- 7722 THEN
            sigmoid_f := 45;
        ELSIF x =- 7721 THEN
            sigmoid_f := 45;
        ELSIF x =- 7720 THEN
            sigmoid_f := 45;
        ELSIF x =- 7719 THEN
            sigmoid_f := 46;
        ELSIF x =- 7718 THEN
            sigmoid_f := 46;
        ELSIF x =- 7717 THEN
            sigmoid_f := 46;
        ELSIF x =- 7716 THEN
            sigmoid_f := 46;
        ELSIF x =- 7715 THEN
            sigmoid_f := 46;
        ELSIF x =- 7714 THEN
            sigmoid_f := 46;
        ELSIF x =- 7713 THEN
            sigmoid_f := 46;
        ELSIF x =- 7712 THEN
            sigmoid_f := 46;
        ELSIF x =- 7711 THEN
            sigmoid_f := 46;
        ELSIF x =- 7710 THEN
            sigmoid_f := 46;
        ELSIF x =- 7709 THEN
            sigmoid_f := 46;
        ELSIF x =- 7708 THEN
            sigmoid_f := 46;
        ELSIF x =- 7707 THEN
            sigmoid_f := 46;
        ELSIF x =- 7706 THEN
            sigmoid_f := 46;
        ELSIF x =- 7705 THEN
            sigmoid_f := 46;
        ELSIF x =- 7704 THEN
            sigmoid_f := 46;
        ELSIF x =- 7703 THEN
            sigmoid_f := 46;
        ELSIF x =- 7702 THEN
            sigmoid_f := 46;
        ELSIF x =- 7701 THEN
            sigmoid_f := 46;
        ELSIF x =- 7700 THEN
            sigmoid_f := 46;
        ELSIF x =- 7699 THEN
            sigmoid_f := 46;
        ELSIF x =- 7698 THEN
            sigmoid_f := 46;
        ELSIF x =- 7697 THEN
            sigmoid_f := 46;
        ELSIF x =- 7696 THEN
            sigmoid_f := 46;
        ELSIF x =- 7695 THEN
            sigmoid_f := 46;
        ELSIF x =- 7694 THEN
            sigmoid_f := 46;
        ELSIF x =- 7693 THEN
            sigmoid_f := 46;
        ELSIF x =- 7692 THEN
            sigmoid_f := 46;
        ELSIF x =- 7691 THEN
            sigmoid_f := 46;
        ELSIF x =- 7690 THEN
            sigmoid_f := 46;
        ELSIF x =- 7689 THEN
            sigmoid_f := 46;
        ELSIF x =- 7688 THEN
            sigmoid_f := 46;
        ELSIF x =- 7687 THEN
            sigmoid_f := 46;
        ELSIF x =- 7686 THEN
            sigmoid_f := 46;
        ELSIF x =- 7685 THEN
            sigmoid_f := 46;
        ELSIF x =- 7684 THEN
            sigmoid_f := 46;
        ELSIF x =- 7683 THEN
            sigmoid_f := 46;
        ELSIF x =- 7682 THEN
            sigmoid_f := 46;
        ELSIF x =- 7681 THEN
            sigmoid_f := 46;
        ELSIF x =- 7680 THEN
            sigmoid_f := 46;
        ELSIF x =- 7679 THEN
            sigmoid_f := 46;
        ELSIF x =- 7678 THEN
            sigmoid_f := 46;
        ELSIF x =- 7677 THEN
            sigmoid_f := 46;
        ELSIF x =- 7676 THEN
            sigmoid_f := 46;
        ELSIF x =- 7675 THEN
            sigmoid_f := 46;
        ELSIF x =- 7674 THEN
            sigmoid_f := 46;
        ELSIF x =- 7673 THEN
            sigmoid_f := 46;
        ELSIF x =- 7672 THEN
            sigmoid_f := 46;
        ELSIF x =- 7671 THEN
            sigmoid_f := 46;
        ELSIF x =- 7670 THEN
            sigmoid_f := 46;
        ELSIF x =- 7669 THEN
            sigmoid_f := 46;
        ELSIF x =- 7668 THEN
            sigmoid_f := 46;
        ELSIF x =- 7667 THEN
            sigmoid_f := 46;
        ELSIF x =- 7666 THEN
            sigmoid_f := 46;
        ELSIF x =- 7665 THEN
            sigmoid_f := 46;
        ELSIF x =- 7664 THEN
            sigmoid_f := 46;
        ELSIF x =- 7663 THEN
            sigmoid_f := 46;
        ELSIF x =- 7662 THEN
            sigmoid_f := 46;
        ELSIF x =- 7661 THEN
            sigmoid_f := 47;
        ELSIF x =- 7660 THEN
            sigmoid_f := 47;
        ELSIF x =- 7659 THEN
            sigmoid_f := 47;
        ELSIF x =- 7658 THEN
            sigmoid_f := 47;
        ELSIF x =- 7657 THEN
            sigmoid_f := 47;
        ELSIF x =- 7656 THEN
            sigmoid_f := 47;
        ELSIF x =- 7655 THEN
            sigmoid_f := 47;
        ELSIF x =- 7654 THEN
            sigmoid_f := 47;
        ELSIF x =- 7653 THEN
            sigmoid_f := 47;
        ELSIF x =- 7652 THEN
            sigmoid_f := 47;
        ELSIF x =- 7651 THEN
            sigmoid_f := 47;
        ELSIF x =- 7650 THEN
            sigmoid_f := 47;
        ELSIF x =- 7649 THEN
            sigmoid_f := 47;
        ELSIF x =- 7648 THEN
            sigmoid_f := 47;
        ELSIF x =- 7647 THEN
            sigmoid_f := 47;
        ELSIF x =- 7646 THEN
            sigmoid_f := 47;
        ELSIF x =- 7645 THEN
            sigmoid_f := 47;
        ELSIF x =- 7644 THEN
            sigmoid_f := 47;
        ELSIF x =- 7643 THEN
            sigmoid_f := 47;
        ELSIF x =- 7642 THEN
            sigmoid_f := 47;
        ELSIF x =- 7641 THEN
            sigmoid_f := 47;
        ELSIF x =- 7640 THEN
            sigmoid_f := 47;
        ELSIF x =- 7639 THEN
            sigmoid_f := 47;
        ELSIF x =- 7638 THEN
            sigmoid_f := 47;
        ELSIF x =- 7637 THEN
            sigmoid_f := 47;
        ELSIF x =- 7636 THEN
            sigmoid_f := 47;
        ELSIF x =- 7635 THEN
            sigmoid_f := 47;
        ELSIF x =- 7634 THEN
            sigmoid_f := 47;
        ELSIF x =- 7633 THEN
            sigmoid_f := 47;
        ELSIF x =- 7632 THEN
            sigmoid_f := 47;
        ELSIF x =- 7631 THEN
            sigmoid_f := 47;
        ELSIF x =- 7630 THEN
            sigmoid_f := 47;
        ELSIF x =- 7629 THEN
            sigmoid_f := 47;
        ELSIF x =- 7628 THEN
            sigmoid_f := 47;
        ELSIF x =- 7627 THEN
            sigmoid_f := 47;
        ELSIF x =- 7626 THEN
            sigmoid_f := 47;
        ELSIF x =- 7625 THEN
            sigmoid_f := 47;
        ELSIF x =- 7624 THEN
            sigmoid_f := 47;
        ELSIF x =- 7623 THEN
            sigmoid_f := 48;
        ELSIF x =- 7622 THEN
            sigmoid_f := 48;
        ELSIF x =- 7621 THEN
            sigmoid_f := 48;
        ELSIF x =- 7620 THEN
            sigmoid_f := 48;
        ELSIF x =- 7619 THEN
            sigmoid_f := 48;
        ELSIF x =- 7618 THEN
            sigmoid_f := 48;
        ELSIF x =- 7617 THEN
            sigmoid_f := 48;
        ELSIF x =- 7616 THEN
            sigmoid_f := 48;
        ELSIF x =- 7615 THEN
            sigmoid_f := 48;
        ELSIF x =- 7614 THEN
            sigmoid_f := 48;
        ELSIF x =- 7613 THEN
            sigmoid_f := 48;
        ELSIF x =- 7612 THEN
            sigmoid_f := 48;
        ELSIF x =- 7611 THEN
            sigmoid_f := 48;
        ELSIF x =- 7610 THEN
            sigmoid_f := 48;
        ELSIF x =- 7609 THEN
            sigmoid_f := 48;
        ELSIF x =- 7608 THEN
            sigmoid_f := 48;
        ELSIF x =- 7607 THEN
            sigmoid_f := 48;
        ELSIF x =- 7606 THEN
            sigmoid_f := 48;
        ELSIF x =- 7605 THEN
            sigmoid_f := 48;
        ELSIF x =- 7604 THEN
            sigmoid_f := 48;
        ELSIF x =- 7603 THEN
            sigmoid_f := 48;
        ELSIF x =- 7602 THEN
            sigmoid_f := 48;
        ELSIF x =- 7601 THEN
            sigmoid_f := 48;
        ELSIF x =- 7600 THEN
            sigmoid_f := 48;
        ELSIF x =- 7599 THEN
            sigmoid_f := 48;
        ELSIF x =- 7598 THEN
            sigmoid_f := 48;
        ELSIF x =- 7597 THEN
            sigmoid_f := 48;
        ELSIF x =- 7596 THEN
            sigmoid_f := 48;
        ELSIF x =- 7595 THEN
            sigmoid_f := 48;
        ELSIF x =- 7594 THEN
            sigmoid_f := 48;
        ELSIF x =- 7593 THEN
            sigmoid_f := 48;
        ELSIF x =- 7592 THEN
            sigmoid_f := 48;
        ELSIF x =- 7591 THEN
            sigmoid_f := 48;
        ELSIF x =- 7590 THEN
            sigmoid_f := 48;
        ELSIF x =- 7589 THEN
            sigmoid_f := 48;
        ELSIF x =- 7588 THEN
            sigmoid_f := 48;
        ELSIF x =- 7587 THEN
            sigmoid_f := 48;
        ELSIF x =- 7586 THEN
            sigmoid_f := 48;
        ELSIF x =- 7585 THEN
            sigmoid_f := 49;
        ELSIF x =- 7584 THEN
            sigmoid_f := 49;
        ELSIF x =- 7583 THEN
            sigmoid_f := 49;
        ELSIF x =- 7582 THEN
            sigmoid_f := 49;
        ELSIF x =- 7581 THEN
            sigmoid_f := 49;
        ELSIF x =- 7580 THEN
            sigmoid_f := 49;
        ELSIF x =- 7579 THEN
            sigmoid_f := 49;
        ELSIF x =- 7578 THEN
            sigmoid_f := 49;
        ELSIF x =- 7577 THEN
            sigmoid_f := 49;
        ELSIF x =- 7576 THEN
            sigmoid_f := 49;
        ELSIF x =- 7575 THEN
            sigmoid_f := 49;
        ELSIF x =- 7574 THEN
            sigmoid_f := 49;
        ELSIF x =- 7573 THEN
            sigmoid_f := 49;
        ELSIF x =- 7572 THEN
            sigmoid_f := 49;
        ELSIF x =- 7571 THEN
            sigmoid_f := 49;
        ELSIF x =- 7570 THEN
            sigmoid_f := 49;
        ELSIF x =- 7569 THEN
            sigmoid_f := 49;
        ELSIF x =- 7568 THEN
            sigmoid_f := 49;
        ELSIF x =- 7567 THEN
            sigmoid_f := 49;
        ELSIF x =- 7566 THEN
            sigmoid_f := 49;
        ELSIF x =- 7565 THEN
            sigmoid_f := 49;
        ELSIF x =- 7564 THEN
            sigmoid_f := 49;
        ELSIF x =- 7563 THEN
            sigmoid_f := 49;
        ELSIF x =- 7562 THEN
            sigmoid_f := 49;
        ELSIF x =- 7561 THEN
            sigmoid_f := 49;
        ELSIF x =- 7560 THEN
            sigmoid_f := 49;
        ELSIF x =- 7559 THEN
            sigmoid_f := 49;
        ELSIF x =- 7558 THEN
            sigmoid_f := 49;
        ELSIF x =- 7557 THEN
            sigmoid_f := 49;
        ELSIF x =- 7556 THEN
            sigmoid_f := 49;
        ELSIF x =- 7555 THEN
            sigmoid_f := 49;
        ELSIF x =- 7554 THEN
            sigmoid_f := 49;
        ELSIF x =- 7553 THEN
            sigmoid_f := 49;
        ELSIF x =- 7552 THEN
            sigmoid_f := 49;
        ELSIF x =- 7551 THEN
            sigmoid_f := 49;
        ELSIF x =- 7550 THEN
            sigmoid_f := 49;
        ELSIF x =- 7549 THEN
            sigmoid_f := 49;
        ELSIF x =- 7548 THEN
            sigmoid_f := 49;
        ELSIF x =- 7547 THEN
            sigmoid_f := 50;
        ELSIF x =- 7546 THEN
            sigmoid_f := 50;
        ELSIF x =- 7545 THEN
            sigmoid_f := 50;
        ELSIF x =- 7544 THEN
            sigmoid_f := 50;
        ELSIF x =- 7543 THEN
            sigmoid_f := 50;
        ELSIF x =- 7542 THEN
            sigmoid_f := 50;
        ELSIF x =- 7541 THEN
            sigmoid_f := 50;
        ELSIF x =- 7540 THEN
            sigmoid_f := 50;
        ELSIF x =- 7539 THEN
            sigmoid_f := 50;
        ELSIF x =- 7538 THEN
            sigmoid_f := 50;
        ELSIF x =- 7537 THEN
            sigmoid_f := 50;
        ELSIF x =- 7536 THEN
            sigmoid_f := 50;
        ELSIF x =- 7535 THEN
            sigmoid_f := 50;
        ELSIF x =- 7534 THEN
            sigmoid_f := 50;
        ELSIF x =- 7533 THEN
            sigmoid_f := 50;
        ELSIF x =- 7532 THEN
            sigmoid_f := 50;
        ELSIF x =- 7531 THEN
            sigmoid_f := 50;
        ELSIF x =- 7530 THEN
            sigmoid_f := 50;
        ELSIF x =- 7529 THEN
            sigmoid_f := 50;
        ELSIF x =- 7528 THEN
            sigmoid_f := 50;
        ELSIF x =- 7527 THEN
            sigmoid_f := 50;
        ELSIF x =- 7526 THEN
            sigmoid_f := 50;
        ELSIF x =- 7525 THEN
            sigmoid_f := 50;
        ELSIF x =- 7524 THEN
            sigmoid_f := 50;
        ELSIF x =- 7523 THEN
            sigmoid_f := 50;
        ELSIF x =- 7522 THEN
            sigmoid_f := 50;
        ELSIF x =- 7521 THEN
            sigmoid_f := 50;
        ELSIF x =- 7520 THEN
            sigmoid_f := 50;
        ELSIF x =- 7519 THEN
            sigmoid_f := 50;
        ELSIF x =- 7518 THEN
            sigmoid_f := 50;
        ELSIF x =- 7517 THEN
            sigmoid_f := 50;
        ELSIF x =- 7516 THEN
            sigmoid_f := 50;
        ELSIF x =- 7515 THEN
            sigmoid_f := 50;
        ELSIF x =- 7514 THEN
            sigmoid_f := 50;
        ELSIF x =- 7513 THEN
            sigmoid_f := 50;
        ELSIF x =- 7512 THEN
            sigmoid_f := 50;
        ELSIF x =- 7511 THEN
            sigmoid_f := 50;
        ELSIF x =- 7510 THEN
            sigmoid_f := 50;
        ELSIF x =- 7509 THEN
            sigmoid_f := 51;
        ELSIF x =- 7508 THEN
            sigmoid_f := 51;
        ELSIF x =- 7507 THEN
            sigmoid_f := 51;
        ELSIF x =- 7506 THEN
            sigmoid_f := 51;
        ELSIF x =- 7505 THEN
            sigmoid_f := 51;
        ELSIF x =- 7504 THEN
            sigmoid_f := 51;
        ELSIF x =- 7503 THEN
            sigmoid_f := 51;
        ELSIF x =- 7502 THEN
            sigmoid_f := 51;
        ELSIF x =- 7501 THEN
            sigmoid_f := 51;
        ELSIF x =- 7500 THEN
            sigmoid_f := 51;
        ELSIF x =- 7499 THEN
            sigmoid_f := 51;
        ELSIF x =- 7498 THEN
            sigmoid_f := 51;
        ELSIF x =- 7497 THEN
            sigmoid_f := 51;
        ELSIF x =- 7496 THEN
            sigmoid_f := 51;
        ELSIF x =- 7495 THEN
            sigmoid_f := 51;
        ELSIF x =- 7494 THEN
            sigmoid_f := 51;
        ELSIF x =- 7493 THEN
            sigmoid_f := 51;
        ELSIF x =- 7492 THEN
            sigmoid_f := 51;
        ELSIF x =- 7491 THEN
            sigmoid_f := 51;
        ELSIF x =- 7490 THEN
            sigmoid_f := 51;
        ELSIF x =- 7489 THEN
            sigmoid_f := 51;
        ELSIF x =- 7488 THEN
            sigmoid_f := 51;
        ELSIF x =- 7487 THEN
            sigmoid_f := 51;
        ELSIF x =- 7486 THEN
            sigmoid_f := 51;
        ELSIF x =- 7485 THEN
            sigmoid_f := 51;
        ELSIF x =- 7484 THEN
            sigmoid_f := 51;
        ELSIF x =- 7483 THEN
            sigmoid_f := 51;
        ELSIF x =- 7482 THEN
            sigmoid_f := 51;
        ELSIF x =- 7481 THEN
            sigmoid_f := 51;
        ELSIF x =- 7480 THEN
            sigmoid_f := 51;
        ELSIF x =- 7479 THEN
            sigmoid_f := 51;
        ELSIF x =- 7478 THEN
            sigmoid_f := 51;
        ELSIF x =- 7477 THEN
            sigmoid_f := 51;
        ELSIF x =- 7476 THEN
            sigmoid_f := 51;
        ELSIF x =- 7475 THEN
            sigmoid_f := 51;
        ELSIF x =- 7474 THEN
            sigmoid_f := 51;
        ELSIF x =- 7473 THEN
            sigmoid_f := 51;
        ELSIF x =- 7472 THEN
            sigmoid_f := 51;
        ELSIF x =- 7471 THEN
            sigmoid_f := 52;
        ELSIF x =- 7470 THEN
            sigmoid_f := 52;
        ELSIF x =- 7469 THEN
            sigmoid_f := 52;
        ELSIF x =- 7468 THEN
            sigmoid_f := 52;
        ELSIF x =- 7467 THEN
            sigmoid_f := 52;
        ELSIF x =- 7466 THEN
            sigmoid_f := 52;
        ELSIF x =- 7465 THEN
            sigmoid_f := 52;
        ELSIF x =- 7464 THEN
            sigmoid_f := 52;
        ELSIF x =- 7463 THEN
            sigmoid_f := 52;
        ELSIF x =- 7462 THEN
            sigmoid_f := 52;
        ELSIF x =- 7461 THEN
            sigmoid_f := 52;
        ELSIF x =- 7460 THEN
            sigmoid_f := 52;
        ELSIF x =- 7459 THEN
            sigmoid_f := 52;
        ELSIF x =- 7458 THEN
            sigmoid_f := 52;
        ELSIF x =- 7457 THEN
            sigmoid_f := 52;
        ELSIF x =- 7456 THEN
            sigmoid_f := 52;
        ELSIF x =- 7455 THEN
            sigmoid_f := 52;
        ELSIF x =- 7454 THEN
            sigmoid_f := 52;
        ELSIF x =- 7453 THEN
            sigmoid_f := 52;
        ELSIF x =- 7452 THEN
            sigmoid_f := 52;
        ELSIF x =- 7451 THEN
            sigmoid_f := 52;
        ELSIF x =- 7450 THEN
            sigmoid_f := 52;
        ELSIF x =- 7449 THEN
            sigmoid_f := 52;
        ELSIF x =- 7448 THEN
            sigmoid_f := 52;
        ELSIF x =- 7447 THEN
            sigmoid_f := 52;
        ELSIF x =- 7446 THEN
            sigmoid_f := 52;
        ELSIF x =- 7445 THEN
            sigmoid_f := 52;
        ELSIF x =- 7444 THEN
            sigmoid_f := 52;
        ELSIF x =- 7443 THEN
            sigmoid_f := 52;
        ELSIF x =- 7442 THEN
            sigmoid_f := 52;
        ELSIF x =- 7441 THEN
            sigmoid_f := 52;
        ELSIF x =- 7440 THEN
            sigmoid_f := 52;
        ELSIF x =- 7439 THEN
            sigmoid_f := 52;
        ELSIF x =- 7438 THEN
            sigmoid_f := 52;
        ELSIF x =- 7437 THEN
            sigmoid_f := 52;
        ELSIF x =- 7436 THEN
            sigmoid_f := 52;
        ELSIF x =- 7435 THEN
            sigmoid_f := 52;
        ELSIF x =- 7434 THEN
            sigmoid_f := 52;
        ELSIF x =- 7433 THEN
            sigmoid_f := 53;
        ELSIF x =- 7432 THEN
            sigmoid_f := 53;
        ELSIF x =- 7431 THEN
            sigmoid_f := 53;
        ELSIF x =- 7430 THEN
            sigmoid_f := 53;
        ELSIF x =- 7429 THEN
            sigmoid_f := 53;
        ELSIF x =- 7428 THEN
            sigmoid_f := 53;
        ELSIF x =- 7427 THEN
            sigmoid_f := 53;
        ELSIF x =- 7426 THEN
            sigmoid_f := 53;
        ELSIF x =- 7425 THEN
            sigmoid_f := 53;
        ELSIF x =- 7424 THEN
            sigmoid_f := 53;
        ELSIF x =- 7423 THEN
            sigmoid_f := 53;
        ELSIF x =- 7422 THEN
            sigmoid_f := 53;
        ELSIF x =- 7421 THEN
            sigmoid_f := 53;
        ELSIF x =- 7420 THEN
            sigmoid_f := 53;
        ELSIF x =- 7419 THEN
            sigmoid_f := 53;
        ELSIF x =- 7418 THEN
            sigmoid_f := 53;
        ELSIF x =- 7417 THEN
            sigmoid_f := 53;
        ELSIF x =- 7416 THEN
            sigmoid_f := 53;
        ELSIF x =- 7415 THEN
            sigmoid_f := 53;
        ELSIF x =- 7414 THEN
            sigmoid_f := 53;
        ELSIF x =- 7413 THEN
            sigmoid_f := 53;
        ELSIF x =- 7412 THEN
            sigmoid_f := 53;
        ELSIF x =- 7411 THEN
            sigmoid_f := 53;
        ELSIF x =- 7410 THEN
            sigmoid_f := 53;
        ELSIF x =- 7409 THEN
            sigmoid_f := 53;
        ELSIF x =- 7408 THEN
            sigmoid_f := 53;
        ELSIF x =- 7407 THEN
            sigmoid_f := 53;
        ELSIF x =- 7406 THEN
            sigmoid_f := 53;
        ELSIF x =- 7405 THEN
            sigmoid_f := 53;
        ELSIF x =- 7404 THEN
            sigmoid_f := 53;
        ELSIF x =- 7403 THEN
            sigmoid_f := 53;
        ELSIF x =- 7402 THEN
            sigmoid_f := 53;
        ELSIF x =- 7401 THEN
            sigmoid_f := 53;
        ELSIF x =- 7400 THEN
            sigmoid_f := 53;
        ELSIF x =- 7399 THEN
            sigmoid_f := 53;
        ELSIF x =- 7398 THEN
            sigmoid_f := 53;
        ELSIF x =- 7397 THEN
            sigmoid_f := 53;
        ELSIF x =- 7396 THEN
            sigmoid_f := 53;
        ELSIF x =- 7395 THEN
            sigmoid_f := 54;
        ELSIF x =- 7394 THEN
            sigmoid_f := 54;
        ELSIF x =- 7393 THEN
            sigmoid_f := 54;
        ELSIF x =- 7392 THEN
            sigmoid_f := 54;
        ELSIF x =- 7391 THEN
            sigmoid_f := 54;
        ELSIF x =- 7390 THEN
            sigmoid_f := 54;
        ELSIF x =- 7389 THEN
            sigmoid_f := 54;
        ELSIF x =- 7388 THEN
            sigmoid_f := 54;
        ELSIF x =- 7387 THEN
            sigmoid_f := 54;
        ELSIF x =- 7386 THEN
            sigmoid_f := 54;
        ELSIF x =- 7385 THEN
            sigmoid_f := 54;
        ELSIF x =- 7384 THEN
            sigmoid_f := 54;
        ELSIF x =- 7383 THEN
            sigmoid_f := 54;
        ELSIF x =- 7382 THEN
            sigmoid_f := 54;
        ELSIF x =- 7381 THEN
            sigmoid_f := 54;
        ELSIF x =- 7380 THEN
            sigmoid_f := 54;
        ELSIF x =- 7379 THEN
            sigmoid_f := 54;
        ELSIF x =- 7378 THEN
            sigmoid_f := 54;
        ELSIF x =- 7377 THEN
            sigmoid_f := 54;
        ELSIF x =- 7376 THEN
            sigmoid_f := 54;
        ELSIF x =- 7375 THEN
            sigmoid_f := 54;
        ELSIF x =- 7374 THEN
            sigmoid_f := 54;
        ELSIF x =- 7373 THEN
            sigmoid_f := 54;
        ELSIF x =- 7372 THEN
            sigmoid_f := 54;
        ELSIF x =- 7371 THEN
            sigmoid_f := 54;
        ELSIF x =- 7370 THEN
            sigmoid_f := 54;
        ELSIF x =- 7369 THEN
            sigmoid_f := 54;
        ELSIF x =- 7368 THEN
            sigmoid_f := 54;
        ELSIF x =- 7367 THEN
            sigmoid_f := 54;
        ELSIF x =- 7366 THEN
            sigmoid_f := 54;
        ELSIF x =- 7365 THEN
            sigmoid_f := 54;
        ELSIF x =- 7364 THEN
            sigmoid_f := 54;
        ELSIF x =- 7363 THEN
            sigmoid_f := 54;
        ELSIF x =- 7362 THEN
            sigmoid_f := 54;
        ELSIF x =- 7361 THEN
            sigmoid_f := 54;
        ELSIF x =- 7360 THEN
            sigmoid_f := 54;
        ELSIF x =- 7359 THEN
            sigmoid_f := 54;
        ELSIF x =- 7358 THEN
            sigmoid_f := 54;
        ELSIF x =- 7357 THEN
            sigmoid_f := 55;
        ELSIF x =- 7356 THEN
            sigmoid_f := 55;
        ELSIF x =- 7355 THEN
            sigmoid_f := 55;
        ELSIF x =- 7354 THEN
            sigmoid_f := 55;
        ELSIF x =- 7353 THEN
            sigmoid_f := 55;
        ELSIF x =- 7352 THEN
            sigmoid_f := 55;
        ELSIF x =- 7351 THEN
            sigmoid_f := 55;
        ELSIF x =- 7350 THEN
            sigmoid_f := 55;
        ELSIF x =- 7349 THEN
            sigmoid_f := 55;
        ELSIF x =- 7348 THEN
            sigmoid_f := 55;
        ELSIF x =- 7347 THEN
            sigmoid_f := 55;
        ELSIF x =- 7346 THEN
            sigmoid_f := 55;
        ELSIF x =- 7345 THEN
            sigmoid_f := 55;
        ELSIF x =- 7344 THEN
            sigmoid_f := 55;
        ELSIF x =- 7343 THEN
            sigmoid_f := 55;
        ELSIF x =- 7342 THEN
            sigmoid_f := 55;
        ELSIF x =- 7341 THEN
            sigmoid_f := 55;
        ELSIF x =- 7340 THEN
            sigmoid_f := 55;
        ELSIF x =- 7339 THEN
            sigmoid_f := 55;
        ELSIF x =- 7338 THEN
            sigmoid_f := 55;
        ELSIF x =- 7337 THEN
            sigmoid_f := 55;
        ELSIF x =- 7336 THEN
            sigmoid_f := 55;
        ELSIF x =- 7335 THEN
            sigmoid_f := 55;
        ELSIF x =- 7334 THEN
            sigmoid_f := 55;
        ELSIF x =- 7333 THEN
            sigmoid_f := 55;
        ELSIF x =- 7332 THEN
            sigmoid_f := 55;
        ELSIF x =- 7331 THEN
            sigmoid_f := 55;
        ELSIF x =- 7330 THEN
            sigmoid_f := 55;
        ELSIF x =- 7329 THEN
            sigmoid_f := 55;
        ELSIF x =- 7328 THEN
            sigmoid_f := 55;
        ELSIF x =- 7327 THEN
            sigmoid_f := 55;
        ELSIF x =- 7326 THEN
            sigmoid_f := 55;
        ELSIF x =- 7325 THEN
            sigmoid_f := 55;
        ELSIF x =- 7324 THEN
            sigmoid_f := 55;
        ELSIF x =- 7323 THEN
            sigmoid_f := 55;
        ELSIF x =- 7322 THEN
            sigmoid_f := 55;
        ELSIF x =- 7321 THEN
            sigmoid_f := 55;
        ELSIF x =- 7320 THEN
            sigmoid_f := 55;
        ELSIF x =- 7319 THEN
            sigmoid_f := 56;
        ELSIF x =- 7318 THEN
            sigmoid_f := 56;
        ELSIF x =- 7317 THEN
            sigmoid_f := 56;
        ELSIF x =- 7316 THEN
            sigmoid_f := 56;
        ELSIF x =- 7315 THEN
            sigmoid_f := 56;
        ELSIF x =- 7314 THEN
            sigmoid_f := 56;
        ELSIF x =- 7313 THEN
            sigmoid_f := 56;
        ELSIF x =- 7312 THEN
            sigmoid_f := 56;
        ELSIF x =- 7311 THEN
            sigmoid_f := 56;
        ELSIF x =- 7310 THEN
            sigmoid_f := 56;
        ELSIF x =- 7309 THEN
            sigmoid_f := 56;
        ELSIF x =- 7308 THEN
            sigmoid_f := 56;
        ELSIF x =- 7307 THEN
            sigmoid_f := 56;
        ELSIF x =- 7306 THEN
            sigmoid_f := 56;
        ELSIF x =- 7305 THEN
            sigmoid_f := 56;
        ELSIF x =- 7304 THEN
            sigmoid_f := 56;
        ELSIF x =- 7303 THEN
            sigmoid_f := 56;
        ELSIF x =- 7302 THEN
            sigmoid_f := 56;
        ELSIF x =- 7301 THEN
            sigmoid_f := 56;
        ELSIF x =- 7300 THEN
            sigmoid_f := 56;
        ELSIF x =- 7299 THEN
            sigmoid_f := 56;
        ELSIF x =- 7298 THEN
            sigmoid_f := 56;
        ELSIF x =- 7297 THEN
            sigmoid_f := 56;
        ELSIF x =- 7296 THEN
            sigmoid_f := 56;
        ELSIF x =- 7295 THEN
            sigmoid_f := 56;
        ELSIF x =- 7294 THEN
            sigmoid_f := 56;
        ELSIF x =- 7293 THEN
            sigmoid_f := 56;
        ELSIF x =- 7292 THEN
            sigmoid_f := 56;
        ELSIF x =- 7291 THEN
            sigmoid_f := 56;
        ELSIF x =- 7290 THEN
            sigmoid_f := 56;
        ELSIF x =- 7289 THEN
            sigmoid_f := 56;
        ELSIF x =- 7288 THEN
            sigmoid_f := 56;
        ELSIF x =- 7287 THEN
            sigmoid_f := 56;
        ELSIF x =- 7286 THEN
            sigmoid_f := 56;
        ELSIF x =- 7285 THEN
            sigmoid_f := 56;
        ELSIF x =- 7284 THEN
            sigmoid_f := 56;
        ELSIF x =- 7283 THEN
            sigmoid_f := 56;
        ELSIF x =- 7282 THEN
            sigmoid_f := 56;
        ELSIF x =- 7281 THEN
            sigmoid_f := 57;
        ELSIF x =- 7280 THEN
            sigmoid_f := 57;
        ELSIF x =- 7279 THEN
            sigmoid_f := 57;
        ELSIF x =- 7278 THEN
            sigmoid_f := 57;
        ELSIF x =- 7277 THEN
            sigmoid_f := 57;
        ELSIF x =- 7276 THEN
            sigmoid_f := 57;
        ELSIF x =- 7275 THEN
            sigmoid_f := 57;
        ELSIF x =- 7274 THEN
            sigmoid_f := 57;
        ELSIF x =- 7273 THEN
            sigmoid_f := 57;
        ELSIF x =- 7272 THEN
            sigmoid_f := 57;
        ELSIF x =- 7271 THEN
            sigmoid_f := 57;
        ELSIF x =- 7270 THEN
            sigmoid_f := 57;
        ELSIF x =- 7269 THEN
            sigmoid_f := 57;
        ELSIF x =- 7268 THEN
            sigmoid_f := 57;
        ELSIF x =- 7267 THEN
            sigmoid_f := 57;
        ELSIF x =- 7266 THEN
            sigmoid_f := 57;
        ELSIF x =- 7265 THEN
            sigmoid_f := 57;
        ELSIF x =- 7264 THEN
            sigmoid_f := 57;
        ELSIF x =- 7263 THEN
            sigmoid_f := 57;
        ELSIF x =- 7262 THEN
            sigmoid_f := 57;
        ELSIF x =- 7261 THEN
            sigmoid_f := 57;
        ELSIF x =- 7260 THEN
            sigmoid_f := 57;
        ELSIF x =- 7259 THEN
            sigmoid_f := 57;
        ELSIF x =- 7258 THEN
            sigmoid_f := 57;
        ELSIF x =- 7257 THEN
            sigmoid_f := 57;
        ELSIF x =- 7256 THEN
            sigmoid_f := 57;
        ELSIF x =- 7255 THEN
            sigmoid_f := 57;
        ELSIF x =- 7254 THEN
            sigmoid_f := 57;
        ELSIF x =- 7253 THEN
            sigmoid_f := 57;
        ELSIF x =- 7252 THEN
            sigmoid_f := 57;
        ELSIF x =- 7251 THEN
            sigmoid_f := 57;
        ELSIF x =- 7250 THEN
            sigmoid_f := 57;
        ELSIF x =- 7249 THEN
            sigmoid_f := 57;
        ELSIF x =- 7248 THEN
            sigmoid_f := 57;
        ELSIF x =- 7247 THEN
            sigmoid_f := 57;
        ELSIF x =- 7246 THEN
            sigmoid_f := 57;
        ELSIF x =- 7245 THEN
            sigmoid_f := 57;
        ELSIF x =- 7244 THEN
            sigmoid_f := 57;
        ELSIF x =- 7243 THEN
            sigmoid_f := 58;
        ELSIF x =- 7242 THEN
            sigmoid_f := 58;
        ELSIF x =- 7241 THEN
            sigmoid_f := 58;
        ELSIF x =- 7240 THEN
            sigmoid_f := 58;
        ELSIF x =- 7239 THEN
            sigmoid_f := 58;
        ELSIF x =- 7238 THEN
            sigmoid_f := 58;
        ELSIF x =- 7237 THEN
            sigmoid_f := 58;
        ELSIF x =- 7236 THEN
            sigmoid_f := 58;
        ELSIF x =- 7235 THEN
            sigmoid_f := 58;
        ELSIF x =- 7234 THEN
            sigmoid_f := 58;
        ELSIF x =- 7233 THEN
            sigmoid_f := 58;
        ELSIF x =- 7232 THEN
            sigmoid_f := 58;
        ELSIF x =- 7231 THEN
            sigmoid_f := 58;
        ELSIF x =- 7230 THEN
            sigmoid_f := 58;
        ELSIF x =- 7229 THEN
            sigmoid_f := 58;
        ELSIF x =- 7228 THEN
            sigmoid_f := 58;
        ELSIF x =- 7227 THEN
            sigmoid_f := 58;
        ELSIF x =- 7226 THEN
            sigmoid_f := 58;
        ELSIF x =- 7225 THEN
            sigmoid_f := 58;
        ELSIF x =- 7224 THEN
            sigmoid_f := 58;
        ELSIF x =- 7223 THEN
            sigmoid_f := 58;
        ELSIF x =- 7222 THEN
            sigmoid_f := 58;
        ELSIF x =- 7221 THEN
            sigmoid_f := 58;
        ELSIF x =- 7220 THEN
            sigmoid_f := 58;
        ELSIF x =- 7219 THEN
            sigmoid_f := 58;
        ELSIF x =- 7218 THEN
            sigmoid_f := 58;
        ELSIF x =- 7217 THEN
            sigmoid_f := 58;
        ELSIF x =- 7216 THEN
            sigmoid_f := 58;
        ELSIF x =- 7215 THEN
            sigmoid_f := 58;
        ELSIF x =- 7214 THEN
            sigmoid_f := 58;
        ELSIF x =- 7213 THEN
            sigmoid_f := 58;
        ELSIF x =- 7212 THEN
            sigmoid_f := 58;
        ELSIF x =- 7211 THEN
            sigmoid_f := 58;
        ELSIF x =- 7210 THEN
            sigmoid_f := 58;
        ELSIF x =- 7209 THEN
            sigmoid_f := 58;
        ELSIF x =- 7208 THEN
            sigmoid_f := 58;
        ELSIF x =- 7207 THEN
            sigmoid_f := 58;
        ELSIF x =- 7206 THEN
            sigmoid_f := 58;
        ELSIF x =- 7205 THEN
            sigmoid_f := 59;
        ELSIF x =- 7204 THEN
            sigmoid_f := 59;
        ELSIF x =- 7203 THEN
            sigmoid_f := 59;
        ELSIF x =- 7202 THEN
            sigmoid_f := 59;
        ELSIF x =- 7201 THEN
            sigmoid_f := 59;
        ELSIF x =- 7200 THEN
            sigmoid_f := 59;
        ELSIF x =- 7199 THEN
            sigmoid_f := 59;
        ELSIF x =- 7198 THEN
            sigmoid_f := 59;
        ELSIF x =- 7197 THEN
            sigmoid_f := 59;
        ELSIF x =- 7196 THEN
            sigmoid_f := 59;
        ELSIF x =- 7195 THEN
            sigmoid_f := 59;
        ELSIF x =- 7194 THEN
            sigmoid_f := 59;
        ELSIF x =- 7193 THEN
            sigmoid_f := 59;
        ELSIF x =- 7192 THEN
            sigmoid_f := 59;
        ELSIF x =- 7191 THEN
            sigmoid_f := 59;
        ELSIF x =- 7190 THEN
            sigmoid_f := 59;
        ELSIF x =- 7189 THEN
            sigmoid_f := 59;
        ELSIF x =- 7188 THEN
            sigmoid_f := 59;
        ELSIF x =- 7187 THEN
            sigmoid_f := 59;
        ELSIF x =- 7186 THEN
            sigmoid_f := 59;
        ELSIF x =- 7185 THEN
            sigmoid_f := 59;
        ELSIF x =- 7184 THEN
            sigmoid_f := 59;
        ELSIF x =- 7183 THEN
            sigmoid_f := 59;
        ELSIF x =- 7182 THEN
            sigmoid_f := 59;
        ELSIF x =- 7181 THEN
            sigmoid_f := 59;
        ELSIF x =- 7180 THEN
            sigmoid_f := 59;
        ELSIF x =- 7179 THEN
            sigmoid_f := 59;
        ELSIF x =- 7178 THEN
            sigmoid_f := 59;
        ELSIF x =- 7177 THEN
            sigmoid_f := 59;
        ELSIF x =- 7176 THEN
            sigmoid_f := 59;
        ELSIF x =- 7175 THEN
            sigmoid_f := 59;
        ELSIF x =- 7174 THEN
            sigmoid_f := 59;
        ELSIF x =- 7173 THEN
            sigmoid_f := 59;
        ELSIF x =- 7172 THEN
            sigmoid_f := 59;
        ELSIF x =- 7171 THEN
            sigmoid_f := 59;
        ELSIF x =- 7170 THEN
            sigmoid_f := 59;
        ELSIF x =- 7169 THEN
            sigmoid_f := 59;
        ELSIF x =- 7168 THEN
            sigmoid_f := 60;
        ELSIF x =- 7167 THEN
            sigmoid_f := 60;
        ELSIF x =- 7166 THEN
            sigmoid_f := 60;
        ELSIF x =- 7165 THEN
            sigmoid_f := 60;
        ELSIF x =- 7164 THEN
            sigmoid_f := 60;
        ELSIF x =- 7163 THEN
            sigmoid_f := 60;
        ELSIF x =- 7162 THEN
            sigmoid_f := 60;
        ELSIF x =- 7161 THEN
            sigmoid_f := 60;
        ELSIF x =- 7160 THEN
            sigmoid_f := 60;
        ELSIF x =- 7159 THEN
            sigmoid_f := 60;
        ELSIF x =- 7158 THEN
            sigmoid_f := 60;
        ELSIF x =- 7157 THEN
            sigmoid_f := 60;
        ELSIF x =- 7156 THEN
            sigmoid_f := 60;
        ELSIF x =- 7155 THEN
            sigmoid_f := 60;
        ELSIF x =- 7154 THEN
            sigmoid_f := 60;
        ELSIF x =- 7153 THEN
            sigmoid_f := 60;
        ELSIF x =- 7152 THEN
            sigmoid_f := 60;
        ELSIF x =- 7151 THEN
            sigmoid_f := 60;
        ELSIF x =- 7150 THEN
            sigmoid_f := 60;
        ELSIF x =- 7149 THEN
            sigmoid_f := 60;
        ELSIF x =- 7148 THEN
            sigmoid_f := 60;
        ELSIF x =- 7147 THEN
            sigmoid_f := 60;
        ELSIF x =- 7146 THEN
            sigmoid_f := 60;
        ELSIF x =- 7145 THEN
            sigmoid_f := 60;
        ELSIF x =- 7144 THEN
            sigmoid_f := 60;
        ELSIF x =- 7143 THEN
            sigmoid_f := 60;
        ELSIF x =- 7142 THEN
            sigmoid_f := 60;
        ELSIF x =- 7141 THEN
            sigmoid_f := 60;
        ELSIF x =- 7140 THEN
            sigmoid_f := 60;
        ELSIF x =- 7139 THEN
            sigmoid_f := 60;
        ELSIF x =- 7138 THEN
            sigmoid_f := 60;
        ELSIF x =- 7137 THEN
            sigmoid_f := 60;
        ELSIF x =- 7136 THEN
            sigmoid_f := 61;
        ELSIF x =- 7135 THEN
            sigmoid_f := 61;
        ELSIF x =- 7134 THEN
            sigmoid_f := 61;
        ELSIF x =- 7133 THEN
            sigmoid_f := 61;
        ELSIF x =- 7132 THEN
            sigmoid_f := 61;
        ELSIF x =- 7131 THEN
            sigmoid_f := 61;
        ELSIF x =- 7130 THEN
            sigmoid_f := 61;
        ELSIF x =- 7129 THEN
            sigmoid_f := 61;
        ELSIF x =- 7128 THEN
            sigmoid_f := 61;
        ELSIF x =- 7127 THEN
            sigmoid_f := 61;
        ELSIF x =- 7126 THEN
            sigmoid_f := 61;
        ELSIF x =- 7125 THEN
            sigmoid_f := 61;
        ELSIF x =- 7124 THEN
            sigmoid_f := 61;
        ELSIF x =- 7123 THEN
            sigmoid_f := 61;
        ELSIF x =- 7122 THEN
            sigmoid_f := 61;
        ELSIF x =- 7121 THEN
            sigmoid_f := 61;
        ELSIF x =- 7120 THEN
            sigmoid_f := 61;
        ELSIF x =- 7119 THEN
            sigmoid_f := 61;
        ELSIF x =- 7118 THEN
            sigmoid_f := 61;
        ELSIF x =- 7117 THEN
            sigmoid_f := 61;
        ELSIF x =- 7116 THEN
            sigmoid_f := 61;
        ELSIF x =- 7115 THEN
            sigmoid_f := 61;
        ELSIF x =- 7114 THEN
            sigmoid_f := 61;
        ELSIF x =- 7113 THEN
            sigmoid_f := 61;
        ELSIF x =- 7112 THEN
            sigmoid_f := 61;
        ELSIF x =- 7111 THEN
            sigmoid_f := 61;
        ELSIF x =- 7110 THEN
            sigmoid_f := 61;
        ELSIF x =- 7109 THEN
            sigmoid_f := 61;
        ELSIF x =- 7108 THEN
            sigmoid_f := 61;
        ELSIF x =- 7107 THEN
            sigmoid_f := 61;
        ELSIF x =- 7106 THEN
            sigmoid_f := 61;
        ELSIF x =- 7105 THEN
            sigmoid_f := 61;
        ELSIF x =- 7104 THEN
            sigmoid_f := 62;
        ELSIF x =- 7103 THEN
            sigmoid_f := 62;
        ELSIF x =- 7102 THEN
            sigmoid_f := 62;
        ELSIF x =- 7101 THEN
            sigmoid_f := 62;
        ELSIF x =- 7100 THEN
            sigmoid_f := 62;
        ELSIF x =- 7099 THEN
            sigmoid_f := 62;
        ELSIF x =- 7098 THEN
            sigmoid_f := 62;
        ELSIF x =- 7097 THEN
            sigmoid_f := 62;
        ELSIF x =- 7096 THEN
            sigmoid_f := 62;
        ELSIF x =- 7095 THEN
            sigmoid_f := 62;
        ELSIF x =- 7094 THEN
            sigmoid_f := 62;
        ELSIF x =- 7093 THEN
            sigmoid_f := 62;
        ELSIF x =- 7092 THEN
            sigmoid_f := 62;
        ELSIF x =- 7091 THEN
            sigmoid_f := 62;
        ELSIF x =- 7090 THEN
            sigmoid_f := 62;
        ELSIF x =- 7089 THEN
            sigmoid_f := 62;
        ELSIF x =- 7088 THEN
            sigmoid_f := 62;
        ELSIF x =- 7087 THEN
            sigmoid_f := 62;
        ELSIF x =- 7086 THEN
            sigmoid_f := 62;
        ELSIF x =- 7085 THEN
            sigmoid_f := 62;
        ELSIF x =- 7084 THEN
            sigmoid_f := 62;
        ELSIF x =- 7083 THEN
            sigmoid_f := 62;
        ELSIF x =- 7082 THEN
            sigmoid_f := 62;
        ELSIF x =- 7081 THEN
            sigmoid_f := 62;
        ELSIF x =- 7080 THEN
            sigmoid_f := 62;
        ELSIF x =- 7079 THEN
            sigmoid_f := 62;
        ELSIF x =- 7078 THEN
            sigmoid_f := 62;
        ELSIF x =- 7077 THEN
            sigmoid_f := 62;
        ELSIF x =- 7076 THEN
            sigmoid_f := 62;
        ELSIF x =- 7075 THEN
            sigmoid_f := 62;
        ELSIF x =- 7074 THEN
            sigmoid_f := 62;
        ELSIF x =- 7073 THEN
            sigmoid_f := 62;
        ELSIF x =- 7072 THEN
            sigmoid_f := 63;
        ELSIF x =- 7071 THEN
            sigmoid_f := 63;
        ELSIF x =- 7070 THEN
            sigmoid_f := 63;
        ELSIF x =- 7069 THEN
            sigmoid_f := 63;
        ELSIF x =- 7068 THEN
            sigmoid_f := 63;
        ELSIF x =- 7067 THEN
            sigmoid_f := 63;
        ELSIF x =- 7066 THEN
            sigmoid_f := 63;
        ELSIF x =- 7065 THEN
            sigmoid_f := 63;
        ELSIF x =- 7064 THEN
            sigmoid_f := 63;
        ELSIF x =- 7063 THEN
            sigmoid_f := 63;
        ELSIF x =- 7062 THEN
            sigmoid_f := 63;
        ELSIF x =- 7061 THEN
            sigmoid_f := 63;
        ELSIF x =- 7060 THEN
            sigmoid_f := 63;
        ELSIF x =- 7059 THEN
            sigmoid_f := 63;
        ELSIF x =- 7058 THEN
            sigmoid_f := 63;
        ELSIF x =- 7057 THEN
            sigmoid_f := 63;
        ELSIF x =- 7056 THEN
            sigmoid_f := 63;
        ELSIF x =- 7055 THEN
            sigmoid_f := 63;
        ELSIF x =- 7054 THEN
            sigmoid_f := 63;
        ELSIF x =- 7053 THEN
            sigmoid_f := 63;
        ELSIF x =- 7052 THEN
            sigmoid_f := 63;
        ELSIF x =- 7051 THEN
            sigmoid_f := 63;
        ELSIF x =- 7050 THEN
            sigmoid_f := 63;
        ELSIF x =- 7049 THEN
            sigmoid_f := 63;
        ELSIF x =- 7048 THEN
            sigmoid_f := 63;
        ELSIF x =- 7047 THEN
            sigmoid_f := 63;
        ELSIF x =- 7046 THEN
            sigmoid_f := 63;
        ELSIF x =- 7045 THEN
            sigmoid_f := 63;
        ELSIF x =- 7044 THEN
            sigmoid_f := 63;
        ELSIF x =- 7043 THEN
            sigmoid_f := 63;
        ELSIF x =- 7042 THEN
            sigmoid_f := 63;
        ELSIF x =- 7041 THEN
            sigmoid_f := 63;
        ELSIF x =- 7040 THEN
            sigmoid_f := 64;
        ELSIF x =- 7039 THEN
            sigmoid_f := 64;
        ELSIF x =- 7038 THEN
            sigmoid_f := 64;
        ELSIF x =- 7037 THEN
            sigmoid_f := 64;
        ELSIF x =- 7036 THEN
            sigmoid_f := 64;
        ELSIF x =- 7035 THEN
            sigmoid_f := 64;
        ELSIF x =- 7034 THEN
            sigmoid_f := 64;
        ELSIF x =- 7033 THEN
            sigmoid_f := 64;
        ELSIF x =- 7032 THEN
            sigmoid_f := 64;
        ELSIF x =- 7031 THEN
            sigmoid_f := 64;
        ELSIF x =- 7030 THEN
            sigmoid_f := 64;
        ELSIF x =- 7029 THEN
            sigmoid_f := 64;
        ELSIF x =- 7028 THEN
            sigmoid_f := 64;
        ELSIF x =- 7027 THEN
            sigmoid_f := 64;
        ELSIF x =- 7026 THEN
            sigmoid_f := 64;
        ELSIF x =- 7025 THEN
            sigmoid_f := 64;
        ELSIF x =- 7024 THEN
            sigmoid_f := 64;
        ELSIF x =- 7023 THEN
            sigmoid_f := 64;
        ELSIF x =- 7022 THEN
            sigmoid_f := 64;
        ELSIF x =- 7021 THEN
            sigmoid_f := 64;
        ELSIF x =- 7020 THEN
            sigmoid_f := 64;
        ELSIF x =- 7019 THEN
            sigmoid_f := 64;
        ELSIF x =- 7018 THEN
            sigmoid_f := 64;
        ELSIF x =- 7017 THEN
            sigmoid_f := 64;
        ELSIF x =- 7016 THEN
            sigmoid_f := 64;
        ELSIF x =- 7015 THEN
            sigmoid_f := 64;
        ELSIF x =- 7014 THEN
            sigmoid_f := 64;
        ELSIF x =- 7013 THEN
            sigmoid_f := 64;
        ELSIF x =- 7012 THEN
            sigmoid_f := 64;
        ELSIF x =- 7011 THEN
            sigmoid_f := 64;
        ELSIF x =- 7010 THEN
            sigmoid_f := 64;
        ELSIF x =- 7009 THEN
            sigmoid_f := 64;
        ELSIF x =- 7008 THEN
            sigmoid_f := 65;
        ELSIF x =- 7007 THEN
            sigmoid_f := 65;
        ELSIF x =- 7006 THEN
            sigmoid_f := 65;
        ELSIF x =- 7005 THEN
            sigmoid_f := 65;
        ELSIF x =- 7004 THEN
            sigmoid_f := 65;
        ELSIF x =- 7003 THEN
            sigmoid_f := 65;
        ELSIF x =- 7002 THEN
            sigmoid_f := 65;
        ELSIF x =- 7001 THEN
            sigmoid_f := 65;
        ELSIF x =- 7000 THEN
            sigmoid_f := 65;
        ELSIF x =- 6999 THEN
            sigmoid_f := 65;
        ELSIF x =- 6998 THEN
            sigmoid_f := 65;
        ELSIF x =- 6997 THEN
            sigmoid_f := 65;
        ELSIF x =- 6996 THEN
            sigmoid_f := 65;
        ELSIF x =- 6995 THEN
            sigmoid_f := 65;
        ELSIF x =- 6994 THEN
            sigmoid_f := 65;
        ELSIF x =- 6993 THEN
            sigmoid_f := 65;
        ELSIF x =- 6992 THEN
            sigmoid_f := 65;
        ELSIF x =- 6991 THEN
            sigmoid_f := 65;
        ELSIF x =- 6990 THEN
            sigmoid_f := 65;
        ELSIF x =- 6989 THEN
            sigmoid_f := 65;
        ELSIF x =- 6988 THEN
            sigmoid_f := 65;
        ELSIF x =- 6987 THEN
            sigmoid_f := 65;
        ELSIF x =- 6986 THEN
            sigmoid_f := 65;
        ELSIF x =- 6985 THEN
            sigmoid_f := 65;
        ELSIF x =- 6984 THEN
            sigmoid_f := 65;
        ELSIF x =- 6983 THEN
            sigmoid_f := 65;
        ELSIF x =- 6982 THEN
            sigmoid_f := 65;
        ELSIF x =- 6981 THEN
            sigmoid_f := 65;
        ELSIF x =- 6980 THEN
            sigmoid_f := 65;
        ELSIF x =- 6979 THEN
            sigmoid_f := 65;
        ELSIF x =- 6978 THEN
            sigmoid_f := 65;
        ELSIF x =- 6977 THEN
            sigmoid_f := 65;
        ELSIF x =- 6976 THEN
            sigmoid_f := 66;
        ELSIF x =- 6975 THEN
            sigmoid_f := 66;
        ELSIF x =- 6974 THEN
            sigmoid_f := 66;
        ELSIF x =- 6973 THEN
            sigmoid_f := 66;
        ELSIF x =- 6972 THEN
            sigmoid_f := 66;
        ELSIF x =- 6971 THEN
            sigmoid_f := 66;
        ELSIF x =- 6970 THEN
            sigmoid_f := 66;
        ELSIF x =- 6969 THEN
            sigmoid_f := 66;
        ELSIF x =- 6968 THEN
            sigmoid_f := 66;
        ELSIF x =- 6967 THEN
            sigmoid_f := 66;
        ELSIF x =- 6966 THEN
            sigmoid_f := 66;
        ELSIF x =- 6965 THEN
            sigmoid_f := 66;
        ELSIF x =- 6964 THEN
            sigmoid_f := 66;
        ELSIF x =- 6963 THEN
            sigmoid_f := 66;
        ELSIF x =- 6962 THEN
            sigmoid_f := 66;
        ELSIF x =- 6961 THEN
            sigmoid_f := 66;
        ELSIF x =- 6960 THEN
            sigmoid_f := 66;
        ELSIF x =- 6959 THEN
            sigmoid_f := 66;
        ELSIF x =- 6958 THEN
            sigmoid_f := 66;
        ELSIF x =- 6957 THEN
            sigmoid_f := 66;
        ELSIF x =- 6956 THEN
            sigmoid_f := 66;
        ELSIF x =- 6955 THEN
            sigmoid_f := 66;
        ELSIF x =- 6954 THEN
            sigmoid_f := 66;
        ELSIF x =- 6953 THEN
            sigmoid_f := 66;
        ELSIF x =- 6952 THEN
            sigmoid_f := 66;
        ELSIF x =- 6951 THEN
            sigmoid_f := 66;
        ELSIF x =- 6950 THEN
            sigmoid_f := 66;
        ELSIF x =- 6949 THEN
            sigmoid_f := 66;
        ELSIF x =- 6948 THEN
            sigmoid_f := 66;
        ELSIF x =- 6947 THEN
            sigmoid_f := 66;
        ELSIF x =- 6946 THEN
            sigmoid_f := 66;
        ELSIF x =- 6945 THEN
            sigmoid_f := 66;
        ELSIF x =- 6944 THEN
            sigmoid_f := 67;
        ELSIF x =- 6943 THEN
            sigmoid_f := 67;
        ELSIF x =- 6942 THEN
            sigmoid_f := 67;
        ELSIF x =- 6941 THEN
            sigmoid_f := 67;
        ELSIF x =- 6940 THEN
            sigmoid_f := 67;
        ELSIF x =- 6939 THEN
            sigmoid_f := 67;
        ELSIF x =- 6938 THEN
            sigmoid_f := 67;
        ELSIF x =- 6937 THEN
            sigmoid_f := 67;
        ELSIF x =- 6936 THEN
            sigmoid_f := 67;
        ELSIF x =- 6935 THEN
            sigmoid_f := 67;
        ELSIF x =- 6934 THEN
            sigmoid_f := 67;
        ELSIF x =- 6933 THEN
            sigmoid_f := 67;
        ELSIF x =- 6932 THEN
            sigmoid_f := 67;
        ELSIF x =- 6931 THEN
            sigmoid_f := 67;
        ELSIF x =- 6930 THEN
            sigmoid_f := 67;
        ELSIF x =- 6929 THEN
            sigmoid_f := 67;
        ELSIF x =- 6928 THEN
            sigmoid_f := 67;
        ELSIF x =- 6927 THEN
            sigmoid_f := 67;
        ELSIF x =- 6926 THEN
            sigmoid_f := 67;
        ELSIF x =- 6925 THEN
            sigmoid_f := 67;
        ELSIF x =- 6924 THEN
            sigmoid_f := 67;
        ELSIF x =- 6923 THEN
            sigmoid_f := 67;
        ELSIF x =- 6922 THEN
            sigmoid_f := 67;
        ELSIF x =- 6921 THEN
            sigmoid_f := 67;
        ELSIF x =- 6920 THEN
            sigmoid_f := 67;
        ELSIF x =- 6919 THEN
            sigmoid_f := 67;
        ELSIF x =- 6918 THEN
            sigmoid_f := 67;
        ELSIF x =- 6917 THEN
            sigmoid_f := 67;
        ELSIF x =- 6916 THEN
            sigmoid_f := 67;
        ELSIF x =- 6915 THEN
            sigmoid_f := 67;
        ELSIF x =- 6914 THEN
            sigmoid_f := 67;
        ELSIF x =- 6913 THEN
            sigmoid_f := 67;
        ELSIF x =- 6912 THEN
            sigmoid_f := 68;
        ELSIF x =- 6911 THEN
            sigmoid_f := 68;
        ELSIF x =- 6910 THEN
            sigmoid_f := 68;
        ELSIF x =- 6909 THEN
            sigmoid_f := 68;
        ELSIF x =- 6908 THEN
            sigmoid_f := 68;
        ELSIF x =- 6907 THEN
            sigmoid_f := 68;
        ELSIF x =- 6906 THEN
            sigmoid_f := 68;
        ELSIF x =- 6905 THEN
            sigmoid_f := 68;
        ELSIF x =- 6904 THEN
            sigmoid_f := 68;
        ELSIF x =- 6903 THEN
            sigmoid_f := 68;
        ELSIF x =- 6902 THEN
            sigmoid_f := 68;
        ELSIF x =- 6901 THEN
            sigmoid_f := 68;
        ELSIF x =- 6900 THEN
            sigmoid_f := 68;
        ELSIF x =- 6899 THEN
            sigmoid_f := 68;
        ELSIF x =- 6898 THEN
            sigmoid_f := 68;
        ELSIF x =- 6897 THEN
            sigmoid_f := 68;
        ELSIF x =- 6896 THEN
            sigmoid_f := 68;
        ELSIF x =- 6895 THEN
            sigmoid_f := 68;
        ELSIF x =- 6894 THEN
            sigmoid_f := 68;
        ELSIF x =- 6893 THEN
            sigmoid_f := 68;
        ELSIF x =- 6892 THEN
            sigmoid_f := 68;
        ELSIF x =- 6891 THEN
            sigmoid_f := 68;
        ELSIF x =- 6890 THEN
            sigmoid_f := 68;
        ELSIF x =- 6889 THEN
            sigmoid_f := 68;
        ELSIF x =- 6888 THEN
            sigmoid_f := 68;
        ELSIF x =- 6887 THEN
            sigmoid_f := 68;
        ELSIF x =- 6886 THEN
            sigmoid_f := 68;
        ELSIF x =- 6885 THEN
            sigmoid_f := 68;
        ELSIF x =- 6884 THEN
            sigmoid_f := 68;
        ELSIF x =- 6883 THEN
            sigmoid_f := 68;
        ELSIF x =- 6882 THEN
            sigmoid_f := 68;
        ELSIF x =- 6881 THEN
            sigmoid_f := 68;
        ELSIF x =- 6880 THEN
            sigmoid_f := 69;
        ELSIF x =- 6879 THEN
            sigmoid_f := 69;
        ELSIF x =- 6878 THEN
            sigmoid_f := 69;
        ELSIF x =- 6877 THEN
            sigmoid_f := 69;
        ELSIF x =- 6876 THEN
            sigmoid_f := 69;
        ELSIF x =- 6875 THEN
            sigmoid_f := 69;
        ELSIF x =- 6874 THEN
            sigmoid_f := 69;
        ELSIF x =- 6873 THEN
            sigmoid_f := 69;
        ELSIF x =- 6872 THEN
            sigmoid_f := 69;
        ELSIF x =- 6871 THEN
            sigmoid_f := 69;
        ELSIF x =- 6870 THEN
            sigmoid_f := 69;
        ELSIF x =- 6869 THEN
            sigmoid_f := 69;
        ELSIF x =- 6868 THEN
            sigmoid_f := 69;
        ELSIF x =- 6867 THEN
            sigmoid_f := 69;
        ELSIF x =- 6866 THEN
            sigmoid_f := 69;
        ELSIF x =- 6865 THEN
            sigmoid_f := 69;
        ELSIF x =- 6864 THEN
            sigmoid_f := 69;
        ELSIF x =- 6863 THEN
            sigmoid_f := 69;
        ELSIF x =- 6862 THEN
            sigmoid_f := 69;
        ELSIF x =- 6861 THEN
            sigmoid_f := 69;
        ELSIF x =- 6860 THEN
            sigmoid_f := 69;
        ELSIF x =- 6859 THEN
            sigmoid_f := 69;
        ELSIF x =- 6858 THEN
            sigmoid_f := 69;
        ELSIF x =- 6857 THEN
            sigmoid_f := 69;
        ELSIF x =- 6856 THEN
            sigmoid_f := 69;
        ELSIF x =- 6855 THEN
            sigmoid_f := 69;
        ELSIF x =- 6854 THEN
            sigmoid_f := 69;
        ELSIF x =- 6853 THEN
            sigmoid_f := 69;
        ELSIF x =- 6852 THEN
            sigmoid_f := 69;
        ELSIF x =- 6851 THEN
            sigmoid_f := 69;
        ELSIF x =- 6850 THEN
            sigmoid_f := 69;
        ELSIF x =- 6849 THEN
            sigmoid_f := 69;
        ELSIF x =- 6848 THEN
            sigmoid_f := 70;
        ELSIF x =- 6847 THEN
            sigmoid_f := 70;
        ELSIF x =- 6846 THEN
            sigmoid_f := 70;
        ELSIF x =- 6845 THEN
            sigmoid_f := 70;
        ELSIF x =- 6844 THEN
            sigmoid_f := 70;
        ELSIF x =- 6843 THEN
            sigmoid_f := 70;
        ELSIF x =- 6842 THEN
            sigmoid_f := 70;
        ELSIF x =- 6841 THEN
            sigmoid_f := 70;
        ELSIF x =- 6840 THEN
            sigmoid_f := 70;
        ELSIF x =- 6839 THEN
            sigmoid_f := 70;
        ELSIF x =- 6838 THEN
            sigmoid_f := 70;
        ELSIF x =- 6837 THEN
            sigmoid_f := 70;
        ELSIF x =- 6836 THEN
            sigmoid_f := 70;
        ELSIF x =- 6835 THEN
            sigmoid_f := 70;
        ELSIF x =- 6834 THEN
            sigmoid_f := 70;
        ELSIF x =- 6833 THEN
            sigmoid_f := 70;
        ELSIF x =- 6832 THEN
            sigmoid_f := 70;
        ELSIF x =- 6831 THEN
            sigmoid_f := 70;
        ELSIF x =- 6830 THEN
            sigmoid_f := 70;
        ELSIF x =- 6829 THEN
            sigmoid_f := 70;
        ELSIF x =- 6828 THEN
            sigmoid_f := 70;
        ELSIF x =- 6827 THEN
            sigmoid_f := 70;
        ELSIF x =- 6826 THEN
            sigmoid_f := 70;
        ELSIF x =- 6825 THEN
            sigmoid_f := 70;
        ELSIF x =- 6824 THEN
            sigmoid_f := 70;
        ELSIF x =- 6823 THEN
            sigmoid_f := 70;
        ELSIF x =- 6822 THEN
            sigmoid_f := 70;
        ELSIF x =- 6821 THEN
            sigmoid_f := 70;
        ELSIF x =- 6820 THEN
            sigmoid_f := 70;
        ELSIF x =- 6819 THEN
            sigmoid_f := 70;
        ELSIF x =- 6818 THEN
            sigmoid_f := 70;
        ELSIF x =- 6817 THEN
            sigmoid_f := 70;
        ELSIF x =- 6816 THEN
            sigmoid_f := 71;
        ELSIF x =- 6815 THEN
            sigmoid_f := 71;
        ELSIF x =- 6814 THEN
            sigmoid_f := 71;
        ELSIF x =- 6813 THEN
            sigmoid_f := 71;
        ELSIF x =- 6812 THEN
            sigmoid_f := 71;
        ELSIF x =- 6811 THEN
            sigmoid_f := 71;
        ELSIF x =- 6810 THEN
            sigmoid_f := 71;
        ELSIF x =- 6809 THEN
            sigmoid_f := 71;
        ELSIF x =- 6808 THEN
            sigmoid_f := 71;
        ELSIF x =- 6807 THEN
            sigmoid_f := 71;
        ELSIF x =- 6806 THEN
            sigmoid_f := 71;
        ELSIF x =- 6805 THEN
            sigmoid_f := 71;
        ELSIF x =- 6804 THEN
            sigmoid_f := 71;
        ELSIF x =- 6803 THEN
            sigmoid_f := 71;
        ELSIF x =- 6802 THEN
            sigmoid_f := 71;
        ELSIF x =- 6801 THEN
            sigmoid_f := 71;
        ELSIF x =- 6800 THEN
            sigmoid_f := 71;
        ELSIF x =- 6799 THEN
            sigmoid_f := 71;
        ELSIF x =- 6798 THEN
            sigmoid_f := 71;
        ELSIF x =- 6797 THEN
            sigmoid_f := 71;
        ELSIF x =- 6796 THEN
            sigmoid_f := 71;
        ELSIF x =- 6795 THEN
            sigmoid_f := 71;
        ELSIF x =- 6794 THEN
            sigmoid_f := 71;
        ELSIF x =- 6793 THEN
            sigmoid_f := 71;
        ELSIF x =- 6792 THEN
            sigmoid_f := 71;
        ELSIF x =- 6791 THEN
            sigmoid_f := 71;
        ELSIF x =- 6790 THEN
            sigmoid_f := 71;
        ELSIF x =- 6789 THEN
            sigmoid_f := 71;
        ELSIF x =- 6788 THEN
            sigmoid_f := 71;
        ELSIF x =- 6787 THEN
            sigmoid_f := 71;
        ELSIF x =- 6786 THEN
            sigmoid_f := 71;
        ELSIF x =- 6785 THEN
            sigmoid_f := 71;
        ELSIF x =- 6784 THEN
            sigmoid_f := 72;
        ELSIF x =- 6783 THEN
            sigmoid_f := 72;
        ELSIF x =- 6782 THEN
            sigmoid_f := 72;
        ELSIF x =- 6781 THEN
            sigmoid_f := 72;
        ELSIF x =- 6780 THEN
            sigmoid_f := 72;
        ELSIF x =- 6779 THEN
            sigmoid_f := 72;
        ELSIF x =- 6778 THEN
            sigmoid_f := 72;
        ELSIF x =- 6777 THEN
            sigmoid_f := 72;
        ELSIF x =- 6776 THEN
            sigmoid_f := 72;
        ELSIF x =- 6775 THEN
            sigmoid_f := 72;
        ELSIF x =- 6774 THEN
            sigmoid_f := 72;
        ELSIF x =- 6773 THEN
            sigmoid_f := 72;
        ELSIF x =- 6772 THEN
            sigmoid_f := 72;
        ELSIF x =- 6771 THEN
            sigmoid_f := 72;
        ELSIF x =- 6770 THEN
            sigmoid_f := 72;
        ELSIF x =- 6769 THEN
            sigmoid_f := 72;
        ELSIF x =- 6768 THEN
            sigmoid_f := 72;
        ELSIF x =- 6767 THEN
            sigmoid_f := 72;
        ELSIF x =- 6766 THEN
            sigmoid_f := 72;
        ELSIF x =- 6765 THEN
            sigmoid_f := 72;
        ELSIF x =- 6764 THEN
            sigmoid_f := 72;
        ELSIF x =- 6763 THEN
            sigmoid_f := 72;
        ELSIF x =- 6762 THEN
            sigmoid_f := 72;
        ELSIF x =- 6761 THEN
            sigmoid_f := 72;
        ELSIF x =- 6760 THEN
            sigmoid_f := 72;
        ELSIF x =- 6759 THEN
            sigmoid_f := 72;
        ELSIF x =- 6758 THEN
            sigmoid_f := 72;
        ELSIF x =- 6757 THEN
            sigmoid_f := 72;
        ELSIF x =- 6756 THEN
            sigmoid_f := 72;
        ELSIF x =- 6755 THEN
            sigmoid_f := 72;
        ELSIF x =- 6754 THEN
            sigmoid_f := 72;
        ELSIF x =- 6753 THEN
            sigmoid_f := 72;
        ELSIF x =- 6752 THEN
            sigmoid_f := 73;
        ELSIF x =- 6751 THEN
            sigmoid_f := 73;
        ELSIF x =- 6750 THEN
            sigmoid_f := 73;
        ELSIF x =- 6749 THEN
            sigmoid_f := 73;
        ELSIF x =- 6748 THEN
            sigmoid_f := 73;
        ELSIF x =- 6747 THEN
            sigmoid_f := 73;
        ELSIF x =- 6746 THEN
            sigmoid_f := 73;
        ELSIF x =- 6745 THEN
            sigmoid_f := 73;
        ELSIF x =- 6744 THEN
            sigmoid_f := 73;
        ELSIF x =- 6743 THEN
            sigmoid_f := 73;
        ELSIF x =- 6742 THEN
            sigmoid_f := 73;
        ELSIF x =- 6741 THEN
            sigmoid_f := 73;
        ELSIF x =- 6740 THEN
            sigmoid_f := 73;
        ELSIF x =- 6739 THEN
            sigmoid_f := 73;
        ELSIF x =- 6738 THEN
            sigmoid_f := 73;
        ELSIF x =- 6737 THEN
            sigmoid_f := 73;
        ELSIF x =- 6736 THEN
            sigmoid_f := 73;
        ELSIF x =- 6735 THEN
            sigmoid_f := 73;
        ELSIF x =- 6734 THEN
            sigmoid_f := 73;
        ELSIF x =- 6733 THEN
            sigmoid_f := 73;
        ELSIF x =- 6732 THEN
            sigmoid_f := 73;
        ELSIF x =- 6731 THEN
            sigmoid_f := 73;
        ELSIF x =- 6730 THEN
            sigmoid_f := 73;
        ELSIF x =- 6729 THEN
            sigmoid_f := 73;
        ELSIF x =- 6728 THEN
            sigmoid_f := 73;
        ELSIF x =- 6727 THEN
            sigmoid_f := 73;
        ELSIF x =- 6726 THEN
            sigmoid_f := 73;
        ELSIF x =- 6725 THEN
            sigmoid_f := 73;
        ELSIF x =- 6724 THEN
            sigmoid_f := 73;
        ELSIF x =- 6723 THEN
            sigmoid_f := 73;
        ELSIF x =- 6722 THEN
            sigmoid_f := 73;
        ELSIF x =- 6721 THEN
            sigmoid_f := 73;
        ELSIF x =- 6720 THEN
            sigmoid_f := 74;
        ELSIF x =- 6719 THEN
            sigmoid_f := 74;
        ELSIF x =- 6718 THEN
            sigmoid_f := 74;
        ELSIF x =- 6717 THEN
            sigmoid_f := 74;
        ELSIF x =- 6716 THEN
            sigmoid_f := 74;
        ELSIF x =- 6715 THEN
            sigmoid_f := 74;
        ELSIF x =- 6714 THEN
            sigmoid_f := 74;
        ELSIF x =- 6713 THEN
            sigmoid_f := 74;
        ELSIF x =- 6712 THEN
            sigmoid_f := 74;
        ELSIF x =- 6711 THEN
            sigmoid_f := 74;
        ELSIF x =- 6710 THEN
            sigmoid_f := 74;
        ELSIF x =- 6709 THEN
            sigmoid_f := 74;
        ELSIF x =- 6708 THEN
            sigmoid_f := 74;
        ELSIF x =- 6707 THEN
            sigmoid_f := 74;
        ELSIF x =- 6706 THEN
            sigmoid_f := 74;
        ELSIF x =- 6705 THEN
            sigmoid_f := 74;
        ELSIF x =- 6704 THEN
            sigmoid_f := 74;
        ELSIF x =- 6703 THEN
            sigmoid_f := 74;
        ELSIF x =- 6702 THEN
            sigmoid_f := 74;
        ELSIF x =- 6701 THEN
            sigmoid_f := 74;
        ELSIF x =- 6700 THEN
            sigmoid_f := 74;
        ELSIF x =- 6699 THEN
            sigmoid_f := 74;
        ELSIF x =- 6698 THEN
            sigmoid_f := 74;
        ELSIF x =- 6697 THEN
            sigmoid_f := 74;
        ELSIF x =- 6696 THEN
            sigmoid_f := 74;
        ELSIF x =- 6695 THEN
            sigmoid_f := 74;
        ELSIF x =- 6694 THEN
            sigmoid_f := 74;
        ELSIF x =- 6693 THEN
            sigmoid_f := 74;
        ELSIF x =- 6692 THEN
            sigmoid_f := 74;
        ELSIF x =- 6691 THEN
            sigmoid_f := 74;
        ELSIF x =- 6690 THEN
            sigmoid_f := 74;
        ELSIF x =- 6689 THEN
            sigmoid_f := 74;
        ELSIF x =- 6688 THEN
            sigmoid_f := 75;
        ELSIF x =- 6687 THEN
            sigmoid_f := 75;
        ELSIF x =- 6686 THEN
            sigmoid_f := 75;
        ELSIF x =- 6685 THEN
            sigmoid_f := 75;
        ELSIF x =- 6684 THEN
            sigmoid_f := 75;
        ELSIF x =- 6683 THEN
            sigmoid_f := 75;
        ELSIF x =- 6682 THEN
            sigmoid_f := 75;
        ELSIF x =- 6681 THEN
            sigmoid_f := 75;
        ELSIF x =- 6680 THEN
            sigmoid_f := 75;
        ELSIF x =- 6679 THEN
            sigmoid_f := 75;
        ELSIF x =- 6678 THEN
            sigmoid_f := 75;
        ELSIF x =- 6677 THEN
            sigmoid_f := 75;
        ELSIF x =- 6676 THEN
            sigmoid_f := 75;
        ELSIF x =- 6675 THEN
            sigmoid_f := 75;
        ELSIF x =- 6674 THEN
            sigmoid_f := 75;
        ELSIF x =- 6673 THEN
            sigmoid_f := 75;
        ELSIF x =- 6672 THEN
            sigmoid_f := 75;
        ELSIF x =- 6671 THEN
            sigmoid_f := 75;
        ELSIF x =- 6670 THEN
            sigmoid_f := 75;
        ELSIF x =- 6669 THEN
            sigmoid_f := 75;
        ELSIF x =- 6668 THEN
            sigmoid_f := 75;
        ELSIF x =- 6667 THEN
            sigmoid_f := 75;
        ELSIF x =- 6666 THEN
            sigmoid_f := 75;
        ELSIF x =- 6665 THEN
            sigmoid_f := 75;
        ELSIF x =- 6664 THEN
            sigmoid_f := 75;
        ELSIF x =- 6663 THEN
            sigmoid_f := 75;
        ELSIF x =- 6662 THEN
            sigmoid_f := 75;
        ELSIF x =- 6661 THEN
            sigmoid_f := 75;
        ELSIF x =- 6660 THEN
            sigmoid_f := 75;
        ELSIF x =- 6659 THEN
            sigmoid_f := 75;
        ELSIF x =- 6658 THEN
            sigmoid_f := 75;
        ELSIF x =- 6657 THEN
            sigmoid_f := 75;
        ELSIF x =- 6656 THEN
            sigmoid_f := 76;
        ELSIF x =- 6655 THEN
            sigmoid_f := 76;
        ELSIF x =- 6654 THEN
            sigmoid_f := 76;
        ELSIF x =- 6653 THEN
            sigmoid_f := 76;
        ELSIF x =- 6652 THEN
            sigmoid_f := 76;
        ELSIF x =- 6651 THEN
            sigmoid_f := 76;
        ELSIF x =- 6650 THEN
            sigmoid_f := 76;
        ELSIF x =- 6649 THEN
            sigmoid_f := 76;
        ELSIF x =- 6648 THEN
            sigmoid_f := 76;
        ELSIF x =- 6647 THEN
            sigmoid_f := 76;
        ELSIF x =- 6646 THEN
            sigmoid_f := 76;
        ELSIF x =- 6645 THEN
            sigmoid_f := 76;
        ELSIF x =- 6644 THEN
            sigmoid_f := 76;
        ELSIF x =- 6643 THEN
            sigmoid_f := 76;
        ELSIF x =- 6642 THEN
            sigmoid_f := 76;
        ELSIF x =- 6641 THEN
            sigmoid_f := 76;
        ELSIF x =- 6640 THEN
            sigmoid_f := 76;
        ELSIF x =- 6639 THEN
            sigmoid_f := 76;
        ELSIF x =- 6638 THEN
            sigmoid_f := 76;
        ELSIF x =- 6637 THEN
            sigmoid_f := 76;
        ELSIF x =- 6636 THEN
            sigmoid_f := 76;
        ELSIF x =- 6635 THEN
            sigmoid_f := 76;
        ELSIF x =- 6634 THEN
            sigmoid_f := 76;
        ELSIF x =- 6633 THEN
            sigmoid_f := 76;
        ELSIF x =- 6632 THEN
            sigmoid_f := 76;
        ELSIF x =- 6631 THEN
            sigmoid_f := 77;
        ELSIF x =- 6630 THEN
            sigmoid_f := 77;
        ELSIF x =- 6629 THEN
            sigmoid_f := 77;
        ELSIF x =- 6628 THEN
            sigmoid_f := 77;
        ELSIF x =- 6627 THEN
            sigmoid_f := 77;
        ELSIF x =- 6626 THEN
            sigmoid_f := 77;
        ELSIF x =- 6625 THEN
            sigmoid_f := 77;
        ELSIF x =- 6624 THEN
            sigmoid_f := 77;
        ELSIF x =- 6623 THEN
            sigmoid_f := 77;
        ELSIF x =- 6622 THEN
            sigmoid_f := 77;
        ELSIF x =- 6621 THEN
            sigmoid_f := 77;
        ELSIF x =- 6620 THEN
            sigmoid_f := 77;
        ELSIF x =- 6619 THEN
            sigmoid_f := 77;
        ELSIF x =- 6618 THEN
            sigmoid_f := 77;
        ELSIF x =- 6617 THEN
            sigmoid_f := 77;
        ELSIF x =- 6616 THEN
            sigmoid_f := 77;
        ELSIF x =- 6615 THEN
            sigmoid_f := 77;
        ELSIF x =- 6614 THEN
            sigmoid_f := 77;
        ELSIF x =- 6613 THEN
            sigmoid_f := 77;
        ELSIF x =- 6612 THEN
            sigmoid_f := 77;
        ELSIF x =- 6611 THEN
            sigmoid_f := 77;
        ELSIF x =- 6610 THEN
            sigmoid_f := 77;
        ELSIF x =- 6609 THEN
            sigmoid_f := 77;
        ELSIF x =- 6608 THEN
            sigmoid_f := 77;
        ELSIF x =- 6607 THEN
            sigmoid_f := 78;
        ELSIF x =- 6606 THEN
            sigmoid_f := 78;
        ELSIF x =- 6605 THEN
            sigmoid_f := 78;
        ELSIF x =- 6604 THEN
            sigmoid_f := 78;
        ELSIF x =- 6603 THEN
            sigmoid_f := 78;
        ELSIF x =- 6602 THEN
            sigmoid_f := 78;
        ELSIF x =- 6601 THEN
            sigmoid_f := 78;
        ELSIF x =- 6600 THEN
            sigmoid_f := 78;
        ELSIF x =- 6599 THEN
            sigmoid_f := 78;
        ELSIF x =- 6598 THEN
            sigmoid_f := 78;
        ELSIF x =- 6597 THEN
            sigmoid_f := 78;
        ELSIF x =- 6596 THEN
            sigmoid_f := 78;
        ELSIF x =- 6595 THEN
            sigmoid_f := 78;
        ELSIF x =- 6594 THEN
            sigmoid_f := 78;
        ELSIF x =- 6593 THEN
            sigmoid_f := 78;
        ELSIF x =- 6592 THEN
            sigmoid_f := 78;
        ELSIF x =- 6591 THEN
            sigmoid_f := 78;
        ELSIF x =- 6590 THEN
            sigmoid_f := 78;
        ELSIF x =- 6589 THEN
            sigmoid_f := 78;
        ELSIF x =- 6588 THEN
            sigmoid_f := 78;
        ELSIF x =- 6587 THEN
            sigmoid_f := 78;
        ELSIF x =- 6586 THEN
            sigmoid_f := 78;
        ELSIF x =- 6585 THEN
            sigmoid_f := 78;
        ELSIF x =- 6584 THEN
            sigmoid_f := 78;
        ELSIF x =- 6583 THEN
            sigmoid_f := 78;
        ELSIF x =- 6582 THEN
            sigmoid_f := 79;
        ELSIF x =- 6581 THEN
            sigmoid_f := 79;
        ELSIF x =- 6580 THEN
            sigmoid_f := 79;
        ELSIF x =- 6579 THEN
            sigmoid_f := 79;
        ELSIF x =- 6578 THEN
            sigmoid_f := 79;
        ELSIF x =- 6577 THEN
            sigmoid_f := 79;
        ELSIF x =- 6576 THEN
            sigmoid_f := 79;
        ELSIF x =- 6575 THEN
            sigmoid_f := 79;
        ELSIF x =- 6574 THEN
            sigmoid_f := 79;
        ELSIF x =- 6573 THEN
            sigmoid_f := 79;
        ELSIF x =- 6572 THEN
            sigmoid_f := 79;
        ELSIF x =- 6571 THEN
            sigmoid_f := 79;
        ELSIF x =- 6570 THEN
            sigmoid_f := 79;
        ELSIF x =- 6569 THEN
            sigmoid_f := 79;
        ELSIF x =- 6568 THEN
            sigmoid_f := 79;
        ELSIF x =- 6567 THEN
            sigmoid_f := 79;
        ELSIF x =- 6566 THEN
            sigmoid_f := 79;
        ELSIF x =- 6565 THEN
            sigmoid_f := 79;
        ELSIF x =- 6564 THEN
            sigmoid_f := 79;
        ELSIF x =- 6563 THEN
            sigmoid_f := 79;
        ELSIF x =- 6562 THEN
            sigmoid_f := 79;
        ELSIF x =- 6561 THEN
            sigmoid_f := 79;
        ELSIF x =- 6560 THEN
            sigmoid_f := 79;
        ELSIF x =- 6559 THEN
            sigmoid_f := 79;
        ELSIF x =- 6558 THEN
            sigmoid_f := 80;
        ELSIF x =- 6557 THEN
            sigmoid_f := 80;
        ELSIF x =- 6556 THEN
            sigmoid_f := 80;
        ELSIF x =- 6555 THEN
            sigmoid_f := 80;
        ELSIF x =- 6554 THEN
            sigmoid_f := 80;
        ELSIF x =- 6553 THEN
            sigmoid_f := 80;
        ELSIF x =- 6552 THEN
            sigmoid_f := 80;
        ELSIF x =- 6551 THEN
            sigmoid_f := 80;
        ELSIF x =- 6550 THEN
            sigmoid_f := 80;
        ELSIF x =- 6549 THEN
            sigmoid_f := 80;
        ELSIF x =- 6548 THEN
            sigmoid_f := 80;
        ELSIF x =- 6547 THEN
            sigmoid_f := 80;
        ELSIF x =- 6546 THEN
            sigmoid_f := 80;
        ELSIF x =- 6545 THEN
            sigmoid_f := 80;
        ELSIF x =- 6544 THEN
            sigmoid_f := 80;
        ELSIF x =- 6543 THEN
            sigmoid_f := 80;
        ELSIF x =- 6542 THEN
            sigmoid_f := 80;
        ELSIF x =- 6541 THEN
            sigmoid_f := 80;
        ELSIF x =- 6540 THEN
            sigmoid_f := 80;
        ELSIF x =- 6539 THEN
            sigmoid_f := 80;
        ELSIF x =- 6538 THEN
            sigmoid_f := 80;
        ELSIF x =- 6537 THEN
            sigmoid_f := 80;
        ELSIF x =- 6536 THEN
            sigmoid_f := 80;
        ELSIF x =- 6535 THEN
            sigmoid_f := 80;
        ELSIF x =- 6534 THEN
            sigmoid_f := 81;
        ELSIF x =- 6533 THEN
            sigmoid_f := 81;
        ELSIF x =- 6532 THEN
            sigmoid_f := 81;
        ELSIF x =- 6531 THEN
            sigmoid_f := 81;
        ELSIF x =- 6530 THEN
            sigmoid_f := 81;
        ELSIF x =- 6529 THEN
            sigmoid_f := 81;
        ELSIF x =- 6528 THEN
            sigmoid_f := 81;
        ELSIF x =- 6527 THEN
            sigmoid_f := 81;
        ELSIF x =- 6526 THEN
            sigmoid_f := 81;
        ELSIF x =- 6525 THEN
            sigmoid_f := 81;
        ELSIF x =- 6524 THEN
            sigmoid_f := 81;
        ELSIF x =- 6523 THEN
            sigmoid_f := 81;
        ELSIF x =- 6522 THEN
            sigmoid_f := 81;
        ELSIF x =- 6521 THEN
            sigmoid_f := 81;
        ELSIF x =- 6520 THEN
            sigmoid_f := 81;
        ELSIF x =- 6519 THEN
            sigmoid_f := 81;
        ELSIF x =- 6518 THEN
            sigmoid_f := 81;
        ELSIF x =- 6517 THEN
            sigmoid_f := 81;
        ELSIF x =- 6516 THEN
            sigmoid_f := 81;
        ELSIF x =- 6515 THEN
            sigmoid_f := 81;
        ELSIF x =- 6514 THEN
            sigmoid_f := 81;
        ELSIF x =- 6513 THEN
            sigmoid_f := 81;
        ELSIF x =- 6512 THEN
            sigmoid_f := 81;
        ELSIF x =- 6511 THEN
            sigmoid_f := 81;
        ELSIF x =- 6510 THEN
            sigmoid_f := 81;
        ELSIF x =- 6509 THEN
            sigmoid_f := 82;
        ELSIF x =- 6508 THEN
            sigmoid_f := 82;
        ELSIF x =- 6507 THEN
            sigmoid_f := 82;
        ELSIF x =- 6506 THEN
            sigmoid_f := 82;
        ELSIF x =- 6505 THEN
            sigmoid_f := 82;
        ELSIF x =- 6504 THEN
            sigmoid_f := 82;
        ELSIF x =- 6503 THEN
            sigmoid_f := 82;
        ELSIF x =- 6502 THEN
            sigmoid_f := 82;
        ELSIF x =- 6501 THEN
            sigmoid_f := 82;
        ELSIF x =- 6500 THEN
            sigmoid_f := 82;
        ELSIF x =- 6499 THEN
            sigmoid_f := 82;
        ELSIF x =- 6498 THEN
            sigmoid_f := 82;
        ELSIF x =- 6497 THEN
            sigmoid_f := 82;
        ELSIF x =- 6496 THEN
            sigmoid_f := 82;
        ELSIF x =- 6495 THEN
            sigmoid_f := 82;
        ELSIF x =- 6494 THEN
            sigmoid_f := 82;
        ELSIF x =- 6493 THEN
            sigmoid_f := 82;
        ELSIF x =- 6492 THEN
            sigmoid_f := 82;
        ELSIF x =- 6491 THEN
            sigmoid_f := 82;
        ELSIF x =- 6490 THEN
            sigmoid_f := 82;
        ELSIF x =- 6489 THEN
            sigmoid_f := 82;
        ELSIF x =- 6488 THEN
            sigmoid_f := 82;
        ELSIF x =- 6487 THEN
            sigmoid_f := 82;
        ELSIF x =- 6486 THEN
            sigmoid_f := 82;
        ELSIF x =- 6485 THEN
            sigmoid_f := 83;
        ELSIF x =- 6484 THEN
            sigmoid_f := 83;
        ELSIF x =- 6483 THEN
            sigmoid_f := 83;
        ELSIF x =- 6482 THEN
            sigmoid_f := 83;
        ELSIF x =- 6481 THEN
            sigmoid_f := 83;
        ELSIF x =- 6480 THEN
            sigmoid_f := 83;
        ELSIF x =- 6479 THEN
            sigmoid_f := 83;
        ELSIF x =- 6478 THEN
            sigmoid_f := 83;
        ELSIF x =- 6477 THEN
            sigmoid_f := 83;
        ELSIF x =- 6476 THEN
            sigmoid_f := 83;
        ELSIF x =- 6475 THEN
            sigmoid_f := 83;
        ELSIF x =- 6474 THEN
            sigmoid_f := 83;
        ELSIF x =- 6473 THEN
            sigmoid_f := 83;
        ELSIF x =- 6472 THEN
            sigmoid_f := 83;
        ELSIF x =- 6471 THEN
            sigmoid_f := 83;
        ELSIF x =- 6470 THEN
            sigmoid_f := 83;
        ELSIF x =- 6469 THEN
            sigmoid_f := 83;
        ELSIF x =- 6468 THEN
            sigmoid_f := 83;
        ELSIF x =- 6467 THEN
            sigmoid_f := 83;
        ELSIF x =- 6466 THEN
            sigmoid_f := 83;
        ELSIF x =- 6465 THEN
            sigmoid_f := 83;
        ELSIF x =- 6464 THEN
            sigmoid_f := 83;
        ELSIF x =- 6463 THEN
            sigmoid_f := 83;
        ELSIF x =- 6462 THEN
            sigmoid_f := 83;
        ELSIF x =- 6461 THEN
            sigmoid_f := 83;
        ELSIF x =- 6460 THEN
            sigmoid_f := 84;
        ELSIF x =- 6459 THEN
            sigmoid_f := 84;
        ELSIF x =- 6458 THEN
            sigmoid_f := 84;
        ELSIF x =- 6457 THEN
            sigmoid_f := 84;
        ELSIF x =- 6456 THEN
            sigmoid_f := 84;
        ELSIF x =- 6455 THEN
            sigmoid_f := 84;
        ELSIF x =- 6454 THEN
            sigmoid_f := 84;
        ELSIF x =- 6453 THEN
            sigmoid_f := 84;
        ELSIF x =- 6452 THEN
            sigmoid_f := 84;
        ELSIF x =- 6451 THEN
            sigmoid_f := 84;
        ELSIF x =- 6450 THEN
            sigmoid_f := 84;
        ELSIF x =- 6449 THEN
            sigmoid_f := 84;
        ELSIF x =- 6448 THEN
            sigmoid_f := 84;
        ELSIF x =- 6447 THEN
            sigmoid_f := 84;
        ELSIF x =- 6446 THEN
            sigmoid_f := 84;
        ELSIF x =- 6445 THEN
            sigmoid_f := 84;
        ELSIF x =- 6444 THEN
            sigmoid_f := 84;
        ELSIF x =- 6443 THEN
            sigmoid_f := 84;
        ELSIF x =- 6442 THEN
            sigmoid_f := 84;
        ELSIF x =- 6441 THEN
            sigmoid_f := 84;
        ELSIF x =- 6440 THEN
            sigmoid_f := 84;
        ELSIF x =- 6439 THEN
            sigmoid_f := 84;
        ELSIF x =- 6438 THEN
            sigmoid_f := 84;
        ELSIF x =- 6437 THEN
            sigmoid_f := 84;
        ELSIF x =- 6436 THEN
            sigmoid_f := 85;
        ELSIF x =- 6435 THEN
            sigmoid_f := 85;
        ELSIF x =- 6434 THEN
            sigmoid_f := 85;
        ELSIF x =- 6433 THEN
            sigmoid_f := 85;
        ELSIF x =- 6432 THEN
            sigmoid_f := 85;
        ELSIF x =- 6431 THEN
            sigmoid_f := 85;
        ELSIF x =- 6430 THEN
            sigmoid_f := 85;
        ELSIF x =- 6429 THEN
            sigmoid_f := 85;
        ELSIF x =- 6428 THEN
            sigmoid_f := 85;
        ELSIF x =- 6427 THEN
            sigmoid_f := 85;
        ELSIF x =- 6426 THEN
            sigmoid_f := 85;
        ELSIF x =- 6425 THEN
            sigmoid_f := 85;
        ELSIF x =- 6424 THEN
            sigmoid_f := 85;
        ELSIF x =- 6423 THEN
            sigmoid_f := 85;
        ELSIF x =- 6422 THEN
            sigmoid_f := 85;
        ELSIF x =- 6421 THEN
            sigmoid_f := 85;
        ELSIF x =- 6420 THEN
            sigmoid_f := 85;
        ELSIF x =- 6419 THEN
            sigmoid_f := 85;
        ELSIF x =- 6418 THEN
            sigmoid_f := 85;
        ELSIF x =- 6417 THEN
            sigmoid_f := 85;
        ELSIF x =- 6416 THEN
            sigmoid_f := 85;
        ELSIF x =- 6415 THEN
            sigmoid_f := 85;
        ELSIF x =- 6414 THEN
            sigmoid_f := 85;
        ELSIF x =- 6413 THEN
            sigmoid_f := 85;
        ELSIF x =- 6412 THEN
            sigmoid_f := 86;
        ELSIF x =- 6411 THEN
            sigmoid_f := 86;
        ELSIF x =- 6410 THEN
            sigmoid_f := 86;
        ELSIF x =- 6409 THEN
            sigmoid_f := 86;
        ELSIF x =- 6408 THEN
            sigmoid_f := 86;
        ELSIF x =- 6407 THEN
            sigmoid_f := 86;
        ELSIF x =- 6406 THEN
            sigmoid_f := 86;
        ELSIF x =- 6405 THEN
            sigmoid_f := 86;
        ELSIF x =- 6404 THEN
            sigmoid_f := 86;
        ELSIF x =- 6403 THEN
            sigmoid_f := 86;
        ELSIF x =- 6402 THEN
            sigmoid_f := 86;
        ELSIF x =- 6401 THEN
            sigmoid_f := 86;
        ELSIF x =- 6400 THEN
            sigmoid_f := 86;
        ELSIF x =- 6399 THEN
            sigmoid_f := 86;
        ELSIF x =- 6398 THEN
            sigmoid_f := 86;
        ELSIF x =- 6397 THEN
            sigmoid_f := 86;
        ELSIF x =- 6396 THEN
            sigmoid_f := 86;
        ELSIF x =- 6395 THEN
            sigmoid_f := 86;
        ELSIF x =- 6394 THEN
            sigmoid_f := 86;
        ELSIF x =- 6393 THEN
            sigmoid_f := 86;
        ELSIF x =- 6392 THEN
            sigmoid_f := 86;
        ELSIF x =- 6391 THEN
            sigmoid_f := 86;
        ELSIF x =- 6390 THEN
            sigmoid_f := 86;
        ELSIF x =- 6389 THEN
            sigmoid_f := 86;
        ELSIF x =- 6388 THEN
            sigmoid_f := 86;
        ELSIF x =- 6387 THEN
            sigmoid_f := 87;
        ELSIF x =- 6386 THEN
            sigmoid_f := 87;
        ELSIF x =- 6385 THEN
            sigmoid_f := 87;
        ELSIF x =- 6384 THEN
            sigmoid_f := 87;
        ELSIF x =- 6383 THEN
            sigmoid_f := 87;
        ELSIF x =- 6382 THEN
            sigmoid_f := 87;
        ELSIF x =- 6381 THEN
            sigmoid_f := 87;
        ELSIF x =- 6380 THEN
            sigmoid_f := 87;
        ELSIF x =- 6379 THEN
            sigmoid_f := 87;
        ELSIF x =- 6378 THEN
            sigmoid_f := 87;
        ELSIF x =- 6377 THEN
            sigmoid_f := 87;
        ELSIF x =- 6376 THEN
            sigmoid_f := 87;
        ELSIF x =- 6375 THEN
            sigmoid_f := 87;
        ELSIF x =- 6374 THEN
            sigmoid_f := 87;
        ELSIF x =- 6373 THEN
            sigmoid_f := 87;
        ELSIF x =- 6372 THEN
            sigmoid_f := 87;
        ELSIF x =- 6371 THEN
            sigmoid_f := 87;
        ELSIF x =- 6370 THEN
            sigmoid_f := 87;
        ELSIF x =- 6369 THEN
            sigmoid_f := 87;
        ELSIF x =- 6368 THEN
            sigmoid_f := 87;
        ELSIF x =- 6367 THEN
            sigmoid_f := 87;
        ELSIF x =- 6366 THEN
            sigmoid_f := 87;
        ELSIF x =- 6365 THEN
            sigmoid_f := 87;
        ELSIF x =- 6364 THEN
            sigmoid_f := 87;
        ELSIF x =- 6363 THEN
            sigmoid_f := 88;
        ELSIF x =- 6362 THEN
            sigmoid_f := 88;
        ELSIF x =- 6361 THEN
            sigmoid_f := 88;
        ELSIF x =- 6360 THEN
            sigmoid_f := 88;
        ELSIF x =- 6359 THEN
            sigmoid_f := 88;
        ELSIF x =- 6358 THEN
            sigmoid_f := 88;
        ELSIF x =- 6357 THEN
            sigmoid_f := 88;
        ELSIF x =- 6356 THEN
            sigmoid_f := 88;
        ELSIF x =- 6355 THEN
            sigmoid_f := 88;
        ELSIF x =- 6354 THEN
            sigmoid_f := 88;
        ELSIF x =- 6353 THEN
            sigmoid_f := 88;
        ELSIF x =- 6352 THEN
            sigmoid_f := 88;
        ELSIF x =- 6351 THEN
            sigmoid_f := 88;
        ELSIF x =- 6350 THEN
            sigmoid_f := 88;
        ELSIF x =- 6349 THEN
            sigmoid_f := 88;
        ELSIF x =- 6348 THEN
            sigmoid_f := 88;
        ELSIF x =- 6347 THEN
            sigmoid_f := 88;
        ELSIF x =- 6346 THEN
            sigmoid_f := 88;
        ELSIF x =- 6345 THEN
            sigmoid_f := 88;
        ELSIF x =- 6344 THEN
            sigmoid_f := 88;
        ELSIF x =- 6343 THEN
            sigmoid_f := 88;
        ELSIF x =- 6342 THEN
            sigmoid_f := 88;
        ELSIF x =- 6341 THEN
            sigmoid_f := 88;
        ELSIF x =- 6340 THEN
            sigmoid_f := 88;
        ELSIF x =- 6339 THEN
            sigmoid_f := 89;
        ELSIF x =- 6338 THEN
            sigmoid_f := 89;
        ELSIF x =- 6337 THEN
            sigmoid_f := 89;
        ELSIF x =- 6336 THEN
            sigmoid_f := 89;
        ELSIF x =- 6335 THEN
            sigmoid_f := 89;
        ELSIF x =- 6334 THEN
            sigmoid_f := 89;
        ELSIF x =- 6333 THEN
            sigmoid_f := 89;
        ELSIF x =- 6332 THEN
            sigmoid_f := 89;
        ELSIF x =- 6331 THEN
            sigmoid_f := 89;
        ELSIF x =- 6330 THEN
            sigmoid_f := 89;
        ELSIF x =- 6329 THEN
            sigmoid_f := 89;
        ELSIF x =- 6328 THEN
            sigmoid_f := 89;
        ELSIF x =- 6327 THEN
            sigmoid_f := 89;
        ELSIF x =- 6326 THEN
            sigmoid_f := 89;
        ELSIF x =- 6325 THEN
            sigmoid_f := 89;
        ELSIF x =- 6324 THEN
            sigmoid_f := 89;
        ELSIF x =- 6323 THEN
            sigmoid_f := 89;
        ELSIF x =- 6322 THEN
            sigmoid_f := 89;
        ELSIF x =- 6321 THEN
            sigmoid_f := 89;
        ELSIF x =- 6320 THEN
            sigmoid_f := 89;
        ELSIF x =- 6319 THEN
            sigmoid_f := 89;
        ELSIF x =- 6318 THEN
            sigmoid_f := 89;
        ELSIF x =- 6317 THEN
            sigmoid_f := 89;
        ELSIF x =- 6316 THEN
            sigmoid_f := 89;
        ELSIF x =- 6315 THEN
            sigmoid_f := 89;
        ELSIF x =- 6314 THEN
            sigmoid_f := 90;
        ELSIF x =- 6313 THEN
            sigmoid_f := 90;
        ELSIF x =- 6312 THEN
            sigmoid_f := 90;
        ELSIF x =- 6311 THEN
            sigmoid_f := 90;
        ELSIF x =- 6310 THEN
            sigmoid_f := 90;
        ELSIF x =- 6309 THEN
            sigmoid_f := 90;
        ELSIF x =- 6308 THEN
            sigmoid_f := 90;
        ELSIF x =- 6307 THEN
            sigmoid_f := 90;
        ELSIF x =- 6306 THEN
            sigmoid_f := 90;
        ELSIF x =- 6305 THEN
            sigmoid_f := 90;
        ELSIF x =- 6304 THEN
            sigmoid_f := 90;
        ELSIF x =- 6303 THEN
            sigmoid_f := 90;
        ELSIF x =- 6302 THEN
            sigmoid_f := 90;
        ELSIF x =- 6301 THEN
            sigmoid_f := 90;
        ELSIF x =- 6300 THEN
            sigmoid_f := 90;
        ELSIF x =- 6299 THEN
            sigmoid_f := 90;
        ELSIF x =- 6298 THEN
            sigmoid_f := 90;
        ELSIF x =- 6297 THEN
            sigmoid_f := 90;
        ELSIF x =- 6296 THEN
            sigmoid_f := 90;
        ELSIF x =- 6295 THEN
            sigmoid_f := 90;
        ELSIF x =- 6294 THEN
            sigmoid_f := 90;
        ELSIF x =- 6293 THEN
            sigmoid_f := 90;
        ELSIF x =- 6292 THEN
            sigmoid_f := 90;
        ELSIF x =- 6291 THEN
            sigmoid_f := 90;
        ELSIF x =- 6290 THEN
            sigmoid_f := 91;
        ELSIF x =- 6289 THEN
            sigmoid_f := 91;
        ELSIF x =- 6288 THEN
            sigmoid_f := 91;
        ELSIF x =- 6287 THEN
            sigmoid_f := 91;
        ELSIF x =- 6286 THEN
            sigmoid_f := 91;
        ELSIF x =- 6285 THEN
            sigmoid_f := 91;
        ELSIF x =- 6284 THEN
            sigmoid_f := 91;
        ELSIF x =- 6283 THEN
            sigmoid_f := 91;
        ELSIF x =- 6282 THEN
            sigmoid_f := 91;
        ELSIF x =- 6281 THEN
            sigmoid_f := 91;
        ELSIF x =- 6280 THEN
            sigmoid_f := 91;
        ELSIF x =- 6279 THEN
            sigmoid_f := 91;
        ELSIF x =- 6278 THEN
            sigmoid_f := 91;
        ELSIF x =- 6277 THEN
            sigmoid_f := 91;
        ELSIF x =- 6276 THEN
            sigmoid_f := 91;
        ELSIF x =- 6275 THEN
            sigmoid_f := 91;
        ELSIF x =- 6274 THEN
            sigmoid_f := 91;
        ELSIF x =- 6273 THEN
            sigmoid_f := 91;
        ELSIF x =- 6272 THEN
            sigmoid_f := 91;
        ELSIF x =- 6271 THEN
            sigmoid_f := 91;
        ELSIF x =- 6270 THEN
            sigmoid_f := 91;
        ELSIF x =- 6269 THEN
            sigmoid_f := 91;
        ELSIF x =- 6268 THEN
            sigmoid_f := 91;
        ELSIF x =- 6267 THEN
            sigmoid_f := 91;
        ELSIF x =- 6266 THEN
            sigmoid_f := 91;
        ELSIF x =- 6265 THEN
            sigmoid_f := 92;
        ELSIF x =- 6264 THEN
            sigmoid_f := 92;
        ELSIF x =- 6263 THEN
            sigmoid_f := 92;
        ELSIF x =- 6262 THEN
            sigmoid_f := 92;
        ELSIF x =- 6261 THEN
            sigmoid_f := 92;
        ELSIF x =- 6260 THEN
            sigmoid_f := 92;
        ELSIF x =- 6259 THEN
            sigmoid_f := 92;
        ELSIF x =- 6258 THEN
            sigmoid_f := 92;
        ELSIF x =- 6257 THEN
            sigmoid_f := 92;
        ELSIF x =- 6256 THEN
            sigmoid_f := 92;
        ELSIF x =- 6255 THEN
            sigmoid_f := 92;
        ELSIF x =- 6254 THEN
            sigmoid_f := 92;
        ELSIF x =- 6253 THEN
            sigmoid_f := 92;
        ELSIF x =- 6252 THEN
            sigmoid_f := 92;
        ELSIF x =- 6251 THEN
            sigmoid_f := 92;
        ELSIF x =- 6250 THEN
            sigmoid_f := 92;
        ELSIF x =- 6249 THEN
            sigmoid_f := 92;
        ELSIF x =- 6248 THEN
            sigmoid_f := 92;
        ELSIF x =- 6247 THEN
            sigmoid_f := 92;
        ELSIF x =- 6246 THEN
            sigmoid_f := 92;
        ELSIF x =- 6245 THEN
            sigmoid_f := 92;
        ELSIF x =- 6244 THEN
            sigmoid_f := 92;
        ELSIF x =- 6243 THEN
            sigmoid_f := 92;
        ELSIF x =- 6242 THEN
            sigmoid_f := 92;
        ELSIF x =- 6241 THEN
            sigmoid_f := 93;
        ELSIF x =- 6240 THEN
            sigmoid_f := 93;
        ELSIF x =- 6239 THEN
            sigmoid_f := 93;
        ELSIF x =- 6238 THEN
            sigmoid_f := 93;
        ELSIF x =- 6237 THEN
            sigmoid_f := 93;
        ELSIF x =- 6236 THEN
            sigmoid_f := 93;
        ELSIF x =- 6235 THEN
            sigmoid_f := 93;
        ELSIF x =- 6234 THEN
            sigmoid_f := 93;
        ELSIF x =- 6233 THEN
            sigmoid_f := 93;
        ELSIF x =- 6232 THEN
            sigmoid_f := 93;
        ELSIF x =- 6231 THEN
            sigmoid_f := 93;
        ELSIF x =- 6230 THEN
            sigmoid_f := 93;
        ELSIF x =- 6229 THEN
            sigmoid_f := 93;
        ELSIF x =- 6228 THEN
            sigmoid_f := 93;
        ELSIF x =- 6227 THEN
            sigmoid_f := 93;
        ELSIF x =- 6226 THEN
            sigmoid_f := 93;
        ELSIF x =- 6225 THEN
            sigmoid_f := 93;
        ELSIF x =- 6224 THEN
            sigmoid_f := 93;
        ELSIF x =- 6223 THEN
            sigmoid_f := 93;
        ELSIF x =- 6222 THEN
            sigmoid_f := 93;
        ELSIF x =- 6221 THEN
            sigmoid_f := 93;
        ELSIF x =- 6220 THEN
            sigmoid_f := 93;
        ELSIF x =- 6219 THEN
            sigmoid_f := 93;
        ELSIF x =- 6218 THEN
            sigmoid_f := 93;
        ELSIF x =- 6217 THEN
            sigmoid_f := 94;
        ELSIF x =- 6216 THEN
            sigmoid_f := 94;
        ELSIF x =- 6215 THEN
            sigmoid_f := 94;
        ELSIF x =- 6214 THEN
            sigmoid_f := 94;
        ELSIF x =- 6213 THEN
            sigmoid_f := 94;
        ELSIF x =- 6212 THEN
            sigmoid_f := 94;
        ELSIF x =- 6211 THEN
            sigmoid_f := 94;
        ELSIF x =- 6210 THEN
            sigmoid_f := 94;
        ELSIF x =- 6209 THEN
            sigmoid_f := 94;
        ELSIF x =- 6208 THEN
            sigmoid_f := 94;
        ELSIF x =- 6207 THEN
            sigmoid_f := 94;
        ELSIF x =- 6206 THEN
            sigmoid_f := 94;
        ELSIF x =- 6205 THEN
            sigmoid_f := 94;
        ELSIF x =- 6204 THEN
            sigmoid_f := 94;
        ELSIF x =- 6203 THEN
            sigmoid_f := 94;
        ELSIF x =- 6202 THEN
            sigmoid_f := 94;
        ELSIF x =- 6201 THEN
            sigmoid_f := 94;
        ELSIF x =- 6200 THEN
            sigmoid_f := 94;
        ELSIF x =- 6199 THEN
            sigmoid_f := 94;
        ELSIF x =- 6198 THEN
            sigmoid_f := 94;
        ELSIF x =- 6197 THEN
            sigmoid_f := 94;
        ELSIF x =- 6196 THEN
            sigmoid_f := 94;
        ELSIF x =- 6195 THEN
            sigmoid_f := 94;
        ELSIF x =- 6194 THEN
            sigmoid_f := 94;
        ELSIF x =- 6193 THEN
            sigmoid_f := 94;
        ELSIF x =- 6192 THEN
            sigmoid_f := 95;
        ELSIF x =- 6191 THEN
            sigmoid_f := 95;
        ELSIF x =- 6190 THEN
            sigmoid_f := 95;
        ELSIF x =- 6189 THEN
            sigmoid_f := 95;
        ELSIF x =- 6188 THEN
            sigmoid_f := 95;
        ELSIF x =- 6187 THEN
            sigmoid_f := 95;
        ELSIF x =- 6186 THEN
            sigmoid_f := 95;
        ELSIF x =- 6185 THEN
            sigmoid_f := 95;
        ELSIF x =- 6184 THEN
            sigmoid_f := 95;
        ELSIF x =- 6183 THEN
            sigmoid_f := 95;
        ELSIF x =- 6182 THEN
            sigmoid_f := 95;
        ELSIF x =- 6181 THEN
            sigmoid_f := 95;
        ELSIF x =- 6180 THEN
            sigmoid_f := 95;
        ELSIF x =- 6179 THEN
            sigmoid_f := 95;
        ELSIF x =- 6178 THEN
            sigmoid_f := 95;
        ELSIF x =- 6177 THEN
            sigmoid_f := 95;
        ELSIF x =- 6176 THEN
            sigmoid_f := 95;
        ELSIF x =- 6175 THEN
            sigmoid_f := 95;
        ELSIF x =- 6174 THEN
            sigmoid_f := 95;
        ELSIF x =- 6173 THEN
            sigmoid_f := 95;
        ELSIF x =- 6172 THEN
            sigmoid_f := 95;
        ELSIF x =- 6171 THEN
            sigmoid_f := 95;
        ELSIF x =- 6170 THEN
            sigmoid_f := 95;
        ELSIF x =- 6169 THEN
            sigmoid_f := 95;
        ELSIF x =- 6168 THEN
            sigmoid_f := 96;
        ELSIF x =- 6167 THEN
            sigmoid_f := 96;
        ELSIF x =- 6166 THEN
            sigmoid_f := 96;
        ELSIF x =- 6165 THEN
            sigmoid_f := 96;
        ELSIF x =- 6164 THEN
            sigmoid_f := 96;
        ELSIF x =- 6163 THEN
            sigmoid_f := 96;
        ELSIF x =- 6162 THEN
            sigmoid_f := 96;
        ELSIF x =- 6161 THEN
            sigmoid_f := 96;
        ELSIF x =- 6160 THEN
            sigmoid_f := 96;
        ELSIF x =- 6159 THEN
            sigmoid_f := 96;
        ELSIF x =- 6158 THEN
            sigmoid_f := 96;
        ELSIF x =- 6157 THEN
            sigmoid_f := 96;
        ELSIF x =- 6156 THEN
            sigmoid_f := 96;
        ELSIF x =- 6155 THEN
            sigmoid_f := 96;
        ELSIF x =- 6154 THEN
            sigmoid_f := 96;
        ELSIF x =- 6153 THEN
            sigmoid_f := 96;
        ELSIF x =- 6152 THEN
            sigmoid_f := 96;
        ELSIF x =- 6151 THEN
            sigmoid_f := 96;
        ELSIF x =- 6150 THEN
            sigmoid_f := 96;
        ELSIF x =- 6149 THEN
            sigmoid_f := 96;
        ELSIF x =- 6148 THEN
            sigmoid_f := 96;
        ELSIF x =- 6147 THEN
            sigmoid_f := 96;
        ELSIF x =- 6146 THEN
            sigmoid_f := 96;
        ELSIF x =- 6145 THEN
            sigmoid_f := 96;
        ELSIF x =- 6144 THEN
            sigmoid_f := 97;
        ELSIF x =- 6143 THEN
            sigmoid_f := 97;
        ELSIF x =- 6142 THEN
            sigmoid_f := 97;
        ELSIF x =- 6141 THEN
            sigmoid_f := 97;
        ELSIF x =- 6140 THEN
            sigmoid_f := 97;
        ELSIF x =- 6139 THEN
            sigmoid_f := 97;
        ELSIF x =- 6138 THEN
            sigmoid_f := 97;
        ELSIF x =- 6137 THEN
            sigmoid_f := 97;
        ELSIF x =- 6136 THEN
            sigmoid_f := 97;
        ELSIF x =- 6135 THEN
            sigmoid_f := 97;
        ELSIF x =- 6134 THEN
            sigmoid_f := 97;
        ELSIF x =- 6133 THEN
            sigmoid_f := 97;
        ELSIF x =- 6132 THEN
            sigmoid_f := 97;
        ELSIF x =- 6131 THEN
            sigmoid_f := 97;
        ELSIF x =- 6130 THEN
            sigmoid_f := 97;
        ELSIF x =- 6129 THEN
            sigmoid_f := 97;
        ELSIF x =- 6128 THEN
            sigmoid_f := 97;
        ELSIF x =- 6127 THEN
            sigmoid_f := 97;
        ELSIF x =- 6126 THEN
            sigmoid_f := 97;
        ELSIF x =- 6125 THEN
            sigmoid_f := 97;
        ELSIF x =- 6124 THEN
            sigmoid_f := 97;
        ELSIF x =- 6123 THEN
            sigmoid_f := 98;
        ELSIF x =- 6122 THEN
            sigmoid_f := 98;
        ELSIF x =- 6121 THEN
            sigmoid_f := 98;
        ELSIF x =- 6120 THEN
            sigmoid_f := 98;
        ELSIF x =- 6119 THEN
            sigmoid_f := 98;
        ELSIF x =- 6118 THEN
            sigmoid_f := 98;
        ELSIF x =- 6117 THEN
            sigmoid_f := 98;
        ELSIF x =- 6116 THEN
            sigmoid_f := 98;
        ELSIF x =- 6115 THEN
            sigmoid_f := 98;
        ELSIF x =- 6114 THEN
            sigmoid_f := 98;
        ELSIF x =- 6113 THEN
            sigmoid_f := 98;
        ELSIF x =- 6112 THEN
            sigmoid_f := 98;
        ELSIF x =- 6111 THEN
            sigmoid_f := 98;
        ELSIF x =- 6110 THEN
            sigmoid_f := 98;
        ELSIF x =- 6109 THEN
            sigmoid_f := 98;
        ELSIF x =- 6108 THEN
            sigmoid_f := 98;
        ELSIF x =- 6107 THEN
            sigmoid_f := 98;
        ELSIF x =- 6106 THEN
            sigmoid_f := 98;
        ELSIF x =- 6105 THEN
            sigmoid_f := 98;
        ELSIF x =- 6104 THEN
            sigmoid_f := 98;
        ELSIF x =- 6103 THEN
            sigmoid_f := 99;
        ELSIF x =- 6102 THEN
            sigmoid_f := 99;
        ELSIF x =- 6101 THEN
            sigmoid_f := 99;
        ELSIF x =- 6100 THEN
            sigmoid_f := 99;
        ELSIF x =- 6099 THEN
            sigmoid_f := 99;
        ELSIF x =- 6098 THEN
            sigmoid_f := 99;
        ELSIF x =- 6097 THEN
            sigmoid_f := 99;
        ELSIF x =- 6096 THEN
            sigmoid_f := 99;
        ELSIF x =- 6095 THEN
            sigmoid_f := 99;
        ELSIF x =- 6094 THEN
            sigmoid_f := 99;
        ELSIF x =- 6093 THEN
            sigmoid_f := 99;
        ELSIF x =- 6092 THEN
            sigmoid_f := 99;
        ELSIF x =- 6091 THEN
            sigmoid_f := 99;
        ELSIF x =- 6090 THEN
            sigmoid_f := 99;
        ELSIF x =- 6089 THEN
            sigmoid_f := 99;
        ELSIF x =- 6088 THEN
            sigmoid_f := 99;
        ELSIF x =- 6087 THEN
            sigmoid_f := 99;
        ELSIF x =- 6086 THEN
            sigmoid_f := 99;
        ELSIF x =- 6085 THEN
            sigmoid_f := 99;
        ELSIF x =- 6084 THEN
            sigmoid_f := 99;
        ELSIF x =- 6083 THEN
            sigmoid_f := 100;
        ELSIF x =- 6082 THEN
            sigmoid_f := 100;
        ELSIF x =- 6081 THEN
            sigmoid_f := 100;
        ELSIF x =- 6080 THEN
            sigmoid_f := 100;
        ELSIF x =- 6079 THEN
            sigmoid_f := 100;
        ELSIF x =- 6078 THEN
            sigmoid_f := 100;
        ELSIF x =- 6077 THEN
            sigmoid_f := 100;
        ELSIF x =- 6076 THEN
            sigmoid_f := 100;
        ELSIF x =- 6075 THEN
            sigmoid_f := 100;
        ELSIF x =- 6074 THEN
            sigmoid_f := 100;
        ELSIF x =- 6073 THEN
            sigmoid_f := 100;
        ELSIF x =- 6072 THEN
            sigmoid_f := 100;
        ELSIF x =- 6071 THEN
            sigmoid_f := 100;
        ELSIF x =- 6070 THEN
            sigmoid_f := 100;
        ELSIF x =- 6069 THEN
            sigmoid_f := 100;
        ELSIF x =- 6068 THEN
            sigmoid_f := 100;
        ELSIF x =- 6067 THEN
            sigmoid_f := 100;
        ELSIF x =- 6066 THEN
            sigmoid_f := 100;
        ELSIF x =- 6065 THEN
            sigmoid_f := 100;
        ELSIF x =- 6064 THEN
            sigmoid_f := 100;
        ELSIF x =- 6063 THEN
            sigmoid_f := 101;
        ELSIF x =- 6062 THEN
            sigmoid_f := 101;
        ELSIF x =- 6061 THEN
            sigmoid_f := 101;
        ELSIF x =- 6060 THEN
            sigmoid_f := 101;
        ELSIF x =- 6059 THEN
            sigmoid_f := 101;
        ELSIF x =- 6058 THEN
            sigmoid_f := 101;
        ELSIF x =- 6057 THEN
            sigmoid_f := 101;
        ELSIF x =- 6056 THEN
            sigmoid_f := 101;
        ELSIF x =- 6055 THEN
            sigmoid_f := 101;
        ELSIF x =- 6054 THEN
            sigmoid_f := 101;
        ELSIF x =- 6053 THEN
            sigmoid_f := 101;
        ELSIF x =- 6052 THEN
            sigmoid_f := 101;
        ELSIF x =- 6051 THEN
            sigmoid_f := 101;
        ELSIF x =- 6050 THEN
            sigmoid_f := 101;
        ELSIF x =- 6049 THEN
            sigmoid_f := 101;
        ELSIF x =- 6048 THEN
            sigmoid_f := 101;
        ELSIF x =- 6047 THEN
            sigmoid_f := 101;
        ELSIF x =- 6046 THEN
            sigmoid_f := 101;
        ELSIF x =- 6045 THEN
            sigmoid_f := 101;
        ELSIF x =- 6044 THEN
            sigmoid_f := 101;
        ELSIF x =- 6043 THEN
            sigmoid_f := 102;
        ELSIF x =- 6042 THEN
            sigmoid_f := 102;
        ELSIF x =- 6041 THEN
            sigmoid_f := 102;
        ELSIF x =- 6040 THEN
            sigmoid_f := 102;
        ELSIF x =- 6039 THEN
            sigmoid_f := 102;
        ELSIF x =- 6038 THEN
            sigmoid_f := 102;
        ELSIF x =- 6037 THEN
            sigmoid_f := 102;
        ELSIF x =- 6036 THEN
            sigmoid_f := 102;
        ELSIF x =- 6035 THEN
            sigmoid_f := 102;
        ELSIF x =- 6034 THEN
            sigmoid_f := 102;
        ELSIF x =- 6033 THEN
            sigmoid_f := 102;
        ELSIF x =- 6032 THEN
            sigmoid_f := 102;
        ELSIF x =- 6031 THEN
            sigmoid_f := 102;
        ELSIF x =- 6030 THEN
            sigmoid_f := 102;
        ELSIF x =- 6029 THEN
            sigmoid_f := 102;
        ELSIF x =- 6028 THEN
            sigmoid_f := 102;
        ELSIF x =- 6027 THEN
            sigmoid_f := 102;
        ELSIF x =- 6026 THEN
            sigmoid_f := 102;
        ELSIF x =- 6025 THEN
            sigmoid_f := 102;
        ELSIF x =- 6024 THEN
            sigmoid_f := 102;
        ELSIF x =- 6023 THEN
            sigmoid_f := 103;
        ELSIF x =- 6022 THEN
            sigmoid_f := 103;
        ELSIF x =- 6021 THEN
            sigmoid_f := 103;
        ELSIF x =- 6020 THEN
            sigmoid_f := 103;
        ELSIF x =- 6019 THEN
            sigmoid_f := 103;
        ELSIF x =- 6018 THEN
            sigmoid_f := 103;
        ELSIF x =- 6017 THEN
            sigmoid_f := 103;
        ELSIF x =- 6016 THEN
            sigmoid_f := 103;
        ELSIF x =- 6015 THEN
            sigmoid_f := 103;
        ELSIF x =- 6014 THEN
            sigmoid_f := 103;
        ELSIF x =- 6013 THEN
            sigmoid_f := 103;
        ELSIF x =- 6012 THEN
            sigmoid_f := 103;
        ELSIF x =- 6011 THEN
            sigmoid_f := 103;
        ELSIF x =- 6010 THEN
            sigmoid_f := 103;
        ELSIF x =- 6009 THEN
            sigmoid_f := 103;
        ELSIF x =- 6008 THEN
            sigmoid_f := 103;
        ELSIF x =- 6007 THEN
            sigmoid_f := 103;
        ELSIF x =- 6006 THEN
            sigmoid_f := 103;
        ELSIF x =- 6005 THEN
            sigmoid_f := 103;
        ELSIF x =- 6004 THEN
            sigmoid_f := 103;
        ELSIF x =- 6003 THEN
            sigmoid_f := 104;
        ELSIF x =- 6002 THEN
            sigmoid_f := 104;
        ELSIF x =- 6001 THEN
            sigmoid_f := 104;
        ELSIF x =- 6000 THEN
            sigmoid_f := 104;
        ELSIF x =- 5999 THEN
            sigmoid_f := 104;
        ELSIF x =- 5998 THEN
            sigmoid_f := 104;
        ELSIF x =- 5997 THEN
            sigmoid_f := 104;
        ELSIF x =- 5996 THEN
            sigmoid_f := 104;
        ELSIF x =- 5995 THEN
            sigmoid_f := 104;
        ELSIF x =- 5994 THEN
            sigmoid_f := 104;
        ELSIF x =- 5993 THEN
            sigmoid_f := 104;
        ELSIF x =- 5992 THEN
            sigmoid_f := 104;
        ELSIF x =- 5991 THEN
            sigmoid_f := 104;
        ELSIF x =- 5990 THEN
            sigmoid_f := 104;
        ELSIF x =- 5989 THEN
            sigmoid_f := 104;
        ELSIF x =- 5988 THEN
            sigmoid_f := 104;
        ELSIF x =- 5987 THEN
            sigmoid_f := 104;
        ELSIF x =- 5986 THEN
            sigmoid_f := 104;
        ELSIF x =- 5985 THEN
            sigmoid_f := 104;
        ELSIF x =- 5984 THEN
            sigmoid_f := 104;
        ELSIF x =- 5983 THEN
            sigmoid_f := 105;
        ELSIF x =- 5982 THEN
            sigmoid_f := 105;
        ELSIF x =- 5981 THEN
            sigmoid_f := 105;
        ELSIF x =- 5980 THEN
            sigmoid_f := 105;
        ELSIF x =- 5979 THEN
            sigmoid_f := 105;
        ELSIF x =- 5978 THEN
            sigmoid_f := 105;
        ELSIF x =- 5977 THEN
            sigmoid_f := 105;
        ELSIF x =- 5976 THEN
            sigmoid_f := 105;
        ELSIF x =- 5975 THEN
            sigmoid_f := 105;
        ELSIF x =- 5974 THEN
            sigmoid_f := 105;
        ELSIF x =- 5973 THEN
            sigmoid_f := 105;
        ELSIF x =- 5972 THEN
            sigmoid_f := 105;
        ELSIF x =- 5971 THEN
            sigmoid_f := 105;
        ELSIF x =- 5970 THEN
            sigmoid_f := 105;
        ELSIF x =- 5969 THEN
            sigmoid_f := 105;
        ELSIF x =- 5968 THEN
            sigmoid_f := 105;
        ELSIF x =- 5967 THEN
            sigmoid_f := 105;
        ELSIF x =- 5966 THEN
            sigmoid_f := 105;
        ELSIF x =- 5965 THEN
            sigmoid_f := 105;
        ELSIF x =- 5964 THEN
            sigmoid_f := 105;
        ELSIF x =- 5963 THEN
            sigmoid_f := 106;
        ELSIF x =- 5962 THEN
            sigmoid_f := 106;
        ELSIF x =- 5961 THEN
            sigmoid_f := 106;
        ELSIF x =- 5960 THEN
            sigmoid_f := 106;
        ELSIF x =- 5959 THEN
            sigmoid_f := 106;
        ELSIF x =- 5958 THEN
            sigmoid_f := 106;
        ELSIF x =- 5957 THEN
            sigmoid_f := 106;
        ELSIF x =- 5956 THEN
            sigmoid_f := 106;
        ELSIF x =- 5955 THEN
            sigmoid_f := 106;
        ELSIF x =- 5954 THEN
            sigmoid_f := 106;
        ELSIF x =- 5953 THEN
            sigmoid_f := 106;
        ELSIF x =- 5952 THEN
            sigmoid_f := 106;
        ELSIF x =- 5951 THEN
            sigmoid_f := 106;
        ELSIF x =- 5950 THEN
            sigmoid_f := 106;
        ELSIF x =- 5949 THEN
            sigmoid_f := 106;
        ELSIF x =- 5948 THEN
            sigmoid_f := 106;
        ELSIF x =- 5947 THEN
            sigmoid_f := 106;
        ELSIF x =- 5946 THEN
            sigmoid_f := 106;
        ELSIF x =- 5945 THEN
            sigmoid_f := 106;
        ELSIF x =- 5944 THEN
            sigmoid_f := 106;
        ELSIF x =- 5943 THEN
            sigmoid_f := 107;
        ELSIF x =- 5942 THEN
            sigmoid_f := 107;
        ELSIF x =- 5941 THEN
            sigmoid_f := 107;
        ELSIF x =- 5940 THEN
            sigmoid_f := 107;
        ELSIF x =- 5939 THEN
            sigmoid_f := 107;
        ELSIF x =- 5938 THEN
            sigmoid_f := 107;
        ELSIF x =- 5937 THEN
            sigmoid_f := 107;
        ELSIF x =- 5936 THEN
            sigmoid_f := 107;
        ELSIF x =- 5935 THEN
            sigmoid_f := 107;
        ELSIF x =- 5934 THEN
            sigmoid_f := 107;
        ELSIF x =- 5933 THEN
            sigmoid_f := 107;
        ELSIF x =- 5932 THEN
            sigmoid_f := 107;
        ELSIF x =- 5931 THEN
            sigmoid_f := 107;
        ELSIF x =- 5930 THEN
            sigmoid_f := 107;
        ELSIF x =- 5929 THEN
            sigmoid_f := 107;
        ELSIF x =- 5928 THEN
            sigmoid_f := 107;
        ELSIF x =- 5927 THEN
            sigmoid_f := 107;
        ELSIF x =- 5926 THEN
            sigmoid_f := 107;
        ELSIF x =- 5925 THEN
            sigmoid_f := 107;
        ELSIF x =- 5924 THEN
            sigmoid_f := 107;
        ELSIF x =- 5923 THEN
            sigmoid_f := 108;
        ELSIF x =- 5922 THEN
            sigmoid_f := 108;
        ELSIF x =- 5921 THEN
            sigmoid_f := 108;
        ELSIF x =- 5920 THEN
            sigmoid_f := 108;
        ELSIF x =- 5919 THEN
            sigmoid_f := 108;
        ELSIF x =- 5918 THEN
            sigmoid_f := 108;
        ELSIF x =- 5917 THEN
            sigmoid_f := 108;
        ELSIF x =- 5916 THEN
            sigmoid_f := 108;
        ELSIF x =- 5915 THEN
            sigmoid_f := 108;
        ELSIF x =- 5914 THEN
            sigmoid_f := 108;
        ELSIF x =- 5913 THEN
            sigmoid_f := 108;
        ELSIF x =- 5912 THEN
            sigmoid_f := 108;
        ELSIF x =- 5911 THEN
            sigmoid_f := 108;
        ELSIF x =- 5910 THEN
            sigmoid_f := 108;
        ELSIF x =- 5909 THEN
            sigmoid_f := 108;
        ELSIF x =- 5908 THEN
            sigmoid_f := 108;
        ELSIF x =- 5907 THEN
            sigmoid_f := 108;
        ELSIF x =- 5906 THEN
            sigmoid_f := 108;
        ELSIF x =- 5905 THEN
            sigmoid_f := 108;
        ELSIF x =- 5904 THEN
            sigmoid_f := 108;
        ELSIF x =- 5903 THEN
            sigmoid_f := 109;
        ELSIF x =- 5902 THEN
            sigmoid_f := 109;
        ELSIF x =- 5901 THEN
            sigmoid_f := 109;
        ELSIF x =- 5900 THEN
            sigmoid_f := 109;
        ELSIF x =- 5899 THEN
            sigmoid_f := 109;
        ELSIF x =- 5898 THEN
            sigmoid_f := 109;
        ELSIF x =- 5897 THEN
            sigmoid_f := 109;
        ELSIF x =- 5896 THEN
            sigmoid_f := 109;
        ELSIF x =- 5895 THEN
            sigmoid_f := 109;
        ELSIF x =- 5894 THEN
            sigmoid_f := 109;
        ELSIF x =- 5893 THEN
            sigmoid_f := 109;
        ELSIF x =- 5892 THEN
            sigmoid_f := 109;
        ELSIF x =- 5891 THEN
            sigmoid_f := 109;
        ELSIF x =- 5890 THEN
            sigmoid_f := 109;
        ELSIF x =- 5889 THEN
            sigmoid_f := 109;
        ELSIF x =- 5888 THEN
            sigmoid_f := 109;
        ELSIF x =- 5887 THEN
            sigmoid_f := 109;
        ELSIF x =- 5886 THEN
            sigmoid_f := 109;
        ELSIF x =- 5885 THEN
            sigmoid_f := 109;
        ELSIF x =- 5884 THEN
            sigmoid_f := 109;
        ELSIF x =- 5883 THEN
            sigmoid_f := 109;
        ELSIF x =- 5882 THEN
            sigmoid_f := 110;
        ELSIF x =- 5881 THEN
            sigmoid_f := 110;
        ELSIF x =- 5880 THEN
            sigmoid_f := 110;
        ELSIF x =- 5879 THEN
            sigmoid_f := 110;
        ELSIF x =- 5878 THEN
            sigmoid_f := 110;
        ELSIF x =- 5877 THEN
            sigmoid_f := 110;
        ELSIF x =- 5876 THEN
            sigmoid_f := 110;
        ELSIF x =- 5875 THEN
            sigmoid_f := 110;
        ELSIF x =- 5874 THEN
            sigmoid_f := 110;
        ELSIF x =- 5873 THEN
            sigmoid_f := 110;
        ELSIF x =- 5872 THEN
            sigmoid_f := 110;
        ELSIF x =- 5871 THEN
            sigmoid_f := 110;
        ELSIF x =- 5870 THEN
            sigmoid_f := 110;
        ELSIF x =- 5869 THEN
            sigmoid_f := 110;
        ELSIF x =- 5868 THEN
            sigmoid_f := 110;
        ELSIF x =- 5867 THEN
            sigmoid_f := 110;
        ELSIF x =- 5866 THEN
            sigmoid_f := 110;
        ELSIF x =- 5865 THEN
            sigmoid_f := 110;
        ELSIF x =- 5864 THEN
            sigmoid_f := 110;
        ELSIF x =- 5863 THEN
            sigmoid_f := 110;
        ELSIF x =- 5862 THEN
            sigmoid_f := 111;
        ELSIF x =- 5861 THEN
            sigmoid_f := 111;
        ELSIF x =- 5860 THEN
            sigmoid_f := 111;
        ELSIF x =- 5859 THEN
            sigmoid_f := 111;
        ELSIF x =- 5858 THEN
            sigmoid_f := 111;
        ELSIF x =- 5857 THEN
            sigmoid_f := 111;
        ELSIF x =- 5856 THEN
            sigmoid_f := 111;
        ELSIF x =- 5855 THEN
            sigmoid_f := 111;
        ELSIF x =- 5854 THEN
            sigmoid_f := 111;
        ELSIF x =- 5853 THEN
            sigmoid_f := 111;
        ELSIF x =- 5852 THEN
            sigmoid_f := 111;
        ELSIF x =- 5851 THEN
            sigmoid_f := 111;
        ELSIF x =- 5850 THEN
            sigmoid_f := 111;
        ELSIF x =- 5849 THEN
            sigmoid_f := 111;
        ELSIF x =- 5848 THEN
            sigmoid_f := 111;
        ELSIF x =- 5847 THEN
            sigmoid_f := 111;
        ELSIF x =- 5846 THEN
            sigmoid_f := 111;
        ELSIF x =- 5845 THEN
            sigmoid_f := 111;
        ELSIF x =- 5844 THEN
            sigmoid_f := 111;
        ELSIF x =- 5843 THEN
            sigmoid_f := 111;
        ELSIF x =- 5842 THEN
            sigmoid_f := 112;
        ELSIF x =- 5841 THEN
            sigmoid_f := 112;
        ELSIF x =- 5840 THEN
            sigmoid_f := 112;
        ELSIF x =- 5839 THEN
            sigmoid_f := 112;
        ELSIF x =- 5838 THEN
            sigmoid_f := 112;
        ELSIF x =- 5837 THEN
            sigmoid_f := 112;
        ELSIF x =- 5836 THEN
            sigmoid_f := 112;
        ELSIF x =- 5835 THEN
            sigmoid_f := 112;
        ELSIF x =- 5834 THEN
            sigmoid_f := 112;
        ELSIF x =- 5833 THEN
            sigmoid_f := 112;
        ELSIF x =- 5832 THEN
            sigmoid_f := 112;
        ELSIF x =- 5831 THEN
            sigmoid_f := 112;
        ELSIF x =- 5830 THEN
            sigmoid_f := 112;
        ELSIF x =- 5829 THEN
            sigmoid_f := 112;
        ELSIF x =- 5828 THEN
            sigmoid_f := 112;
        ELSIF x =- 5827 THEN
            sigmoid_f := 112;
        ELSIF x =- 5826 THEN
            sigmoid_f := 112;
        ELSIF x =- 5825 THEN
            sigmoid_f := 112;
        ELSIF x =- 5824 THEN
            sigmoid_f := 112;
        ELSIF x =- 5823 THEN
            sigmoid_f := 112;
        ELSIF x =- 5822 THEN
            sigmoid_f := 113;
        ELSIF x =- 5821 THEN
            sigmoid_f := 113;
        ELSIF x =- 5820 THEN
            sigmoid_f := 113;
        ELSIF x =- 5819 THEN
            sigmoid_f := 113;
        ELSIF x =- 5818 THEN
            sigmoid_f := 113;
        ELSIF x =- 5817 THEN
            sigmoid_f := 113;
        ELSIF x =- 5816 THEN
            sigmoid_f := 113;
        ELSIF x =- 5815 THEN
            sigmoid_f := 113;
        ELSIF x =- 5814 THEN
            sigmoid_f := 113;
        ELSIF x =- 5813 THEN
            sigmoid_f := 113;
        ELSIF x =- 5812 THEN
            sigmoid_f := 113;
        ELSIF x =- 5811 THEN
            sigmoid_f := 113;
        ELSIF x =- 5810 THEN
            sigmoid_f := 113;
        ELSIF x =- 5809 THEN
            sigmoid_f := 113;
        ELSIF x =- 5808 THEN
            sigmoid_f := 113;
        ELSIF x =- 5807 THEN
            sigmoid_f := 113;
        ELSIF x =- 5806 THEN
            sigmoid_f := 113;
        ELSIF x =- 5805 THEN
            sigmoid_f := 113;
        ELSIF x =- 5804 THEN
            sigmoid_f := 113;
        ELSIF x =- 5803 THEN
            sigmoid_f := 113;
        ELSIF x =- 5802 THEN
            sigmoid_f := 114;
        ELSIF x =- 5801 THEN
            sigmoid_f := 114;
        ELSIF x =- 5800 THEN
            sigmoid_f := 114;
        ELSIF x =- 5799 THEN
            sigmoid_f := 114;
        ELSIF x =- 5798 THEN
            sigmoid_f := 114;
        ELSIF x =- 5797 THEN
            sigmoid_f := 114;
        ELSIF x =- 5796 THEN
            sigmoid_f := 114;
        ELSIF x =- 5795 THEN
            sigmoid_f := 114;
        ELSIF x =- 5794 THEN
            sigmoid_f := 114;
        ELSIF x =- 5793 THEN
            sigmoid_f := 114;
        ELSIF x =- 5792 THEN
            sigmoid_f := 114;
        ELSIF x =- 5791 THEN
            sigmoid_f := 114;
        ELSIF x =- 5790 THEN
            sigmoid_f := 114;
        ELSIF x =- 5789 THEN
            sigmoid_f := 114;
        ELSIF x =- 5788 THEN
            sigmoid_f := 114;
        ELSIF x =- 5787 THEN
            sigmoid_f := 114;
        ELSIF x =- 5786 THEN
            sigmoid_f := 114;
        ELSIF x =- 5785 THEN
            sigmoid_f := 114;
        ELSIF x =- 5784 THEN
            sigmoid_f := 114;
        ELSIF x =- 5783 THEN
            sigmoid_f := 114;
        ELSIF x =- 5782 THEN
            sigmoid_f := 115;
        ELSIF x =- 5781 THEN
            sigmoid_f := 115;
        ELSIF x =- 5780 THEN
            sigmoid_f := 115;
        ELSIF x =- 5779 THEN
            sigmoid_f := 115;
        ELSIF x =- 5778 THEN
            sigmoid_f := 115;
        ELSIF x =- 5777 THEN
            sigmoid_f := 115;
        ELSIF x =- 5776 THEN
            sigmoid_f := 115;
        ELSIF x =- 5775 THEN
            sigmoid_f := 115;
        ELSIF x =- 5774 THEN
            sigmoid_f := 115;
        ELSIF x =- 5773 THEN
            sigmoid_f := 115;
        ELSIF x =- 5772 THEN
            sigmoid_f := 115;
        ELSIF x =- 5771 THEN
            sigmoid_f := 115;
        ELSIF x =- 5770 THEN
            sigmoid_f := 115;
        ELSIF x =- 5769 THEN
            sigmoid_f := 115;
        ELSIF x =- 5768 THEN
            sigmoid_f := 115;
        ELSIF x =- 5767 THEN
            sigmoid_f := 115;
        ELSIF x =- 5766 THEN
            sigmoid_f := 115;
        ELSIF x =- 5765 THEN
            sigmoid_f := 115;
        ELSIF x =- 5764 THEN
            sigmoid_f := 115;
        ELSIF x =- 5763 THEN
            sigmoid_f := 115;
        ELSIF x =- 5762 THEN
            sigmoid_f := 116;
        ELSIF x =- 5761 THEN
            sigmoid_f := 116;
        ELSIF x =- 5760 THEN
            sigmoid_f := 116;
        ELSIF x =- 5759 THEN
            sigmoid_f := 116;
        ELSIF x =- 5758 THEN
            sigmoid_f := 116;
        ELSIF x =- 5757 THEN
            sigmoid_f := 116;
        ELSIF x =- 5756 THEN
            sigmoid_f := 116;
        ELSIF x =- 5755 THEN
            sigmoid_f := 116;
        ELSIF x =- 5754 THEN
            sigmoid_f := 116;
        ELSIF x =- 5753 THEN
            sigmoid_f := 116;
        ELSIF x =- 5752 THEN
            sigmoid_f := 116;
        ELSIF x =- 5751 THEN
            sigmoid_f := 116;
        ELSIF x =- 5750 THEN
            sigmoid_f := 116;
        ELSIF x =- 5749 THEN
            sigmoid_f := 116;
        ELSIF x =- 5748 THEN
            sigmoid_f := 116;
        ELSIF x =- 5747 THEN
            sigmoid_f := 116;
        ELSIF x =- 5746 THEN
            sigmoid_f := 116;
        ELSIF x =- 5745 THEN
            sigmoid_f := 116;
        ELSIF x =- 5744 THEN
            sigmoid_f := 116;
        ELSIF x =- 5743 THEN
            sigmoid_f := 116;
        ELSIF x =- 5742 THEN
            sigmoid_f := 117;
        ELSIF x =- 5741 THEN
            sigmoid_f := 117;
        ELSIF x =- 5740 THEN
            sigmoid_f := 117;
        ELSIF x =- 5739 THEN
            sigmoid_f := 117;
        ELSIF x =- 5738 THEN
            sigmoid_f := 117;
        ELSIF x =- 5737 THEN
            sigmoid_f := 117;
        ELSIF x =- 5736 THEN
            sigmoid_f := 117;
        ELSIF x =- 5735 THEN
            sigmoid_f := 117;
        ELSIF x =- 5734 THEN
            sigmoid_f := 117;
        ELSIF x =- 5733 THEN
            sigmoid_f := 117;
        ELSIF x =- 5732 THEN
            sigmoid_f := 117;
        ELSIF x =- 5731 THEN
            sigmoid_f := 117;
        ELSIF x =- 5730 THEN
            sigmoid_f := 117;
        ELSIF x =- 5729 THEN
            sigmoid_f := 117;
        ELSIF x =- 5728 THEN
            sigmoid_f := 117;
        ELSIF x =- 5727 THEN
            sigmoid_f := 117;
        ELSIF x =- 5726 THEN
            sigmoid_f := 117;
        ELSIF x =- 5725 THEN
            sigmoid_f := 117;
        ELSIF x =- 5724 THEN
            sigmoid_f := 117;
        ELSIF x =- 5723 THEN
            sigmoid_f := 117;
        ELSIF x =- 5722 THEN
            sigmoid_f := 118;
        ELSIF x =- 5721 THEN
            sigmoid_f := 118;
        ELSIF x =- 5720 THEN
            sigmoid_f := 118;
        ELSIF x =- 5719 THEN
            sigmoid_f := 118;
        ELSIF x =- 5718 THEN
            sigmoid_f := 118;
        ELSIF x =- 5717 THEN
            sigmoid_f := 118;
        ELSIF x =- 5716 THEN
            sigmoid_f := 118;
        ELSIF x =- 5715 THEN
            sigmoid_f := 118;
        ELSIF x =- 5714 THEN
            sigmoid_f := 118;
        ELSIF x =- 5713 THEN
            sigmoid_f := 118;
        ELSIF x =- 5712 THEN
            sigmoid_f := 118;
        ELSIF x =- 5711 THEN
            sigmoid_f := 118;
        ELSIF x =- 5710 THEN
            sigmoid_f := 118;
        ELSIF x =- 5709 THEN
            sigmoid_f := 118;
        ELSIF x =- 5708 THEN
            sigmoid_f := 118;
        ELSIF x =- 5707 THEN
            sigmoid_f := 118;
        ELSIF x =- 5706 THEN
            sigmoid_f := 118;
        ELSIF x =- 5705 THEN
            sigmoid_f := 118;
        ELSIF x =- 5704 THEN
            sigmoid_f := 118;
        ELSIF x =- 5703 THEN
            sigmoid_f := 118;
        ELSIF x =- 5702 THEN
            sigmoid_f := 119;
        ELSIF x =- 5701 THEN
            sigmoid_f := 119;
        ELSIF x =- 5700 THEN
            sigmoid_f := 119;
        ELSIF x =- 5699 THEN
            sigmoid_f := 119;
        ELSIF x =- 5698 THEN
            sigmoid_f := 119;
        ELSIF x =- 5697 THEN
            sigmoid_f := 119;
        ELSIF x =- 5696 THEN
            sigmoid_f := 119;
        ELSIF x =- 5695 THEN
            sigmoid_f := 119;
        ELSIF x =- 5694 THEN
            sigmoid_f := 119;
        ELSIF x =- 5693 THEN
            sigmoid_f := 119;
        ELSIF x =- 5692 THEN
            sigmoid_f := 119;
        ELSIF x =- 5691 THEN
            sigmoid_f := 119;
        ELSIF x =- 5690 THEN
            sigmoid_f := 119;
        ELSIF x =- 5689 THEN
            sigmoid_f := 119;
        ELSIF x =- 5688 THEN
            sigmoid_f := 119;
        ELSIF x =- 5687 THEN
            sigmoid_f := 119;
        ELSIF x =- 5686 THEN
            sigmoid_f := 119;
        ELSIF x =- 5685 THEN
            sigmoid_f := 119;
        ELSIF x =- 5684 THEN
            sigmoid_f := 119;
        ELSIF x =- 5683 THEN
            sigmoid_f := 119;
        ELSIF x =- 5682 THEN
            sigmoid_f := 120;
        ELSIF x =- 5681 THEN
            sigmoid_f := 120;
        ELSIF x =- 5680 THEN
            sigmoid_f := 120;
        ELSIF x =- 5679 THEN
            sigmoid_f := 120;
        ELSIF x =- 5678 THEN
            sigmoid_f := 120;
        ELSIF x =- 5677 THEN
            sigmoid_f := 120;
        ELSIF x =- 5676 THEN
            sigmoid_f := 120;
        ELSIF x =- 5675 THEN
            sigmoid_f := 120;
        ELSIF x =- 5674 THEN
            sigmoid_f := 120;
        ELSIF x =- 5673 THEN
            sigmoid_f := 120;
        ELSIF x =- 5672 THEN
            sigmoid_f := 120;
        ELSIF x =- 5671 THEN
            sigmoid_f := 120;
        ELSIF x =- 5670 THEN
            sigmoid_f := 120;
        ELSIF x =- 5669 THEN
            sigmoid_f := 120;
        ELSIF x =- 5668 THEN
            sigmoid_f := 120;
        ELSIF x =- 5667 THEN
            sigmoid_f := 120;
        ELSIF x =- 5666 THEN
            sigmoid_f := 120;
        ELSIF x =- 5665 THEN
            sigmoid_f := 120;
        ELSIF x =- 5664 THEN
            sigmoid_f := 120;
        ELSIF x =- 5663 THEN
            sigmoid_f := 120;
        ELSIF x =- 5662 THEN
            sigmoid_f := 121;
        ELSIF x =- 5661 THEN
            sigmoid_f := 121;
        ELSIF x =- 5660 THEN
            sigmoid_f := 121;
        ELSIF x =- 5659 THEN
            sigmoid_f := 121;
        ELSIF x =- 5658 THEN
            sigmoid_f := 121;
        ELSIF x =- 5657 THEN
            sigmoid_f := 121;
        ELSIF x =- 5656 THEN
            sigmoid_f := 121;
        ELSIF x =- 5655 THEN
            sigmoid_f := 121;
        ELSIF x =- 5654 THEN
            sigmoid_f := 121;
        ELSIF x =- 5653 THEN
            sigmoid_f := 121;
        ELSIF x =- 5652 THEN
            sigmoid_f := 121;
        ELSIF x =- 5651 THEN
            sigmoid_f := 121;
        ELSIF x =- 5650 THEN
            sigmoid_f := 121;
        ELSIF x =- 5649 THEN
            sigmoid_f := 121;
        ELSIF x =- 5648 THEN
            sigmoid_f := 121;
        ELSIF x =- 5647 THEN
            sigmoid_f := 121;
        ELSIF x =- 5646 THEN
            sigmoid_f := 121;
        ELSIF x =- 5645 THEN
            sigmoid_f := 121;
        ELSIF x =- 5644 THEN
            sigmoid_f := 121;
        ELSIF x =- 5643 THEN
            sigmoid_f := 121;
        ELSIF x =- 5642 THEN
            sigmoid_f := 122;
        ELSIF x =- 5641 THEN
            sigmoid_f := 122;
        ELSIF x =- 5640 THEN
            sigmoid_f := 122;
        ELSIF x =- 5639 THEN
            sigmoid_f := 122;
        ELSIF x =- 5638 THEN
            sigmoid_f := 122;
        ELSIF x =- 5637 THEN
            sigmoid_f := 122;
        ELSIF x =- 5636 THEN
            sigmoid_f := 122;
        ELSIF x =- 5635 THEN
            sigmoid_f := 122;
        ELSIF x =- 5634 THEN
            sigmoid_f := 122;
        ELSIF x =- 5633 THEN
            sigmoid_f := 122;
        ELSIF x =- 5632 THEN
            sigmoid_f := 122;
        ELSIF x =- 5631 THEN
            sigmoid_f := 122;
        ELSIF x =- 5630 THEN
            sigmoid_f := 122;
        ELSIF x =- 5629 THEN
            sigmoid_f := 122;
        ELSIF x =- 5628 THEN
            sigmoid_f := 122;
        ELSIF x =- 5627 THEN
            sigmoid_f := 123;
        ELSIF x =- 5626 THEN
            sigmoid_f := 123;
        ELSIF x =- 5625 THEN
            sigmoid_f := 123;
        ELSIF x =- 5624 THEN
            sigmoid_f := 123;
        ELSIF x =- 5623 THEN
            sigmoid_f := 123;
        ELSIF x =- 5622 THEN
            sigmoid_f := 123;
        ELSIF x =- 5621 THEN
            sigmoid_f := 123;
        ELSIF x =- 5620 THEN
            sigmoid_f := 123;
        ELSIF x =- 5619 THEN
            sigmoid_f := 123;
        ELSIF x =- 5618 THEN
            sigmoid_f := 123;
        ELSIF x =- 5617 THEN
            sigmoid_f := 123;
        ELSIF x =- 5616 THEN
            sigmoid_f := 123;
        ELSIF x =- 5615 THEN
            sigmoid_f := 123;
        ELSIF x =- 5614 THEN
            sigmoid_f := 123;
        ELSIF x =- 5613 THEN
            sigmoid_f := 123;
        ELSIF x =- 5612 THEN
            sigmoid_f := 123;
        ELSIF x =- 5611 THEN
            sigmoid_f := 124;
        ELSIF x =- 5610 THEN
            sigmoid_f := 124;
        ELSIF x =- 5609 THEN
            sigmoid_f := 124;
        ELSIF x =- 5608 THEN
            sigmoid_f := 124;
        ELSIF x =- 5607 THEN
            sigmoid_f := 124;
        ELSIF x =- 5606 THEN
            sigmoid_f := 124;
        ELSIF x =- 5605 THEN
            sigmoid_f := 124;
        ELSIF x =- 5604 THEN
            sigmoid_f := 124;
        ELSIF x =- 5603 THEN
            sigmoid_f := 124;
        ELSIF x =- 5602 THEN
            sigmoid_f := 124;
        ELSIF x =- 5601 THEN
            sigmoid_f := 124;
        ELSIF x =- 5600 THEN
            sigmoid_f := 124;
        ELSIF x =- 5599 THEN
            sigmoid_f := 124;
        ELSIF x =- 5598 THEN
            sigmoid_f := 124;
        ELSIF x =- 5597 THEN
            sigmoid_f := 124;
        ELSIF x =- 5596 THEN
            sigmoid_f := 124;
        ELSIF x =- 5595 THEN
            sigmoid_f := 125;
        ELSIF x =- 5594 THEN
            sigmoid_f := 125;
        ELSIF x =- 5593 THEN
            sigmoid_f := 125;
        ELSIF x =- 5592 THEN
            sigmoid_f := 125;
        ELSIF x =- 5591 THEN
            sigmoid_f := 125;
        ELSIF x =- 5590 THEN
            sigmoid_f := 125;
        ELSIF x =- 5589 THEN
            sigmoid_f := 125;
        ELSIF x =- 5588 THEN
            sigmoid_f := 125;
        ELSIF x =- 5587 THEN
            sigmoid_f := 125;
        ELSIF x =- 5586 THEN
            sigmoid_f := 125;
        ELSIF x =- 5585 THEN
            sigmoid_f := 125;
        ELSIF x =- 5584 THEN
            sigmoid_f := 125;
        ELSIF x =- 5583 THEN
            sigmoid_f := 125;
        ELSIF x =- 5582 THEN
            sigmoid_f := 125;
        ELSIF x =- 5581 THEN
            sigmoid_f := 125;
        ELSIF x =- 5580 THEN
            sigmoid_f := 125;
        ELSIF x =- 5579 THEN
            sigmoid_f := 126;
        ELSIF x =- 5578 THEN
            sigmoid_f := 126;
        ELSIF x =- 5577 THEN
            sigmoid_f := 126;
        ELSIF x =- 5576 THEN
            sigmoid_f := 126;
        ELSIF x =- 5575 THEN
            sigmoid_f := 126;
        ELSIF x =- 5574 THEN
            sigmoid_f := 126;
        ELSIF x =- 5573 THEN
            sigmoid_f := 126;
        ELSIF x =- 5572 THEN
            sigmoid_f := 126;
        ELSIF x =- 5571 THEN
            sigmoid_f := 126;
        ELSIF x =- 5570 THEN
            sigmoid_f := 126;
        ELSIF x =- 5569 THEN
            sigmoid_f := 126;
        ELSIF x =- 5568 THEN
            sigmoid_f := 126;
        ELSIF x =- 5567 THEN
            sigmoid_f := 126;
        ELSIF x =- 5566 THEN
            sigmoid_f := 126;
        ELSIF x =- 5565 THEN
            sigmoid_f := 126;
        ELSIF x =- 5564 THEN
            sigmoid_f := 126;
        ELSIF x =- 5563 THEN
            sigmoid_f := 127;
        ELSIF x =- 5562 THEN
            sigmoid_f := 127;
        ELSIF x =- 5561 THEN
            sigmoid_f := 127;
        ELSIF x =- 5560 THEN
            sigmoid_f := 127;
        ELSIF x =- 5559 THEN
            sigmoid_f := 127;
        ELSIF x =- 5558 THEN
            sigmoid_f := 127;
        ELSIF x =- 5557 THEN
            sigmoid_f := 127;
        ELSIF x =- 5556 THEN
            sigmoid_f := 127;
        ELSIF x =- 5555 THEN
            sigmoid_f := 127;
        ELSIF x =- 5554 THEN
            sigmoid_f := 127;
        ELSIF x =- 5553 THEN
            sigmoid_f := 127;
        ELSIF x =- 5552 THEN
            sigmoid_f := 127;
        ELSIF x =- 5551 THEN
            sigmoid_f := 127;
        ELSIF x =- 5550 THEN
            sigmoid_f := 127;
        ELSIF x =- 5549 THEN
            sigmoid_f := 127;
        ELSIF x =- 5548 THEN
            sigmoid_f := 127;
        ELSIF x =- 5547 THEN
            sigmoid_f := 128;
        ELSIF x =- 5546 THEN
            sigmoid_f := 128;
        ELSIF x =- 5545 THEN
            sigmoid_f := 128;
        ELSIF x =- 5544 THEN
            sigmoid_f := 128;
        ELSIF x =- 5543 THEN
            sigmoid_f := 128;
        ELSIF x =- 5542 THEN
            sigmoid_f := 128;
        ELSIF x =- 5541 THEN
            sigmoid_f := 128;
        ELSIF x =- 5540 THEN
            sigmoid_f := 128;
        ELSIF x =- 5539 THEN
            sigmoid_f := 128;
        ELSIF x =- 5538 THEN
            sigmoid_f := 128;
        ELSIF x =- 5537 THEN
            sigmoid_f := 128;
        ELSIF x =- 5536 THEN
            sigmoid_f := 128;
        ELSIF x =- 5535 THEN
            sigmoid_f := 128;
        ELSIF x =- 5534 THEN
            sigmoid_f := 128;
        ELSIF x =- 5533 THEN
            sigmoid_f := 128;
        ELSIF x =- 5532 THEN
            sigmoid_f := 128;
        ELSIF x =- 5531 THEN
            sigmoid_f := 129;
        ELSIF x =- 5530 THEN
            sigmoid_f := 129;
        ELSIF x =- 5529 THEN
            sigmoid_f := 129;
        ELSIF x =- 5528 THEN
            sigmoid_f := 129;
        ELSIF x =- 5527 THEN
            sigmoid_f := 129;
        ELSIF x =- 5526 THEN
            sigmoid_f := 129;
        ELSIF x =- 5525 THEN
            sigmoid_f := 129;
        ELSIF x =- 5524 THEN
            sigmoid_f := 129;
        ELSIF x =- 5523 THEN
            sigmoid_f := 129;
        ELSIF x =- 5522 THEN
            sigmoid_f := 129;
        ELSIF x =- 5521 THEN
            sigmoid_f := 129;
        ELSIF x =- 5520 THEN
            sigmoid_f := 129;
        ELSIF x =- 5519 THEN
            sigmoid_f := 129;
        ELSIF x =- 5518 THEN
            sigmoid_f := 129;
        ELSIF x =- 5517 THEN
            sigmoid_f := 129;
        ELSIF x =- 5516 THEN
            sigmoid_f := 129;
        ELSIF x =- 5515 THEN
            sigmoid_f := 130;
        ELSIF x =- 5514 THEN
            sigmoid_f := 130;
        ELSIF x =- 5513 THEN
            sigmoid_f := 130;
        ELSIF x =- 5512 THEN
            sigmoid_f := 130;
        ELSIF x =- 5511 THEN
            sigmoid_f := 130;
        ELSIF x =- 5510 THEN
            sigmoid_f := 130;
        ELSIF x =- 5509 THEN
            sigmoid_f := 130;
        ELSIF x =- 5508 THEN
            sigmoid_f := 130;
        ELSIF x =- 5507 THEN
            sigmoid_f := 130;
        ELSIF x =- 5506 THEN
            sigmoid_f := 130;
        ELSIF x =- 5505 THEN
            sigmoid_f := 130;
        ELSIF x =- 5504 THEN
            sigmoid_f := 130;
        ELSIF x =- 5503 THEN
            sigmoid_f := 130;
        ELSIF x =- 5502 THEN
            sigmoid_f := 130;
        ELSIF x =- 5501 THEN
            sigmoid_f := 130;
        ELSIF x =- 5500 THEN
            sigmoid_f := 130;
        ELSIF x =- 5499 THEN
            sigmoid_f := 130;
        ELSIF x =- 5498 THEN
            sigmoid_f := 131;
        ELSIF x =- 5497 THEN
            sigmoid_f := 131;
        ELSIF x =- 5496 THEN
            sigmoid_f := 131;
        ELSIF x =- 5495 THEN
            sigmoid_f := 131;
        ELSIF x =- 5494 THEN
            sigmoid_f := 131;
        ELSIF x =- 5493 THEN
            sigmoid_f := 131;
        ELSIF x =- 5492 THEN
            sigmoid_f := 131;
        ELSIF x =- 5491 THEN
            sigmoid_f := 131;
        ELSIF x =- 5490 THEN
            sigmoid_f := 131;
        ELSIF x =- 5489 THEN
            sigmoid_f := 131;
        ELSIF x =- 5488 THEN
            sigmoid_f := 131;
        ELSIF x =- 5487 THEN
            sigmoid_f := 131;
        ELSIF x =- 5486 THEN
            sigmoid_f := 131;
        ELSIF x =- 5485 THEN
            sigmoid_f := 131;
        ELSIF x =- 5484 THEN
            sigmoid_f := 131;
        ELSIF x =- 5483 THEN
            sigmoid_f := 131;
        ELSIF x =- 5482 THEN
            sigmoid_f := 132;
        ELSIF x =- 5481 THEN
            sigmoid_f := 132;
        ELSIF x =- 5480 THEN
            sigmoid_f := 132;
        ELSIF x =- 5479 THEN
            sigmoid_f := 132;
        ELSIF x =- 5478 THEN
            sigmoid_f := 132;
        ELSIF x =- 5477 THEN
            sigmoid_f := 132;
        ELSIF x =- 5476 THEN
            sigmoid_f := 132;
        ELSIF x =- 5475 THEN
            sigmoid_f := 132;
        ELSIF x =- 5474 THEN
            sigmoid_f := 132;
        ELSIF x =- 5473 THEN
            sigmoid_f := 132;
        ELSIF x =- 5472 THEN
            sigmoid_f := 132;
        ELSIF x =- 5471 THEN
            sigmoid_f := 132;
        ELSIF x =- 5470 THEN
            sigmoid_f := 132;
        ELSIF x =- 5469 THEN
            sigmoid_f := 132;
        ELSIF x =- 5468 THEN
            sigmoid_f := 132;
        ELSIF x =- 5467 THEN
            sigmoid_f := 132;
        ELSIF x =- 5466 THEN
            sigmoid_f := 133;
        ELSIF x =- 5465 THEN
            sigmoid_f := 133;
        ELSIF x =- 5464 THEN
            sigmoid_f := 133;
        ELSIF x =- 5463 THEN
            sigmoid_f := 133;
        ELSIF x =- 5462 THEN
            sigmoid_f := 133;
        ELSIF x =- 5461 THEN
            sigmoid_f := 133;
        ELSIF x =- 5460 THEN
            sigmoid_f := 133;
        ELSIF x =- 5459 THEN
            sigmoid_f := 133;
        ELSIF x =- 5458 THEN
            sigmoid_f := 133;
        ELSIF x =- 5457 THEN
            sigmoid_f := 133;
        ELSIF x =- 5456 THEN
            sigmoid_f := 133;
        ELSIF x =- 5455 THEN
            sigmoid_f := 133;
        ELSIF x =- 5454 THEN
            sigmoid_f := 133;
        ELSIF x =- 5453 THEN
            sigmoid_f := 133;
        ELSIF x =- 5452 THEN
            sigmoid_f := 133;
        ELSIF x =- 5451 THEN
            sigmoid_f := 133;
        ELSIF x =- 5450 THEN
            sigmoid_f := 134;
        ELSIF x =- 5449 THEN
            sigmoid_f := 134;
        ELSIF x =- 5448 THEN
            sigmoid_f := 134;
        ELSIF x =- 5447 THEN
            sigmoid_f := 134;
        ELSIF x =- 5446 THEN
            sigmoid_f := 134;
        ELSIF x =- 5445 THEN
            sigmoid_f := 134;
        ELSIF x =- 5444 THEN
            sigmoid_f := 134;
        ELSIF x =- 5443 THEN
            sigmoid_f := 134;
        ELSIF x =- 5442 THEN
            sigmoid_f := 134;
        ELSIF x =- 5441 THEN
            sigmoid_f := 134;
        ELSIF x =- 5440 THEN
            sigmoid_f := 134;
        ELSIF x =- 5439 THEN
            sigmoid_f := 134;
        ELSIF x =- 5438 THEN
            sigmoid_f := 134;
        ELSIF x =- 5437 THEN
            sigmoid_f := 134;
        ELSIF x =- 5436 THEN
            sigmoid_f := 134;
        ELSIF x =- 5435 THEN
            sigmoid_f := 134;
        ELSIF x =- 5434 THEN
            sigmoid_f := 135;
        ELSIF x =- 5433 THEN
            sigmoid_f := 135;
        ELSIF x =- 5432 THEN
            sigmoid_f := 135;
        ELSIF x =- 5431 THEN
            sigmoid_f := 135;
        ELSIF x =- 5430 THEN
            sigmoid_f := 135;
        ELSIF x =- 5429 THEN
            sigmoid_f := 135;
        ELSIF x =- 5428 THEN
            sigmoid_f := 135;
        ELSIF x =- 5427 THEN
            sigmoid_f := 135;
        ELSIF x =- 5426 THEN
            sigmoid_f := 135;
        ELSIF x =- 5425 THEN
            sigmoid_f := 135;
        ELSIF x =- 5424 THEN
            sigmoid_f := 135;
        ELSIF x =- 5423 THEN
            sigmoid_f := 135;
        ELSIF x =- 5422 THEN
            sigmoid_f := 135;
        ELSIF x =- 5421 THEN
            sigmoid_f := 135;
        ELSIF x =- 5420 THEN
            sigmoid_f := 135;
        ELSIF x =- 5419 THEN
            sigmoid_f := 135;
        ELSIF x =- 5418 THEN
            sigmoid_f := 136;
        ELSIF x =- 5417 THEN
            sigmoid_f := 136;
        ELSIF x =- 5416 THEN
            sigmoid_f := 136;
        ELSIF x =- 5415 THEN
            sigmoid_f := 136;
        ELSIF x =- 5414 THEN
            sigmoid_f := 136;
        ELSIF x =- 5413 THEN
            sigmoid_f := 136;
        ELSIF x =- 5412 THEN
            sigmoid_f := 136;
        ELSIF x =- 5411 THEN
            sigmoid_f := 136;
        ELSIF x =- 5410 THEN
            sigmoid_f := 136;
        ELSIF x =- 5409 THEN
            sigmoid_f := 136;
        ELSIF x =- 5408 THEN
            sigmoid_f := 136;
        ELSIF x =- 5407 THEN
            sigmoid_f := 136;
        ELSIF x =- 5406 THEN
            sigmoid_f := 136;
        ELSIF x =- 5405 THEN
            sigmoid_f := 136;
        ELSIF x =- 5404 THEN
            sigmoid_f := 136;
        ELSIF x =- 5403 THEN
            sigmoid_f := 136;
        ELSIF x =- 5402 THEN
            sigmoid_f := 137;
        ELSIF x =- 5401 THEN
            sigmoid_f := 137;
        ELSIF x =- 5400 THEN
            sigmoid_f := 137;
        ELSIF x =- 5399 THEN
            sigmoid_f := 137;
        ELSIF x =- 5398 THEN
            sigmoid_f := 137;
        ELSIF x =- 5397 THEN
            sigmoid_f := 137;
        ELSIF x =- 5396 THEN
            sigmoid_f := 137;
        ELSIF x =- 5395 THEN
            sigmoid_f := 137;
        ELSIF x =- 5394 THEN
            sigmoid_f := 137;
        ELSIF x =- 5393 THEN
            sigmoid_f := 137;
        ELSIF x =- 5392 THEN
            sigmoid_f := 137;
        ELSIF x =- 5391 THEN
            sigmoid_f := 137;
        ELSIF x =- 5390 THEN
            sigmoid_f := 137;
        ELSIF x =- 5389 THEN
            sigmoid_f := 137;
        ELSIF x =- 5388 THEN
            sigmoid_f := 137;
        ELSIF x =- 5387 THEN
            sigmoid_f := 137;
        ELSIF x =- 5386 THEN
            sigmoid_f := 138;
        ELSIF x =- 5385 THEN
            sigmoid_f := 138;
        ELSIF x =- 5384 THEN
            sigmoid_f := 138;
        ELSIF x =- 5383 THEN
            sigmoid_f := 138;
        ELSIF x =- 5382 THEN
            sigmoid_f := 138;
        ELSIF x =- 5381 THEN
            sigmoid_f := 138;
        ELSIF x =- 5380 THEN
            sigmoid_f := 138;
        ELSIF x =- 5379 THEN
            sigmoid_f := 138;
        ELSIF x =- 5378 THEN
            sigmoid_f := 138;
        ELSIF x =- 5377 THEN
            sigmoid_f := 138;
        ELSIF x =- 5376 THEN
            sigmoid_f := 138;
        ELSIF x =- 5375 THEN
            sigmoid_f := 138;
        ELSIF x =- 5374 THEN
            sigmoid_f := 138;
        ELSIF x =- 5373 THEN
            sigmoid_f := 138;
        ELSIF x =- 5372 THEN
            sigmoid_f := 138;
        ELSIF x =- 5371 THEN
            sigmoid_f := 138;
        ELSIF x =- 5370 THEN
            sigmoid_f := 138;
        ELSIF x =- 5369 THEN
            sigmoid_f := 139;
        ELSIF x =- 5368 THEN
            sigmoid_f := 139;
        ELSIF x =- 5367 THEN
            sigmoid_f := 139;
        ELSIF x =- 5366 THEN
            sigmoid_f := 139;
        ELSIF x =- 5365 THEN
            sigmoid_f := 139;
        ELSIF x =- 5364 THEN
            sigmoid_f := 139;
        ELSIF x =- 5363 THEN
            sigmoid_f := 139;
        ELSIF x =- 5362 THEN
            sigmoid_f := 139;
        ELSIF x =- 5361 THEN
            sigmoid_f := 139;
        ELSIF x =- 5360 THEN
            sigmoid_f := 139;
        ELSIF x =- 5359 THEN
            sigmoid_f := 139;
        ELSIF x =- 5358 THEN
            sigmoid_f := 139;
        ELSIF x =- 5357 THEN
            sigmoid_f := 139;
        ELSIF x =- 5356 THEN
            sigmoid_f := 139;
        ELSIF x =- 5355 THEN
            sigmoid_f := 139;
        ELSIF x =- 5354 THEN
            sigmoid_f := 139;
        ELSIF x =- 5353 THEN
            sigmoid_f := 140;
        ELSIF x =- 5352 THEN
            sigmoid_f := 140;
        ELSIF x =- 5351 THEN
            sigmoid_f := 140;
        ELSIF x =- 5350 THEN
            sigmoid_f := 140;
        ELSIF x =- 5349 THEN
            sigmoid_f := 140;
        ELSIF x =- 5348 THEN
            sigmoid_f := 140;
        ELSIF x =- 5347 THEN
            sigmoid_f := 140;
        ELSIF x =- 5346 THEN
            sigmoid_f := 140;
        ELSIF x =- 5345 THEN
            sigmoid_f := 140;
        ELSIF x =- 5344 THEN
            sigmoid_f := 140;
        ELSIF x =- 5343 THEN
            sigmoid_f := 140;
        ELSIF x =- 5342 THEN
            sigmoid_f := 140;
        ELSIF x =- 5341 THEN
            sigmoid_f := 140;
        ELSIF x =- 5340 THEN
            sigmoid_f := 140;
        ELSIF x =- 5339 THEN
            sigmoid_f := 140;
        ELSIF x =- 5338 THEN
            sigmoid_f := 140;
        ELSIF x =- 5337 THEN
            sigmoid_f := 141;
        ELSIF x =- 5336 THEN
            sigmoid_f := 141;
        ELSIF x =- 5335 THEN
            sigmoid_f := 141;
        ELSIF x =- 5334 THEN
            sigmoid_f := 141;
        ELSIF x =- 5333 THEN
            sigmoid_f := 141;
        ELSIF x =- 5332 THEN
            sigmoid_f := 141;
        ELSIF x =- 5331 THEN
            sigmoid_f := 141;
        ELSIF x =- 5330 THEN
            sigmoid_f := 141;
        ELSIF x =- 5329 THEN
            sigmoid_f := 141;
        ELSIF x =- 5328 THEN
            sigmoid_f := 141;
        ELSIF x =- 5327 THEN
            sigmoid_f := 141;
        ELSIF x =- 5326 THEN
            sigmoid_f := 141;
        ELSIF x =- 5325 THEN
            sigmoid_f := 141;
        ELSIF x =- 5324 THEN
            sigmoid_f := 141;
        ELSIF x =- 5323 THEN
            sigmoid_f := 141;
        ELSIF x =- 5322 THEN
            sigmoid_f := 141;
        ELSIF x =- 5321 THEN
            sigmoid_f := 142;
        ELSIF x =- 5320 THEN
            sigmoid_f := 142;
        ELSIF x =- 5319 THEN
            sigmoid_f := 142;
        ELSIF x =- 5318 THEN
            sigmoid_f := 142;
        ELSIF x =- 5317 THEN
            sigmoid_f := 142;
        ELSIF x =- 5316 THEN
            sigmoid_f := 142;
        ELSIF x =- 5315 THEN
            sigmoid_f := 142;
        ELSIF x =- 5314 THEN
            sigmoid_f := 142;
        ELSIF x =- 5313 THEN
            sigmoid_f := 142;
        ELSIF x =- 5312 THEN
            sigmoid_f := 142;
        ELSIF x =- 5311 THEN
            sigmoid_f := 142;
        ELSIF x =- 5310 THEN
            sigmoid_f := 142;
        ELSIF x =- 5309 THEN
            sigmoid_f := 142;
        ELSIF x =- 5308 THEN
            sigmoid_f := 142;
        ELSIF x =- 5307 THEN
            sigmoid_f := 142;
        ELSIF x =- 5306 THEN
            sigmoid_f := 142;
        ELSIF x =- 5305 THEN
            sigmoid_f := 143;
        ELSIF x =- 5304 THEN
            sigmoid_f := 143;
        ELSIF x =- 5303 THEN
            sigmoid_f := 143;
        ELSIF x =- 5302 THEN
            sigmoid_f := 143;
        ELSIF x =- 5301 THEN
            sigmoid_f := 143;
        ELSIF x =- 5300 THEN
            sigmoid_f := 143;
        ELSIF x =- 5299 THEN
            sigmoid_f := 143;
        ELSIF x =- 5298 THEN
            sigmoid_f := 143;
        ELSIF x =- 5297 THEN
            sigmoid_f := 143;
        ELSIF x =- 5296 THEN
            sigmoid_f := 143;
        ELSIF x =- 5295 THEN
            sigmoid_f := 143;
        ELSIF x =- 5294 THEN
            sigmoid_f := 143;
        ELSIF x =- 5293 THEN
            sigmoid_f := 143;
        ELSIF x =- 5292 THEN
            sigmoid_f := 143;
        ELSIF x =- 5291 THEN
            sigmoid_f := 143;
        ELSIF x =- 5290 THEN
            sigmoid_f := 143;
        ELSIF x =- 5289 THEN
            sigmoid_f := 144;
        ELSIF x =- 5288 THEN
            sigmoid_f := 144;
        ELSIF x =- 5287 THEN
            sigmoid_f := 144;
        ELSIF x =- 5286 THEN
            sigmoid_f := 144;
        ELSIF x =- 5285 THEN
            sigmoid_f := 144;
        ELSIF x =- 5284 THEN
            sigmoid_f := 144;
        ELSIF x =- 5283 THEN
            sigmoid_f := 144;
        ELSIF x =- 5282 THEN
            sigmoid_f := 144;
        ELSIF x =- 5281 THEN
            sigmoid_f := 144;
        ELSIF x =- 5280 THEN
            sigmoid_f := 144;
        ELSIF x =- 5279 THEN
            sigmoid_f := 144;
        ELSIF x =- 5278 THEN
            sigmoid_f := 144;
        ELSIF x =- 5277 THEN
            sigmoid_f := 144;
        ELSIF x =- 5276 THEN
            sigmoid_f := 144;
        ELSIF x =- 5275 THEN
            sigmoid_f := 144;
        ELSIF x =- 5274 THEN
            sigmoid_f := 144;
        ELSIF x =- 5273 THEN
            sigmoid_f := 145;
        ELSIF x =- 5272 THEN
            sigmoid_f := 145;
        ELSIF x =- 5271 THEN
            sigmoid_f := 145;
        ELSIF x =- 5270 THEN
            sigmoid_f := 145;
        ELSIF x =- 5269 THEN
            sigmoid_f := 145;
        ELSIF x =- 5268 THEN
            sigmoid_f := 145;
        ELSIF x =- 5267 THEN
            sigmoid_f := 145;
        ELSIF x =- 5266 THEN
            sigmoid_f := 145;
        ELSIF x =- 5265 THEN
            sigmoid_f := 145;
        ELSIF x =- 5264 THEN
            sigmoid_f := 145;
        ELSIF x =- 5263 THEN
            sigmoid_f := 145;
        ELSIF x =- 5262 THEN
            sigmoid_f := 145;
        ELSIF x =- 5261 THEN
            sigmoid_f := 145;
        ELSIF x =- 5260 THEN
            sigmoid_f := 145;
        ELSIF x =- 5259 THEN
            sigmoid_f := 145;
        ELSIF x =- 5258 THEN
            sigmoid_f := 145;
        ELSIF x =- 5257 THEN
            sigmoid_f := 146;
        ELSIF x =- 5256 THEN
            sigmoid_f := 146;
        ELSIF x =- 5255 THEN
            sigmoid_f := 146;
        ELSIF x =- 5254 THEN
            sigmoid_f := 146;
        ELSIF x =- 5253 THEN
            sigmoid_f := 146;
        ELSIF x =- 5252 THEN
            sigmoid_f := 146;
        ELSIF x =- 5251 THEN
            sigmoid_f := 146;
        ELSIF x =- 5250 THEN
            sigmoid_f := 146;
        ELSIF x =- 5249 THEN
            sigmoid_f := 146;
        ELSIF x =- 5248 THEN
            sigmoid_f := 146;
        ELSIF x =- 5247 THEN
            sigmoid_f := 146;
        ELSIF x =- 5246 THEN
            sigmoid_f := 146;
        ELSIF x =- 5245 THEN
            sigmoid_f := 146;
        ELSIF x =- 5244 THEN
            sigmoid_f := 146;
        ELSIF x =- 5243 THEN
            sigmoid_f := 146;
        ELSIF x =- 5242 THEN
            sigmoid_f := 146;
        ELSIF x =- 5241 THEN
            sigmoid_f := 146;
        ELSIF x =- 5240 THEN
            sigmoid_f := 147;
        ELSIF x =- 5239 THEN
            sigmoid_f := 147;
        ELSIF x =- 5238 THEN
            sigmoid_f := 147;
        ELSIF x =- 5237 THEN
            sigmoid_f := 147;
        ELSIF x =- 5236 THEN
            sigmoid_f := 147;
        ELSIF x =- 5235 THEN
            sigmoid_f := 147;
        ELSIF x =- 5234 THEN
            sigmoid_f := 147;
        ELSIF x =- 5233 THEN
            sigmoid_f := 147;
        ELSIF x =- 5232 THEN
            sigmoid_f := 147;
        ELSIF x =- 5231 THEN
            sigmoid_f := 147;
        ELSIF x =- 5230 THEN
            sigmoid_f := 147;
        ELSIF x =- 5229 THEN
            sigmoid_f := 147;
        ELSIF x =- 5228 THEN
            sigmoid_f := 147;
        ELSIF x =- 5227 THEN
            sigmoid_f := 147;
        ELSIF x =- 5226 THEN
            sigmoid_f := 147;
        ELSIF x =- 5225 THEN
            sigmoid_f := 147;
        ELSIF x =- 5224 THEN
            sigmoid_f := 148;
        ELSIF x =- 5223 THEN
            sigmoid_f := 148;
        ELSIF x =- 5222 THEN
            sigmoid_f := 148;
        ELSIF x =- 5221 THEN
            sigmoid_f := 148;
        ELSIF x =- 5220 THEN
            sigmoid_f := 148;
        ELSIF x =- 5219 THEN
            sigmoid_f := 148;
        ELSIF x =- 5218 THEN
            sigmoid_f := 148;
        ELSIF x =- 5217 THEN
            sigmoid_f := 148;
        ELSIF x =- 5216 THEN
            sigmoid_f := 148;
        ELSIF x =- 5215 THEN
            sigmoid_f := 148;
        ELSIF x =- 5214 THEN
            sigmoid_f := 148;
        ELSIF x =- 5213 THEN
            sigmoid_f := 148;
        ELSIF x =- 5212 THEN
            sigmoid_f := 148;
        ELSIF x =- 5211 THEN
            sigmoid_f := 148;
        ELSIF x =- 5210 THEN
            sigmoid_f := 148;
        ELSIF x =- 5209 THEN
            sigmoid_f := 148;
        ELSIF x =- 5208 THEN
            sigmoid_f := 149;
        ELSIF x =- 5207 THEN
            sigmoid_f := 149;
        ELSIF x =- 5206 THEN
            sigmoid_f := 149;
        ELSIF x =- 5205 THEN
            sigmoid_f := 149;
        ELSIF x =- 5204 THEN
            sigmoid_f := 149;
        ELSIF x =- 5203 THEN
            sigmoid_f := 149;
        ELSIF x =- 5202 THEN
            sigmoid_f := 149;
        ELSIF x =- 5201 THEN
            sigmoid_f := 149;
        ELSIF x =- 5200 THEN
            sigmoid_f := 149;
        ELSIF x =- 5199 THEN
            sigmoid_f := 149;
        ELSIF x =- 5198 THEN
            sigmoid_f := 149;
        ELSIF x =- 5197 THEN
            sigmoid_f := 149;
        ELSIF x =- 5196 THEN
            sigmoid_f := 149;
        ELSIF x =- 5195 THEN
            sigmoid_f := 149;
        ELSIF x =- 5194 THEN
            sigmoid_f := 149;
        ELSIF x =- 5193 THEN
            sigmoid_f := 149;
        ELSIF x =- 5192 THEN
            sigmoid_f := 150;
        ELSIF x =- 5191 THEN
            sigmoid_f := 150;
        ELSIF x =- 5190 THEN
            sigmoid_f := 150;
        ELSIF x =- 5189 THEN
            sigmoid_f := 150;
        ELSIF x =- 5188 THEN
            sigmoid_f := 150;
        ELSIF x =- 5187 THEN
            sigmoid_f := 150;
        ELSIF x =- 5186 THEN
            sigmoid_f := 150;
        ELSIF x =- 5185 THEN
            sigmoid_f := 150;
        ELSIF x =- 5184 THEN
            sigmoid_f := 150;
        ELSIF x =- 5183 THEN
            sigmoid_f := 150;
        ELSIF x =- 5182 THEN
            sigmoid_f := 150;
        ELSIF x =- 5181 THEN
            sigmoid_f := 150;
        ELSIF x =- 5180 THEN
            sigmoid_f := 150;
        ELSIF x =- 5179 THEN
            sigmoid_f := 150;
        ELSIF x =- 5178 THEN
            sigmoid_f := 150;
        ELSIF x =- 5177 THEN
            sigmoid_f := 150;
        ELSIF x =- 5176 THEN
            sigmoid_f := 151;
        ELSIF x =- 5175 THEN
            sigmoid_f := 151;
        ELSIF x =- 5174 THEN
            sigmoid_f := 151;
        ELSIF x =- 5173 THEN
            sigmoid_f := 151;
        ELSIF x =- 5172 THEN
            sigmoid_f := 151;
        ELSIF x =- 5171 THEN
            sigmoid_f := 151;
        ELSIF x =- 5170 THEN
            sigmoid_f := 151;
        ELSIF x =- 5169 THEN
            sigmoid_f := 151;
        ELSIF x =- 5168 THEN
            sigmoid_f := 151;
        ELSIF x =- 5167 THEN
            sigmoid_f := 151;
        ELSIF x =- 5166 THEN
            sigmoid_f := 151;
        ELSIF x =- 5165 THEN
            sigmoid_f := 151;
        ELSIF x =- 5164 THEN
            sigmoid_f := 151;
        ELSIF x =- 5163 THEN
            sigmoid_f := 151;
        ELSIF x =- 5162 THEN
            sigmoid_f := 151;
        ELSIF x =- 5161 THEN
            sigmoid_f := 151;
        ELSIF x =- 5160 THEN
            sigmoid_f := 152;
        ELSIF x =- 5159 THEN
            sigmoid_f := 152;
        ELSIF x =- 5158 THEN
            sigmoid_f := 152;
        ELSIF x =- 5157 THEN
            sigmoid_f := 152;
        ELSIF x =- 5156 THEN
            sigmoid_f := 152;
        ELSIF x =- 5155 THEN
            sigmoid_f := 152;
        ELSIF x =- 5154 THEN
            sigmoid_f := 152;
        ELSIF x =- 5153 THEN
            sigmoid_f := 152;
        ELSIF x =- 5152 THEN
            sigmoid_f := 152;
        ELSIF x =- 5151 THEN
            sigmoid_f := 152;
        ELSIF x =- 5150 THEN
            sigmoid_f := 152;
        ELSIF x =- 5149 THEN
            sigmoid_f := 152;
        ELSIF x =- 5148 THEN
            sigmoid_f := 152;
        ELSIF x =- 5147 THEN
            sigmoid_f := 152;
        ELSIF x =- 5146 THEN
            sigmoid_f := 152;
        ELSIF x =- 5145 THEN
            sigmoid_f := 152;
        ELSIF x =- 5144 THEN
            sigmoid_f := 153;
        ELSIF x =- 5143 THEN
            sigmoid_f := 153;
        ELSIF x =- 5142 THEN
            sigmoid_f := 153;
        ELSIF x =- 5141 THEN
            sigmoid_f := 153;
        ELSIF x =- 5140 THEN
            sigmoid_f := 153;
        ELSIF x =- 5139 THEN
            sigmoid_f := 153;
        ELSIF x =- 5138 THEN
            sigmoid_f := 153;
        ELSIF x =- 5137 THEN
            sigmoid_f := 153;
        ELSIF x =- 5136 THEN
            sigmoid_f := 153;
        ELSIF x =- 5135 THEN
            sigmoid_f := 153;
        ELSIF x =- 5134 THEN
            sigmoid_f := 153;
        ELSIF x =- 5133 THEN
            sigmoid_f := 153;
        ELSIF x =- 5132 THEN
            sigmoid_f := 153;
        ELSIF x =- 5131 THEN
            sigmoid_f := 153;
        ELSIF x =- 5130 THEN
            sigmoid_f := 153;
        ELSIF x =- 5129 THEN
            sigmoid_f := 153;
        ELSIF x =- 5128 THEN
            sigmoid_f := 154;
        ELSIF x =- 5127 THEN
            sigmoid_f := 154;
        ELSIF x =- 5126 THEN
            sigmoid_f := 154;
        ELSIF x =- 5125 THEN
            sigmoid_f := 154;
        ELSIF x =- 5124 THEN
            sigmoid_f := 154;
        ELSIF x =- 5123 THEN
            sigmoid_f := 154;
        ELSIF x =- 5122 THEN
            sigmoid_f := 154;
        ELSIF x =- 5121 THEN
            sigmoid_f := 154;
        ELSIF x =- 5120 THEN
            sigmoid_f := 154;
        ELSIF x =- 5119 THEN
            sigmoid_f := 154;
        ELSIF x =- 5118 THEN
            sigmoid_f := 154;
        ELSIF x =- 5117 THEN
            sigmoid_f := 154;
        ELSIF x =- 5116 THEN
            sigmoid_f := 154;
        ELSIF x =- 5115 THEN
            sigmoid_f := 154;
        ELSIF x =- 5114 THEN
            sigmoid_f := 154;
        ELSIF x =- 5113 THEN
            sigmoid_f := 155;
        ELSIF x =- 5112 THEN
            sigmoid_f := 155;
        ELSIF x =- 5111 THEN
            sigmoid_f := 155;
        ELSIF x =- 5110 THEN
            sigmoid_f := 155;
        ELSIF x =- 5109 THEN
            sigmoid_f := 155;
        ELSIF x =- 5108 THEN
            sigmoid_f := 155;
        ELSIF x =- 5107 THEN
            sigmoid_f := 155;
        ELSIF x =- 5106 THEN
            sigmoid_f := 155;
        ELSIF x =- 5105 THEN
            sigmoid_f := 155;
        ELSIF x =- 5104 THEN
            sigmoid_f := 155;
        ELSIF x =- 5103 THEN
            sigmoid_f := 155;
        ELSIF x =- 5102 THEN
            sigmoid_f := 155;
        ELSIF x =- 5101 THEN
            sigmoid_f := 155;
        ELSIF x =- 5100 THEN
            sigmoid_f := 156;
        ELSIF x =- 5099 THEN
            sigmoid_f := 156;
        ELSIF x =- 5098 THEN
            sigmoid_f := 156;
        ELSIF x =- 5097 THEN
            sigmoid_f := 156;
        ELSIF x =- 5096 THEN
            sigmoid_f := 156;
        ELSIF x =- 5095 THEN
            sigmoid_f := 156;
        ELSIF x =- 5094 THEN
            sigmoid_f := 156;
        ELSIF x =- 5093 THEN
            sigmoid_f := 156;
        ELSIF x =- 5092 THEN
            sigmoid_f := 156;
        ELSIF x =- 5091 THEN
            sigmoid_f := 156;
        ELSIF x =- 5090 THEN
            sigmoid_f := 156;
        ELSIF x =- 5089 THEN
            sigmoid_f := 156;
        ELSIF x =- 5088 THEN
            sigmoid_f := 157;
        ELSIF x =- 5087 THEN
            sigmoid_f := 157;
        ELSIF x =- 5086 THEN
            sigmoid_f := 157;
        ELSIF x =- 5085 THEN
            sigmoid_f := 157;
        ELSIF x =- 5084 THEN
            sigmoid_f := 157;
        ELSIF x =- 5083 THEN
            sigmoid_f := 157;
        ELSIF x =- 5082 THEN
            sigmoid_f := 157;
        ELSIF x =- 5081 THEN
            sigmoid_f := 157;
        ELSIF x =- 5080 THEN
            sigmoid_f := 157;
        ELSIF x =- 5079 THEN
            sigmoid_f := 157;
        ELSIF x =- 5078 THEN
            sigmoid_f := 157;
        ELSIF x =- 5077 THEN
            sigmoid_f := 157;
        ELSIF x =- 5076 THEN
            sigmoid_f := 157;
        ELSIF x =- 5075 THEN
            sigmoid_f := 158;
        ELSIF x =- 5074 THEN
            sigmoid_f := 158;
        ELSIF x =- 5073 THEN
            sigmoid_f := 158;
        ELSIF x =- 5072 THEN
            sigmoid_f := 158;
        ELSIF x =- 5071 THEN
            sigmoid_f := 158;
        ELSIF x =- 5070 THEN
            sigmoid_f := 158;
        ELSIF x =- 5069 THEN
            sigmoid_f := 158;
        ELSIF x =- 5068 THEN
            sigmoid_f := 158;
        ELSIF x =- 5067 THEN
            sigmoid_f := 158;
        ELSIF x =- 5066 THEN
            sigmoid_f := 158;
        ELSIF x =- 5065 THEN
            sigmoid_f := 158;
        ELSIF x =- 5064 THEN
            sigmoid_f := 158;
        ELSIF x =- 5063 THEN
            sigmoid_f := 158;
        ELSIF x =- 5062 THEN
            sigmoid_f := 159;
        ELSIF x =- 5061 THEN
            sigmoid_f := 159;
        ELSIF x =- 5060 THEN
            sigmoid_f := 159;
        ELSIF x =- 5059 THEN
            sigmoid_f := 159;
        ELSIF x =- 5058 THEN
            sigmoid_f := 159;
        ELSIF x =- 5057 THEN
            sigmoid_f := 159;
        ELSIF x =- 5056 THEN
            sigmoid_f := 159;
        ELSIF x =- 5055 THEN
            sigmoid_f := 159;
        ELSIF x =- 5054 THEN
            sigmoid_f := 159;
        ELSIF x =- 5053 THEN
            sigmoid_f := 159;
        ELSIF x =- 5052 THEN
            sigmoid_f := 159;
        ELSIF x =- 5051 THEN
            sigmoid_f := 159;
        ELSIF x =- 5050 THEN
            sigmoid_f := 160;
        ELSIF x =- 5049 THEN
            sigmoid_f := 160;
        ELSIF x =- 5048 THEN
            sigmoid_f := 160;
        ELSIF x =- 5047 THEN
            sigmoid_f := 160;
        ELSIF x =- 5046 THEN
            sigmoid_f := 160;
        ELSIF x =- 5045 THEN
            sigmoid_f := 160;
        ELSIF x =- 5044 THEN
            sigmoid_f := 160;
        ELSIF x =- 5043 THEN
            sigmoid_f := 160;
        ELSIF x =- 5042 THEN
            sigmoid_f := 160;
        ELSIF x =- 5041 THEN
            sigmoid_f := 160;
        ELSIF x =- 5040 THEN
            sigmoid_f := 160;
        ELSIF x =- 5039 THEN
            sigmoid_f := 160;
        ELSIF x =- 5038 THEN
            sigmoid_f := 160;
        ELSIF x =- 5037 THEN
            sigmoid_f := 161;
        ELSIF x =- 5036 THEN
            sigmoid_f := 161;
        ELSIF x =- 5035 THEN
            sigmoid_f := 161;
        ELSIF x =- 5034 THEN
            sigmoid_f := 161;
        ELSIF x =- 5033 THEN
            sigmoid_f := 161;
        ELSIF x =- 5032 THEN
            sigmoid_f := 161;
        ELSIF x =- 5031 THEN
            sigmoid_f := 161;
        ELSIF x =- 5030 THEN
            sigmoid_f := 161;
        ELSIF x =- 5029 THEN
            sigmoid_f := 161;
        ELSIF x =- 5028 THEN
            sigmoid_f := 161;
        ELSIF x =- 5027 THEN
            sigmoid_f := 161;
        ELSIF x =- 5026 THEN
            sigmoid_f := 161;
        ELSIF x =- 5025 THEN
            sigmoid_f := 161;
        ELSIF x =- 5024 THEN
            sigmoid_f := 162;
        ELSIF x =- 5023 THEN
            sigmoid_f := 162;
        ELSIF x =- 5022 THEN
            sigmoid_f := 162;
        ELSIF x =- 5021 THEN
            sigmoid_f := 162;
        ELSIF x =- 5020 THEN
            sigmoid_f := 162;
        ELSIF x =- 5019 THEN
            sigmoid_f := 162;
        ELSIF x =- 5018 THEN
            sigmoid_f := 162;
        ELSIF x =- 5017 THEN
            sigmoid_f := 162;
        ELSIF x =- 5016 THEN
            sigmoid_f := 162;
        ELSIF x =- 5015 THEN
            sigmoid_f := 162;
        ELSIF x =- 5014 THEN
            sigmoid_f := 162;
        ELSIF x =- 5013 THEN
            sigmoid_f := 162;
        ELSIF x =- 5012 THEN
            sigmoid_f := 162;
        ELSIF x =- 5011 THEN
            sigmoid_f := 163;
        ELSIF x =- 5010 THEN
            sigmoid_f := 163;
        ELSIF x =- 5009 THEN
            sigmoid_f := 163;
        ELSIF x =- 5008 THEN
            sigmoid_f := 163;
        ELSIF x =- 5007 THEN
            sigmoid_f := 163;
        ELSIF x =- 5006 THEN
            sigmoid_f := 163;
        ELSIF x =- 5005 THEN
            sigmoid_f := 163;
        ELSIF x =- 5004 THEN
            sigmoid_f := 163;
        ELSIF x =- 5003 THEN
            sigmoid_f := 163;
        ELSIF x =- 5002 THEN
            sigmoid_f := 163;
        ELSIF x =- 5001 THEN
            sigmoid_f := 163;
        ELSIF x =- 5000 THEN
            sigmoid_f := 163;
        ELSIF x =- 4999 THEN
            sigmoid_f := 164;
        ELSIF x =- 4998 THEN
            sigmoid_f := 164;
        ELSIF x =- 4997 THEN
            sigmoid_f := 164;
        ELSIF x =- 4996 THEN
            sigmoid_f := 164;
        ELSIF x =- 4995 THEN
            sigmoid_f := 164;
        ELSIF x =- 4994 THEN
            sigmoid_f := 164;
        ELSIF x =- 4993 THEN
            sigmoid_f := 164;
        ELSIF x =- 4992 THEN
            sigmoid_f := 164;
        ELSIF x =- 4991 THEN
            sigmoid_f := 164;
        ELSIF x =- 4990 THEN
            sigmoid_f := 164;
        ELSIF x =- 4989 THEN
            sigmoid_f := 164;
        ELSIF x =- 4988 THEN
            sigmoid_f := 164;
        ELSIF x =- 4987 THEN
            sigmoid_f := 164;
        ELSIF x =- 4986 THEN
            sigmoid_f := 165;
        ELSIF x =- 4985 THEN
            sigmoid_f := 165;
        ELSIF x =- 4984 THEN
            sigmoid_f := 165;
        ELSIF x =- 4983 THEN
            sigmoid_f := 165;
        ELSIF x =- 4982 THEN
            sigmoid_f := 165;
        ELSIF x =- 4981 THEN
            sigmoid_f := 165;
        ELSIF x =- 4980 THEN
            sigmoid_f := 165;
        ELSIF x =- 4979 THEN
            sigmoid_f := 165;
        ELSIF x =- 4978 THEN
            sigmoid_f := 165;
        ELSIF x =- 4977 THEN
            sigmoid_f := 165;
        ELSIF x =- 4976 THEN
            sigmoid_f := 165;
        ELSIF x =- 4975 THEN
            sigmoid_f := 165;
        ELSIF x =- 4974 THEN
            sigmoid_f := 165;
        ELSIF x =- 4973 THEN
            sigmoid_f := 166;
        ELSIF x =- 4972 THEN
            sigmoid_f := 166;
        ELSIF x =- 4971 THEN
            sigmoid_f := 166;
        ELSIF x =- 4970 THEN
            sigmoid_f := 166;
        ELSIF x =- 4969 THEN
            sigmoid_f := 166;
        ELSIF x =- 4968 THEN
            sigmoid_f := 166;
        ELSIF x =- 4967 THEN
            sigmoid_f := 166;
        ELSIF x =- 4966 THEN
            sigmoid_f := 166;
        ELSIF x =- 4965 THEN
            sigmoid_f := 166;
        ELSIF x =- 4964 THEN
            sigmoid_f := 166;
        ELSIF x =- 4963 THEN
            sigmoid_f := 166;
        ELSIF x =- 4962 THEN
            sigmoid_f := 166;
        ELSIF x =- 4961 THEN
            sigmoid_f := 166;
        ELSIF x =- 4960 THEN
            sigmoid_f := 167;
        ELSIF x =- 4959 THEN
            sigmoid_f := 167;
        ELSIF x =- 4958 THEN
            sigmoid_f := 167;
        ELSIF x =- 4957 THEN
            sigmoid_f := 167;
        ELSIF x =- 4956 THEN
            sigmoid_f := 167;
        ELSIF x =- 4955 THEN
            sigmoid_f := 167;
        ELSIF x =- 4954 THEN
            sigmoid_f := 167;
        ELSIF x =- 4953 THEN
            sigmoid_f := 167;
        ELSIF x =- 4952 THEN
            sigmoid_f := 167;
        ELSIF x =- 4951 THEN
            sigmoid_f := 167;
        ELSIF x =- 4950 THEN
            sigmoid_f := 167;
        ELSIF x =- 4949 THEN
            sigmoid_f := 167;
        ELSIF x =- 4948 THEN
            sigmoid_f := 168;
        ELSIF x =- 4947 THEN
            sigmoid_f := 168;
        ELSIF x =- 4946 THEN
            sigmoid_f := 168;
        ELSIF x =- 4945 THEN
            sigmoid_f := 168;
        ELSIF x =- 4944 THEN
            sigmoid_f := 168;
        ELSIF x =- 4943 THEN
            sigmoid_f := 168;
        ELSIF x =- 4942 THEN
            sigmoid_f := 168;
        ELSIF x =- 4941 THEN
            sigmoid_f := 168;
        ELSIF x =- 4940 THEN
            sigmoid_f := 168;
        ELSIF x =- 4939 THEN
            sigmoid_f := 168;
        ELSIF x =- 4938 THEN
            sigmoid_f := 168;
        ELSIF x =- 4937 THEN
            sigmoid_f := 168;
        ELSIF x =- 4936 THEN
            sigmoid_f := 168;
        ELSIF x =- 4935 THEN
            sigmoid_f := 169;
        ELSIF x =- 4934 THEN
            sigmoid_f := 169;
        ELSIF x =- 4933 THEN
            sigmoid_f := 169;
        ELSIF x =- 4932 THEN
            sigmoid_f := 169;
        ELSIF x =- 4931 THEN
            sigmoid_f := 169;
        ELSIF x =- 4930 THEN
            sigmoid_f := 169;
        ELSIF x =- 4929 THEN
            sigmoid_f := 169;
        ELSIF x =- 4928 THEN
            sigmoid_f := 169;
        ELSIF x =- 4927 THEN
            sigmoid_f := 169;
        ELSIF x =- 4926 THEN
            sigmoid_f := 169;
        ELSIF x =- 4925 THEN
            sigmoid_f := 169;
        ELSIF x =- 4924 THEN
            sigmoid_f := 169;
        ELSIF x =- 4923 THEN
            sigmoid_f := 169;
        ELSIF x =- 4922 THEN
            sigmoid_f := 170;
        ELSIF x =- 4921 THEN
            sigmoid_f := 170;
        ELSIF x =- 4920 THEN
            sigmoid_f := 170;
        ELSIF x =- 4919 THEN
            sigmoid_f := 170;
        ELSIF x =- 4918 THEN
            sigmoid_f := 170;
        ELSIF x =- 4917 THEN
            sigmoid_f := 170;
        ELSIF x =- 4916 THEN
            sigmoid_f := 170;
        ELSIF x =- 4915 THEN
            sigmoid_f := 170;
        ELSIF x =- 4914 THEN
            sigmoid_f := 170;
        ELSIF x =- 4913 THEN
            sigmoid_f := 170;
        ELSIF x =- 4912 THEN
            sigmoid_f := 170;
        ELSIF x =- 4911 THEN
            sigmoid_f := 170;
        ELSIF x =- 4910 THEN
            sigmoid_f := 171;
        ELSIF x =- 4909 THEN
            sigmoid_f := 171;
        ELSIF x =- 4908 THEN
            sigmoid_f := 171;
        ELSIF x =- 4907 THEN
            sigmoid_f := 171;
        ELSIF x =- 4906 THEN
            sigmoid_f := 171;
        ELSIF x =- 4905 THEN
            sigmoid_f := 171;
        ELSIF x =- 4904 THEN
            sigmoid_f := 171;
        ELSIF x =- 4903 THEN
            sigmoid_f := 171;
        ELSIF x =- 4902 THEN
            sigmoid_f := 171;
        ELSIF x =- 4901 THEN
            sigmoid_f := 171;
        ELSIF x =- 4900 THEN
            sigmoid_f := 171;
        ELSIF x =- 4899 THEN
            sigmoid_f := 171;
        ELSIF x =- 4898 THEN
            sigmoid_f := 171;
        ELSIF x =- 4897 THEN
            sigmoid_f := 172;
        ELSIF x =- 4896 THEN
            sigmoid_f := 172;
        ELSIF x =- 4895 THEN
            sigmoid_f := 172;
        ELSIF x =- 4894 THEN
            sigmoid_f := 172;
        ELSIF x =- 4893 THEN
            sigmoid_f := 172;
        ELSIF x =- 4892 THEN
            sigmoid_f := 172;
        ELSIF x =- 4891 THEN
            sigmoid_f := 172;
        ELSIF x =- 4890 THEN
            sigmoid_f := 172;
        ELSIF x =- 4889 THEN
            sigmoid_f := 172;
        ELSIF x =- 4888 THEN
            sigmoid_f := 172;
        ELSIF x =- 4887 THEN
            sigmoid_f := 172;
        ELSIF x =- 4886 THEN
            sigmoid_f := 172;
        ELSIF x =- 4885 THEN
            sigmoid_f := 172;
        ELSIF x =- 4884 THEN
            sigmoid_f := 173;
        ELSIF x =- 4883 THEN
            sigmoid_f := 173;
        ELSIF x =- 4882 THEN
            sigmoid_f := 173;
        ELSIF x =- 4881 THEN
            sigmoid_f := 173;
        ELSIF x =- 4880 THEN
            sigmoid_f := 173;
        ELSIF x =- 4879 THEN
            sigmoid_f := 173;
        ELSIF x =- 4878 THEN
            sigmoid_f := 173;
        ELSIF x =- 4877 THEN
            sigmoid_f := 173;
        ELSIF x =- 4876 THEN
            sigmoid_f := 173;
        ELSIF x =- 4875 THEN
            sigmoid_f := 173;
        ELSIF x =- 4874 THEN
            sigmoid_f := 173;
        ELSIF x =- 4873 THEN
            sigmoid_f := 173;
        ELSIF x =- 4872 THEN
            sigmoid_f := 173;
        ELSIF x =- 4871 THEN
            sigmoid_f := 174;
        ELSIF x =- 4870 THEN
            sigmoid_f := 174;
        ELSIF x =- 4869 THEN
            sigmoid_f := 174;
        ELSIF x =- 4868 THEN
            sigmoid_f := 174;
        ELSIF x =- 4867 THEN
            sigmoid_f := 174;
        ELSIF x =- 4866 THEN
            sigmoid_f := 174;
        ELSIF x =- 4865 THEN
            sigmoid_f := 174;
        ELSIF x =- 4864 THEN
            sigmoid_f := 174;
        ELSIF x =- 4863 THEN
            sigmoid_f := 174;
        ELSIF x =- 4862 THEN
            sigmoid_f := 174;
        ELSIF x =- 4861 THEN
            sigmoid_f := 174;
        ELSIF x =- 4860 THEN
            sigmoid_f := 174;
        ELSIF x =- 4859 THEN
            sigmoid_f := 175;
        ELSIF x =- 4858 THEN
            sigmoid_f := 175;
        ELSIF x =- 4857 THEN
            sigmoid_f := 175;
        ELSIF x =- 4856 THEN
            sigmoid_f := 175;
        ELSIF x =- 4855 THEN
            sigmoid_f := 175;
        ELSIF x =- 4854 THEN
            sigmoid_f := 175;
        ELSIF x =- 4853 THEN
            sigmoid_f := 175;
        ELSIF x =- 4852 THEN
            sigmoid_f := 175;
        ELSIF x =- 4851 THEN
            sigmoid_f := 175;
        ELSIF x =- 4850 THEN
            sigmoid_f := 175;
        ELSIF x =- 4849 THEN
            sigmoid_f := 175;
        ELSIF x =- 4848 THEN
            sigmoid_f := 175;
        ELSIF x =- 4847 THEN
            sigmoid_f := 175;
        ELSIF x =- 4846 THEN
            sigmoid_f := 176;
        ELSIF x =- 4845 THEN
            sigmoid_f := 176;
        ELSIF x =- 4844 THEN
            sigmoid_f := 176;
        ELSIF x =- 4843 THEN
            sigmoid_f := 176;
        ELSIF x =- 4842 THEN
            sigmoid_f := 176;
        ELSIF x =- 4841 THEN
            sigmoid_f := 176;
        ELSIF x =- 4840 THEN
            sigmoid_f := 176;
        ELSIF x =- 4839 THEN
            sigmoid_f := 176;
        ELSIF x =- 4838 THEN
            sigmoid_f := 176;
        ELSIF x =- 4837 THEN
            sigmoid_f := 176;
        ELSIF x =- 4836 THEN
            sigmoid_f := 176;
        ELSIF x =- 4835 THEN
            sigmoid_f := 176;
        ELSIF x =- 4834 THEN
            sigmoid_f := 176;
        ELSIF x =- 4833 THEN
            sigmoid_f := 177;
        ELSIF x =- 4832 THEN
            sigmoid_f := 177;
        ELSIF x =- 4831 THEN
            sigmoid_f := 177;
        ELSIF x =- 4830 THEN
            sigmoid_f := 177;
        ELSIF x =- 4829 THEN
            sigmoid_f := 177;
        ELSIF x =- 4828 THEN
            sigmoid_f := 177;
        ELSIF x =- 4827 THEN
            sigmoid_f := 177;
        ELSIF x =- 4826 THEN
            sigmoid_f := 177;
        ELSIF x =- 4825 THEN
            sigmoid_f := 177;
        ELSIF x =- 4824 THEN
            sigmoid_f := 177;
        ELSIF x =- 4823 THEN
            sigmoid_f := 177;
        ELSIF x =- 4822 THEN
            sigmoid_f := 177;
        ELSIF x =- 4821 THEN
            sigmoid_f := 178;
        ELSIF x =- 4820 THEN
            sigmoid_f := 178;
        ELSIF x =- 4819 THEN
            sigmoid_f := 178;
        ELSIF x =- 4818 THEN
            sigmoid_f := 178;
        ELSIF x =- 4817 THEN
            sigmoid_f := 178;
        ELSIF x =- 4816 THEN
            sigmoid_f := 178;
        ELSIF x =- 4815 THEN
            sigmoid_f := 178;
        ELSIF x =- 4814 THEN
            sigmoid_f := 178;
        ELSIF x =- 4813 THEN
            sigmoid_f := 178;
        ELSIF x =- 4812 THEN
            sigmoid_f := 178;
        ELSIF x =- 4811 THEN
            sigmoid_f := 178;
        ELSIF x =- 4810 THEN
            sigmoid_f := 178;
        ELSIF x =- 4809 THEN
            sigmoid_f := 178;
        ELSIF x =- 4808 THEN
            sigmoid_f := 179;
        ELSIF x =- 4807 THEN
            sigmoid_f := 179;
        ELSIF x =- 4806 THEN
            sigmoid_f := 179;
        ELSIF x =- 4805 THEN
            sigmoid_f := 179;
        ELSIF x =- 4804 THEN
            sigmoid_f := 179;
        ELSIF x =- 4803 THEN
            sigmoid_f := 179;
        ELSIF x =- 4802 THEN
            sigmoid_f := 179;
        ELSIF x =- 4801 THEN
            sigmoid_f := 179;
        ELSIF x =- 4800 THEN
            sigmoid_f := 179;
        ELSIF x =- 4799 THEN
            sigmoid_f := 179;
        ELSIF x =- 4798 THEN
            sigmoid_f := 179;
        ELSIF x =- 4797 THEN
            sigmoid_f := 179;
        ELSIF x =- 4796 THEN
            sigmoid_f := 179;
        ELSIF x =- 4795 THEN
            sigmoid_f := 180;
        ELSIF x =- 4794 THEN
            sigmoid_f := 180;
        ELSIF x =- 4793 THEN
            sigmoid_f := 180;
        ELSIF x =- 4792 THEN
            sigmoid_f := 180;
        ELSIF x =- 4791 THEN
            sigmoid_f := 180;
        ELSIF x =- 4790 THEN
            sigmoid_f := 180;
        ELSIF x =- 4789 THEN
            sigmoid_f := 180;
        ELSIF x =- 4788 THEN
            sigmoid_f := 180;
        ELSIF x =- 4787 THEN
            sigmoid_f := 180;
        ELSIF x =- 4786 THEN
            sigmoid_f := 180;
        ELSIF x =- 4785 THEN
            sigmoid_f := 180;
        ELSIF x =- 4784 THEN
            sigmoid_f := 180;
        ELSIF x =- 4783 THEN
            sigmoid_f := 180;
        ELSIF x =- 4782 THEN
            sigmoid_f := 181;
        ELSIF x =- 4781 THEN
            sigmoid_f := 181;
        ELSIF x =- 4780 THEN
            sigmoid_f := 181;
        ELSIF x =- 4779 THEN
            sigmoid_f := 181;
        ELSIF x =- 4778 THEN
            sigmoid_f := 181;
        ELSIF x =- 4777 THEN
            sigmoid_f := 181;
        ELSIF x =- 4776 THEN
            sigmoid_f := 181;
        ELSIF x =- 4775 THEN
            sigmoid_f := 181;
        ELSIF x =- 4774 THEN
            sigmoid_f := 181;
        ELSIF x =- 4773 THEN
            sigmoid_f := 181;
        ELSIF x =- 4772 THEN
            sigmoid_f := 181;
        ELSIF x =- 4771 THEN
            sigmoid_f := 181;
        ELSIF x =- 4770 THEN
            sigmoid_f := 182;
        ELSIF x =- 4769 THEN
            sigmoid_f := 182;
        ELSIF x =- 4768 THEN
            sigmoid_f := 182;
        ELSIF x =- 4767 THEN
            sigmoid_f := 182;
        ELSIF x =- 4766 THEN
            sigmoid_f := 182;
        ELSIF x =- 4765 THEN
            sigmoid_f := 182;
        ELSIF x =- 4764 THEN
            sigmoid_f := 182;
        ELSIF x =- 4763 THEN
            sigmoid_f := 182;
        ELSIF x =- 4762 THEN
            sigmoid_f := 182;
        ELSIF x =- 4761 THEN
            sigmoid_f := 182;
        ELSIF x =- 4760 THEN
            sigmoid_f := 182;
        ELSIF x =- 4759 THEN
            sigmoid_f := 182;
        ELSIF x =- 4758 THEN
            sigmoid_f := 182;
        ELSIF x =- 4757 THEN
            sigmoid_f := 183;
        ELSIF x =- 4756 THEN
            sigmoid_f := 183;
        ELSIF x =- 4755 THEN
            sigmoid_f := 183;
        ELSIF x =- 4754 THEN
            sigmoid_f := 183;
        ELSIF x =- 4753 THEN
            sigmoid_f := 183;
        ELSIF x =- 4752 THEN
            sigmoid_f := 183;
        ELSIF x =- 4751 THEN
            sigmoid_f := 183;
        ELSIF x =- 4750 THEN
            sigmoid_f := 183;
        ELSIF x =- 4749 THEN
            sigmoid_f := 183;
        ELSIF x =- 4748 THEN
            sigmoid_f := 183;
        ELSIF x =- 4747 THEN
            sigmoid_f := 183;
        ELSIF x =- 4746 THEN
            sigmoid_f := 183;
        ELSIF x =- 4745 THEN
            sigmoid_f := 183;
        ELSIF x =- 4744 THEN
            sigmoid_f := 184;
        ELSIF x =- 4743 THEN
            sigmoid_f := 184;
        ELSIF x =- 4742 THEN
            sigmoid_f := 184;
        ELSIF x =- 4741 THEN
            sigmoid_f := 184;
        ELSIF x =- 4740 THEN
            sigmoid_f := 184;
        ELSIF x =- 4739 THEN
            sigmoid_f := 184;
        ELSIF x =- 4738 THEN
            sigmoid_f := 184;
        ELSIF x =- 4737 THEN
            sigmoid_f := 184;
        ELSIF x =- 4736 THEN
            sigmoid_f := 184;
        ELSIF x =- 4735 THEN
            sigmoid_f := 184;
        ELSIF x =- 4734 THEN
            sigmoid_f := 184;
        ELSIF x =- 4733 THEN
            sigmoid_f := 184;
        ELSIF x =- 4732 THEN
            sigmoid_f := 185;
        ELSIF x =- 4731 THEN
            sigmoid_f := 185;
        ELSIF x =- 4730 THEN
            sigmoid_f := 185;
        ELSIF x =- 4729 THEN
            sigmoid_f := 185;
        ELSIF x =- 4728 THEN
            sigmoid_f := 185;
        ELSIF x =- 4727 THEN
            sigmoid_f := 185;
        ELSIF x =- 4726 THEN
            sigmoid_f := 185;
        ELSIF x =- 4725 THEN
            sigmoid_f := 185;
        ELSIF x =- 4724 THEN
            sigmoid_f := 185;
        ELSIF x =- 4723 THEN
            sigmoid_f := 185;
        ELSIF x =- 4722 THEN
            sigmoid_f := 185;
        ELSIF x =- 4721 THEN
            sigmoid_f := 185;
        ELSIF x =- 4720 THEN
            sigmoid_f := 185;
        ELSIF x =- 4719 THEN
            sigmoid_f := 186;
        ELSIF x =- 4718 THEN
            sigmoid_f := 186;
        ELSIF x =- 4717 THEN
            sigmoid_f := 186;
        ELSIF x =- 4716 THEN
            sigmoid_f := 186;
        ELSIF x =- 4715 THEN
            sigmoid_f := 186;
        ELSIF x =- 4714 THEN
            sigmoid_f := 186;
        ELSIF x =- 4713 THEN
            sigmoid_f := 186;
        ELSIF x =- 4712 THEN
            sigmoid_f := 186;
        ELSIF x =- 4711 THEN
            sigmoid_f := 186;
        ELSIF x =- 4710 THEN
            sigmoid_f := 186;
        ELSIF x =- 4709 THEN
            sigmoid_f := 186;
        ELSIF x =- 4708 THEN
            sigmoid_f := 186;
        ELSIF x =- 4707 THEN
            sigmoid_f := 186;
        ELSIF x =- 4706 THEN
            sigmoid_f := 187;
        ELSIF x =- 4705 THEN
            sigmoid_f := 187;
        ELSIF x =- 4704 THEN
            sigmoid_f := 187;
        ELSIF x =- 4703 THEN
            sigmoid_f := 187;
        ELSIF x =- 4702 THEN
            sigmoid_f := 187;
        ELSIF x =- 4701 THEN
            sigmoid_f := 187;
        ELSIF x =- 4700 THEN
            sigmoid_f := 187;
        ELSIF x =- 4699 THEN
            sigmoid_f := 187;
        ELSIF x =- 4698 THEN
            sigmoid_f := 187;
        ELSIF x =- 4697 THEN
            sigmoid_f := 187;
        ELSIF x =- 4696 THEN
            sigmoid_f := 187;
        ELSIF x =- 4695 THEN
            sigmoid_f := 187;
        ELSIF x =- 4694 THEN
            sigmoid_f := 187;
        ELSIF x =- 4693 THEN
            sigmoid_f := 188;
        ELSIF x =- 4692 THEN
            sigmoid_f := 188;
        ELSIF x =- 4691 THEN
            sigmoid_f := 188;
        ELSIF x =- 4690 THEN
            sigmoid_f := 188;
        ELSIF x =- 4689 THEN
            sigmoid_f := 188;
        ELSIF x =- 4688 THEN
            sigmoid_f := 188;
        ELSIF x =- 4687 THEN
            sigmoid_f := 188;
        ELSIF x =- 4686 THEN
            sigmoid_f := 188;
        ELSIF x =- 4685 THEN
            sigmoid_f := 188;
        ELSIF x =- 4684 THEN
            sigmoid_f := 188;
        ELSIF x =- 4683 THEN
            sigmoid_f := 188;
        ELSIF x =- 4682 THEN
            sigmoid_f := 188;
        ELSIF x =- 4681 THEN
            sigmoid_f := 189;
        ELSIF x =- 4680 THEN
            sigmoid_f := 189;
        ELSIF x =- 4679 THEN
            sigmoid_f := 189;
        ELSIF x =- 4678 THEN
            sigmoid_f := 189;
        ELSIF x =- 4677 THEN
            sigmoid_f := 189;
        ELSIF x =- 4676 THEN
            sigmoid_f := 189;
        ELSIF x =- 4675 THEN
            sigmoid_f := 189;
        ELSIF x =- 4674 THEN
            sigmoid_f := 189;
        ELSIF x =- 4673 THEN
            sigmoid_f := 189;
        ELSIF x =- 4672 THEN
            sigmoid_f := 189;
        ELSIF x =- 4671 THEN
            sigmoid_f := 189;
        ELSIF x =- 4670 THEN
            sigmoid_f := 189;
        ELSIF x =- 4669 THEN
            sigmoid_f := 189;
        ELSIF x =- 4668 THEN
            sigmoid_f := 190;
        ELSIF x =- 4667 THEN
            sigmoid_f := 190;
        ELSIF x =- 4666 THEN
            sigmoid_f := 190;
        ELSIF x =- 4665 THEN
            sigmoid_f := 190;
        ELSIF x =- 4664 THEN
            sigmoid_f := 190;
        ELSIF x =- 4663 THEN
            sigmoid_f := 190;
        ELSIF x =- 4662 THEN
            sigmoid_f := 190;
        ELSIF x =- 4661 THEN
            sigmoid_f := 190;
        ELSIF x =- 4660 THEN
            sigmoid_f := 190;
        ELSIF x =- 4659 THEN
            sigmoid_f := 190;
        ELSIF x =- 4658 THEN
            sigmoid_f := 190;
        ELSIF x =- 4657 THEN
            sigmoid_f := 190;
        ELSIF x =- 4656 THEN
            sigmoid_f := 190;
        ELSIF x =- 4655 THEN
            sigmoid_f := 191;
        ELSIF x =- 4654 THEN
            sigmoid_f := 191;
        ELSIF x =- 4653 THEN
            sigmoid_f := 191;
        ELSIF x =- 4652 THEN
            sigmoid_f := 191;
        ELSIF x =- 4651 THEN
            sigmoid_f := 191;
        ELSIF x =- 4650 THEN
            sigmoid_f := 191;
        ELSIF x =- 4649 THEN
            sigmoid_f := 191;
        ELSIF x =- 4648 THEN
            sigmoid_f := 191;
        ELSIF x =- 4647 THEN
            sigmoid_f := 191;
        ELSIF x =- 4646 THEN
            sigmoid_f := 191;
        ELSIF x =- 4645 THEN
            sigmoid_f := 191;
        ELSIF x =- 4644 THEN
            sigmoid_f := 191;
        ELSIF x =- 4643 THEN
            sigmoid_f := 191;
        ELSIF x =- 4642 THEN
            sigmoid_f := 192;
        ELSIF x =- 4641 THEN
            sigmoid_f := 192;
        ELSIF x =- 4640 THEN
            sigmoid_f := 192;
        ELSIF x =- 4639 THEN
            sigmoid_f := 192;
        ELSIF x =- 4638 THEN
            sigmoid_f := 192;
        ELSIF x =- 4637 THEN
            sigmoid_f := 192;
        ELSIF x =- 4636 THEN
            sigmoid_f := 192;
        ELSIF x =- 4635 THEN
            sigmoid_f := 192;
        ELSIF x =- 4634 THEN
            sigmoid_f := 192;
        ELSIF x =- 4633 THEN
            sigmoid_f := 192;
        ELSIF x =- 4632 THEN
            sigmoid_f := 192;
        ELSIF x =- 4631 THEN
            sigmoid_f := 192;
        ELSIF x =- 4630 THEN
            sigmoid_f := 193;
        ELSIF x =- 4629 THEN
            sigmoid_f := 193;
        ELSIF x =- 4628 THEN
            sigmoid_f := 193;
        ELSIF x =- 4627 THEN
            sigmoid_f := 193;
        ELSIF x =- 4626 THEN
            sigmoid_f := 193;
        ELSIF x =- 4625 THEN
            sigmoid_f := 193;
        ELSIF x =- 4624 THEN
            sigmoid_f := 193;
        ELSIF x =- 4623 THEN
            sigmoid_f := 193;
        ELSIF x =- 4622 THEN
            sigmoid_f := 193;
        ELSIF x =- 4621 THEN
            sigmoid_f := 193;
        ELSIF x =- 4620 THEN
            sigmoid_f := 193;
        ELSIF x =- 4619 THEN
            sigmoid_f := 193;
        ELSIF x =- 4618 THEN
            sigmoid_f := 193;
        ELSIF x =- 4617 THEN
            sigmoid_f := 194;
        ELSIF x =- 4616 THEN
            sigmoid_f := 194;
        ELSIF x =- 4615 THEN
            sigmoid_f := 194;
        ELSIF x =- 4614 THEN
            sigmoid_f := 194;
        ELSIF x =- 4613 THEN
            sigmoid_f := 194;
        ELSIF x =- 4612 THEN
            sigmoid_f := 194;
        ELSIF x =- 4611 THEN
            sigmoid_f := 194;
        ELSIF x =- 4610 THEN
            sigmoid_f := 194;
        ELSIF x =- 4609 THEN
            sigmoid_f := 194;
        ELSIF x =- 4608 THEN
            sigmoid_f := 194;
        ELSIF x =- 4607 THEN
            sigmoid_f := 194;
        ELSIF x =- 4606 THEN
            sigmoid_f := 194;
        ELSIF x =- 4605 THEN
            sigmoid_f := 195;
        ELSIF x =- 4604 THEN
            sigmoid_f := 195;
        ELSIF x =- 4603 THEN
            sigmoid_f := 195;
        ELSIF x =- 4602 THEN
            sigmoid_f := 195;
        ELSIF x =- 4601 THEN
            sigmoid_f := 195;
        ELSIF x =- 4600 THEN
            sigmoid_f := 195;
        ELSIF x =- 4599 THEN
            sigmoid_f := 195;
        ELSIF x =- 4598 THEN
            sigmoid_f := 195;
        ELSIF x =- 4597 THEN
            sigmoid_f := 195;
        ELSIF x =- 4596 THEN
            sigmoid_f := 195;
        ELSIF x =- 4595 THEN
            sigmoid_f := 195;
        ELSIF x =- 4594 THEN
            sigmoid_f := 196;
        ELSIF x =- 4593 THEN
            sigmoid_f := 196;
        ELSIF x =- 4592 THEN
            sigmoid_f := 196;
        ELSIF x =- 4591 THEN
            sigmoid_f := 196;
        ELSIF x =- 4590 THEN
            sigmoid_f := 196;
        ELSIF x =- 4589 THEN
            sigmoid_f := 196;
        ELSIF x =- 4588 THEN
            sigmoid_f := 196;
        ELSIF x =- 4587 THEN
            sigmoid_f := 196;
        ELSIF x =- 4586 THEN
            sigmoid_f := 196;
        ELSIF x =- 4585 THEN
            sigmoid_f := 196;
        ELSIF x =- 4584 THEN
            sigmoid_f := 197;
        ELSIF x =- 4583 THEN
            sigmoid_f := 197;
        ELSIF x =- 4582 THEN
            sigmoid_f := 197;
        ELSIF x =- 4581 THEN
            sigmoid_f := 197;
        ELSIF x =- 4580 THEN
            sigmoid_f := 197;
        ELSIF x =- 4579 THEN
            sigmoid_f := 197;
        ELSIF x =- 4578 THEN
            sigmoid_f := 197;
        ELSIF x =- 4577 THEN
            sigmoid_f := 197;
        ELSIF x =- 4576 THEN
            sigmoid_f := 197;
        ELSIF x =- 4575 THEN
            sigmoid_f := 197;
        ELSIF x =- 4574 THEN
            sigmoid_f := 197;
        ELSIF x =- 4573 THEN
            sigmoid_f := 198;
        ELSIF x =- 4572 THEN
            sigmoid_f := 198;
        ELSIF x =- 4571 THEN
            sigmoid_f := 198;
        ELSIF x =- 4570 THEN
            sigmoid_f := 198;
        ELSIF x =- 4569 THEN
            sigmoid_f := 198;
        ELSIF x =- 4568 THEN
            sigmoid_f := 198;
        ELSIF x =- 4567 THEN
            sigmoid_f := 198;
        ELSIF x =- 4566 THEN
            sigmoid_f := 198;
        ELSIF x =- 4565 THEN
            sigmoid_f := 198;
        ELSIF x =- 4564 THEN
            sigmoid_f := 198;
        ELSIF x =- 4563 THEN
            sigmoid_f := 198;
        ELSIF x =- 4562 THEN
            sigmoid_f := 199;
        ELSIF x =- 4561 THEN
            sigmoid_f := 199;
        ELSIF x =- 4560 THEN
            sigmoid_f := 199;
        ELSIF x =- 4559 THEN
            sigmoid_f := 199;
        ELSIF x =- 4558 THEN
            sigmoid_f := 199;
        ELSIF x =- 4557 THEN
            sigmoid_f := 199;
        ELSIF x =- 4556 THEN
            sigmoid_f := 199;
        ELSIF x =- 4555 THEN
            sigmoid_f := 199;
        ELSIF x =- 4554 THEN
            sigmoid_f := 199;
        ELSIF x =- 4553 THEN
            sigmoid_f := 199;
        ELSIF x =- 4552 THEN
            sigmoid_f := 200;
        ELSIF x =- 4551 THEN
            sigmoid_f := 200;
        ELSIF x =- 4550 THEN
            sigmoid_f := 200;
        ELSIF x =- 4549 THEN
            sigmoid_f := 200;
        ELSIF x =- 4548 THEN
            sigmoid_f := 200;
        ELSIF x =- 4547 THEN
            sigmoid_f := 200;
        ELSIF x =- 4546 THEN
            sigmoid_f := 200;
        ELSIF x =- 4545 THEN
            sigmoid_f := 200;
        ELSIF x =- 4544 THEN
            sigmoid_f := 200;
        ELSIF x =- 4543 THEN
            sigmoid_f := 200;
        ELSIF x =- 4542 THEN
            sigmoid_f := 200;
        ELSIF x =- 4541 THEN
            sigmoid_f := 201;
        ELSIF x =- 4540 THEN
            sigmoid_f := 201;
        ELSIF x =- 4539 THEN
            sigmoid_f := 201;
        ELSIF x =- 4538 THEN
            sigmoid_f := 201;
        ELSIF x =- 4537 THEN
            sigmoid_f := 201;
        ELSIF x =- 4536 THEN
            sigmoid_f := 201;
        ELSIF x =- 4535 THEN
            sigmoid_f := 201;
        ELSIF x =- 4534 THEN
            sigmoid_f := 201;
        ELSIF x =- 4533 THEN
            sigmoid_f := 201;
        ELSIF x =- 4532 THEN
            sigmoid_f := 201;
        ELSIF x =- 4531 THEN
            sigmoid_f := 202;
        ELSIF x =- 4530 THEN
            sigmoid_f := 202;
        ELSIF x =- 4529 THEN
            sigmoid_f := 202;
        ELSIF x =- 4528 THEN
            sigmoid_f := 202;
        ELSIF x =- 4527 THEN
            sigmoid_f := 202;
        ELSIF x =- 4526 THEN
            sigmoid_f := 202;
        ELSIF x =- 4525 THEN
            sigmoid_f := 202;
        ELSIF x =- 4524 THEN
            sigmoid_f := 202;
        ELSIF x =- 4523 THEN
            sigmoid_f := 202;
        ELSIF x =- 4522 THEN
            sigmoid_f := 202;
        ELSIF x =- 4521 THEN
            sigmoid_f := 202;
        ELSIF x =- 4520 THEN
            sigmoid_f := 203;
        ELSIF x =- 4519 THEN
            sigmoid_f := 203;
        ELSIF x =- 4518 THEN
            sigmoid_f := 203;
        ELSIF x =- 4517 THEN
            sigmoid_f := 203;
        ELSIF x =- 4516 THEN
            sigmoid_f := 203;
        ELSIF x =- 4515 THEN
            sigmoid_f := 203;
        ELSIF x =- 4514 THEN
            sigmoid_f := 203;
        ELSIF x =- 4513 THEN
            sigmoid_f := 203;
        ELSIF x =- 4512 THEN
            sigmoid_f := 203;
        ELSIF x =- 4511 THEN
            sigmoid_f := 203;
        ELSIF x =- 4510 THEN
            sigmoid_f := 203;
        ELSIF x =- 4509 THEN
            sigmoid_f := 204;
        ELSIF x =- 4508 THEN
            sigmoid_f := 204;
        ELSIF x =- 4507 THEN
            sigmoid_f := 204;
        ELSIF x =- 4506 THEN
            sigmoid_f := 204;
        ELSIF x =- 4505 THEN
            sigmoid_f := 204;
        ELSIF x =- 4504 THEN
            sigmoid_f := 204;
        ELSIF x =- 4503 THEN
            sigmoid_f := 204;
        ELSIF x =- 4502 THEN
            sigmoid_f := 204;
        ELSIF x =- 4501 THEN
            sigmoid_f := 204;
        ELSIF x =- 4500 THEN
            sigmoid_f := 204;
        ELSIF x =- 4499 THEN
            sigmoid_f := 205;
        ELSIF x =- 4498 THEN
            sigmoid_f := 205;
        ELSIF x =- 4497 THEN
            sigmoid_f := 205;
        ELSIF x =- 4496 THEN
            sigmoid_f := 205;
        ELSIF x =- 4495 THEN
            sigmoid_f := 205;
        ELSIF x =- 4494 THEN
            sigmoid_f := 205;
        ELSIF x =- 4493 THEN
            sigmoid_f := 205;
        ELSIF x =- 4492 THEN
            sigmoid_f := 205;
        ELSIF x =- 4491 THEN
            sigmoid_f := 205;
        ELSIF x =- 4490 THEN
            sigmoid_f := 205;
        ELSIF x =- 4489 THEN
            sigmoid_f := 205;
        ELSIF x =- 4488 THEN
            sigmoid_f := 206;
        ELSIF x =- 4487 THEN
            sigmoid_f := 206;
        ELSIF x =- 4486 THEN
            sigmoid_f := 206;
        ELSIF x =- 4485 THEN
            sigmoid_f := 206;
        ELSIF x =- 4484 THEN
            sigmoid_f := 206;
        ELSIF x =- 4483 THEN
            sigmoid_f := 206;
        ELSIF x =- 4482 THEN
            sigmoid_f := 206;
        ELSIF x =- 4481 THEN
            sigmoid_f := 206;
        ELSIF x =- 4480 THEN
            sigmoid_f := 206;
        ELSIF x =- 4479 THEN
            sigmoid_f := 206;
        ELSIF x =- 4478 THEN
            sigmoid_f := 207;
        ELSIF x =- 4477 THEN
            sigmoid_f := 207;
        ELSIF x =- 4476 THEN
            sigmoid_f := 207;
        ELSIF x =- 4475 THEN
            sigmoid_f := 207;
        ELSIF x =- 4474 THEN
            sigmoid_f := 207;
        ELSIF x =- 4473 THEN
            sigmoid_f := 207;
        ELSIF x =- 4472 THEN
            sigmoid_f := 207;
        ELSIF x =- 4471 THEN
            sigmoid_f := 207;
        ELSIF x =- 4470 THEN
            sigmoid_f := 207;
        ELSIF x =- 4469 THEN
            sigmoid_f := 207;
        ELSIF x =- 4468 THEN
            sigmoid_f := 207;
        ELSIF x =- 4467 THEN
            sigmoid_f := 208;
        ELSIF x =- 4466 THEN
            sigmoid_f := 208;
        ELSIF x =- 4465 THEN
            sigmoid_f := 208;
        ELSIF x =- 4464 THEN
            sigmoid_f := 208;
        ELSIF x =- 4463 THEN
            sigmoid_f := 208;
        ELSIF x =- 4462 THEN
            sigmoid_f := 208;
        ELSIF x =- 4461 THEN
            sigmoid_f := 208;
        ELSIF x =- 4460 THEN
            sigmoid_f := 208;
        ELSIF x =- 4459 THEN
            sigmoid_f := 208;
        ELSIF x =- 4458 THEN
            sigmoid_f := 208;
        ELSIF x =- 4457 THEN
            sigmoid_f := 208;
        ELSIF x =- 4456 THEN
            sigmoid_f := 209;
        ELSIF x =- 4455 THEN
            sigmoid_f := 209;
        ELSIF x =- 4454 THEN
            sigmoid_f := 209;
        ELSIF x =- 4453 THEN
            sigmoid_f := 209;
        ELSIF x =- 4452 THEN
            sigmoid_f := 209;
        ELSIF x =- 4451 THEN
            sigmoid_f := 209;
        ELSIF x =- 4450 THEN
            sigmoid_f := 209;
        ELSIF x =- 4449 THEN
            sigmoid_f := 209;
        ELSIF x =- 4448 THEN
            sigmoid_f := 209;
        ELSIF x =- 4447 THEN
            sigmoid_f := 209;
        ELSIF x =- 4446 THEN
            sigmoid_f := 210;
        ELSIF x =- 4445 THEN
            sigmoid_f := 210;
        ELSIF x =- 4444 THEN
            sigmoid_f := 210;
        ELSIF x =- 4443 THEN
            sigmoid_f := 210;
        ELSIF x =- 4442 THEN
            sigmoid_f := 210;
        ELSIF x =- 4441 THEN
            sigmoid_f := 210;
        ELSIF x =- 4440 THEN
            sigmoid_f := 210;
        ELSIF x =- 4439 THEN
            sigmoid_f := 210;
        ELSIF x =- 4438 THEN
            sigmoid_f := 210;
        ELSIF x =- 4437 THEN
            sigmoid_f := 210;
        ELSIF x =- 4436 THEN
            sigmoid_f := 210;
        ELSIF x =- 4435 THEN
            sigmoid_f := 211;
        ELSIF x =- 4434 THEN
            sigmoid_f := 211;
        ELSIF x =- 4433 THEN
            sigmoid_f := 211;
        ELSIF x =- 4432 THEN
            sigmoid_f := 211;
        ELSIF x =- 4431 THEN
            sigmoid_f := 211;
        ELSIF x =- 4430 THEN
            sigmoid_f := 211;
        ELSIF x =- 4429 THEN
            sigmoid_f := 211;
        ELSIF x =- 4428 THEN
            sigmoid_f := 211;
        ELSIF x =- 4427 THEN
            sigmoid_f := 211;
        ELSIF x =- 4426 THEN
            sigmoid_f := 211;
        ELSIF x =- 4425 THEN
            sigmoid_f := 211;
        ELSIF x =- 4424 THEN
            sigmoid_f := 212;
        ELSIF x =- 4423 THEN
            sigmoid_f := 212;
        ELSIF x =- 4422 THEN
            sigmoid_f := 212;
        ELSIF x =- 4421 THEN
            sigmoid_f := 212;
        ELSIF x =- 4420 THEN
            sigmoid_f := 212;
        ELSIF x =- 4419 THEN
            sigmoid_f := 212;
        ELSIF x =- 4418 THEN
            sigmoid_f := 212;
        ELSIF x =- 4417 THEN
            sigmoid_f := 212;
        ELSIF x =- 4416 THEN
            sigmoid_f := 212;
        ELSIF x =- 4415 THEN
            sigmoid_f := 212;
        ELSIF x =- 4414 THEN
            sigmoid_f := 213;
        ELSIF x =- 4413 THEN
            sigmoid_f := 213;
        ELSIF x =- 4412 THEN
            sigmoid_f := 213;
        ELSIF x =- 4411 THEN
            sigmoid_f := 213;
        ELSIF x =- 4410 THEN
            sigmoid_f := 213;
        ELSIF x =- 4409 THEN
            sigmoid_f := 213;
        ELSIF x =- 4408 THEN
            sigmoid_f := 213;
        ELSIF x =- 4407 THEN
            sigmoid_f := 213;
        ELSIF x =- 4406 THEN
            sigmoid_f := 213;
        ELSIF x =- 4405 THEN
            sigmoid_f := 213;
        ELSIF x =- 4404 THEN
            sigmoid_f := 213;
        ELSIF x =- 4403 THEN
            sigmoid_f := 214;
        ELSIF x =- 4402 THEN
            sigmoid_f := 214;
        ELSIF x =- 4401 THEN
            sigmoid_f := 214;
        ELSIF x =- 4400 THEN
            sigmoid_f := 214;
        ELSIF x =- 4399 THEN
            sigmoid_f := 214;
        ELSIF x =- 4398 THEN
            sigmoid_f := 214;
        ELSIF x =- 4397 THEN
            sigmoid_f := 214;
        ELSIF x =- 4396 THEN
            sigmoid_f := 214;
        ELSIF x =- 4395 THEN
            sigmoid_f := 214;
        ELSIF x =- 4394 THEN
            sigmoid_f := 214;
        ELSIF x =- 4393 THEN
            sigmoid_f := 215;
        ELSIF x =- 4392 THEN
            sigmoid_f := 215;
        ELSIF x =- 4391 THEN
            sigmoid_f := 215;
        ELSIF x =- 4390 THEN
            sigmoid_f := 215;
        ELSIF x =- 4389 THEN
            sigmoid_f := 215;
        ELSIF x =- 4388 THEN
            sigmoid_f := 215;
        ELSIF x =- 4387 THEN
            sigmoid_f := 215;
        ELSIF x =- 4386 THEN
            sigmoid_f := 215;
        ELSIF x =- 4385 THEN
            sigmoid_f := 215;
        ELSIF x =- 4384 THEN
            sigmoid_f := 215;
        ELSIF x =- 4383 THEN
            sigmoid_f := 215;
        ELSIF x =- 4382 THEN
            sigmoid_f := 216;
        ELSIF x =- 4381 THEN
            sigmoid_f := 216;
        ELSIF x =- 4380 THEN
            sigmoid_f := 216;
        ELSIF x =- 4379 THEN
            sigmoid_f := 216;
        ELSIF x =- 4378 THEN
            sigmoid_f := 216;
        ELSIF x =- 4377 THEN
            sigmoid_f := 216;
        ELSIF x =- 4376 THEN
            sigmoid_f := 216;
        ELSIF x =- 4375 THEN
            sigmoid_f := 216;
        ELSIF x =- 4374 THEN
            sigmoid_f := 216;
        ELSIF x =- 4373 THEN
            sigmoid_f := 216;
        ELSIF x =- 4372 THEN
            sigmoid_f := 216;
        ELSIF x =- 4371 THEN
            sigmoid_f := 217;
        ELSIF x =- 4370 THEN
            sigmoid_f := 217;
        ELSIF x =- 4369 THEN
            sigmoid_f := 217;
        ELSIF x =- 4368 THEN
            sigmoid_f := 217;
        ELSIF x =- 4367 THEN
            sigmoid_f := 217;
        ELSIF x =- 4366 THEN
            sigmoid_f := 217;
        ELSIF x =- 4365 THEN
            sigmoid_f := 217;
        ELSIF x =- 4364 THEN
            sigmoid_f := 217;
        ELSIF x =- 4363 THEN
            sigmoid_f := 217;
        ELSIF x =- 4362 THEN
            sigmoid_f := 217;
        ELSIF x =- 4361 THEN
            sigmoid_f := 218;
        ELSIF x =- 4360 THEN
            sigmoid_f := 218;
        ELSIF x =- 4359 THEN
            sigmoid_f := 218;
        ELSIF x =- 4358 THEN
            sigmoid_f := 218;
        ELSIF x =- 4357 THEN
            sigmoid_f := 218;
        ELSIF x =- 4356 THEN
            sigmoid_f := 218;
        ELSIF x =- 4355 THEN
            sigmoid_f := 218;
        ELSIF x =- 4354 THEN
            sigmoid_f := 218;
        ELSIF x =- 4353 THEN
            sigmoid_f := 218;
        ELSIF x =- 4352 THEN
            sigmoid_f := 218;
        ELSIF x =- 4351 THEN
            sigmoid_f := 218;
        ELSIF x =- 4350 THEN
            sigmoid_f := 219;
        ELSIF x =- 4349 THEN
            sigmoid_f := 219;
        ELSIF x =- 4348 THEN
            sigmoid_f := 219;
        ELSIF x =- 4347 THEN
            sigmoid_f := 219;
        ELSIF x =- 4346 THEN
            sigmoid_f := 219;
        ELSIF x =- 4345 THEN
            sigmoid_f := 219;
        ELSIF x =- 4344 THEN
            sigmoid_f := 219;
        ELSIF x =- 4343 THEN
            sigmoid_f := 219;
        ELSIF x =- 4342 THEN
            sigmoid_f := 219;
        ELSIF x =- 4341 THEN
            sigmoid_f := 219;
        ELSIF x =- 4340 THEN
            sigmoid_f := 220;
        ELSIF x =- 4339 THEN
            sigmoid_f := 220;
        ELSIF x =- 4338 THEN
            sigmoid_f := 220;
        ELSIF x =- 4337 THEN
            sigmoid_f := 220;
        ELSIF x =- 4336 THEN
            sigmoid_f := 220;
        ELSIF x =- 4335 THEN
            sigmoid_f := 220;
        ELSIF x =- 4334 THEN
            sigmoid_f := 220;
        ELSIF x =- 4333 THEN
            sigmoid_f := 220;
        ELSIF x =- 4332 THEN
            sigmoid_f := 220;
        ELSIF x =- 4331 THEN
            sigmoid_f := 220;
        ELSIF x =- 4330 THEN
            sigmoid_f := 220;
        ELSIF x =- 4329 THEN
            sigmoid_f := 221;
        ELSIF x =- 4328 THEN
            sigmoid_f := 221;
        ELSIF x =- 4327 THEN
            sigmoid_f := 221;
        ELSIF x =- 4326 THEN
            sigmoid_f := 221;
        ELSIF x =- 4325 THEN
            sigmoid_f := 221;
        ELSIF x =- 4324 THEN
            sigmoid_f := 221;
        ELSIF x =- 4323 THEN
            sigmoid_f := 221;
        ELSIF x =- 4322 THEN
            sigmoid_f := 221;
        ELSIF x =- 4321 THEN
            sigmoid_f := 221;
        ELSIF x =- 4320 THEN
            sigmoid_f := 221;
        ELSIF x =- 4319 THEN
            sigmoid_f := 221;
        ELSIF x =- 4318 THEN
            sigmoid_f := 222;
        ELSIF x =- 4317 THEN
            sigmoid_f := 222;
        ELSIF x =- 4316 THEN
            sigmoid_f := 222;
        ELSIF x =- 4315 THEN
            sigmoid_f := 222;
        ELSIF x =- 4314 THEN
            sigmoid_f := 222;
        ELSIF x =- 4313 THEN
            sigmoid_f := 222;
        ELSIF x =- 4312 THEN
            sigmoid_f := 222;
        ELSIF x =- 4311 THEN
            sigmoid_f := 222;
        ELSIF x =- 4310 THEN
            sigmoid_f := 222;
        ELSIF x =- 4309 THEN
            sigmoid_f := 222;
        ELSIF x =- 4308 THEN
            sigmoid_f := 223;
        ELSIF x =- 4307 THEN
            sigmoid_f := 223;
        ELSIF x =- 4306 THEN
            sigmoid_f := 223;
        ELSIF x =- 4305 THEN
            sigmoid_f := 223;
        ELSIF x =- 4304 THEN
            sigmoid_f := 223;
        ELSIF x =- 4303 THEN
            sigmoid_f := 223;
        ELSIF x =- 4302 THEN
            sigmoid_f := 223;
        ELSIF x =- 4301 THEN
            sigmoid_f := 223;
        ELSIF x =- 4300 THEN
            sigmoid_f := 223;
        ELSIF x =- 4299 THEN
            sigmoid_f := 223;
        ELSIF x =- 4298 THEN
            sigmoid_f := 223;
        ELSIF x =- 4297 THEN
            sigmoid_f := 224;
        ELSIF x =- 4296 THEN
            sigmoid_f := 224;
        ELSIF x =- 4295 THEN
            sigmoid_f := 224;
        ELSIF x =- 4294 THEN
            sigmoid_f := 224;
        ELSIF x =- 4293 THEN
            sigmoid_f := 224;
        ELSIF x =- 4292 THEN
            sigmoid_f := 224;
        ELSIF x =- 4291 THEN
            sigmoid_f := 224;
        ELSIF x =- 4290 THEN
            sigmoid_f := 224;
        ELSIF x =- 4289 THEN
            sigmoid_f := 224;
        ELSIF x =- 4288 THEN
            sigmoid_f := 224;
        ELSIF x =- 4287 THEN
            sigmoid_f := 225;
        ELSIF x =- 4286 THEN
            sigmoid_f := 225;
        ELSIF x =- 4285 THEN
            sigmoid_f := 225;
        ELSIF x =- 4284 THEN
            sigmoid_f := 225;
        ELSIF x =- 4283 THEN
            sigmoid_f := 225;
        ELSIF x =- 4282 THEN
            sigmoid_f := 225;
        ELSIF x =- 4281 THEN
            sigmoid_f := 225;
        ELSIF x =- 4280 THEN
            sigmoid_f := 225;
        ELSIF x =- 4279 THEN
            sigmoid_f := 225;
        ELSIF x =- 4278 THEN
            sigmoid_f := 225;
        ELSIF x =- 4277 THEN
            sigmoid_f := 225;
        ELSIF x =- 4276 THEN
            sigmoid_f := 226;
        ELSIF x =- 4275 THEN
            sigmoid_f := 226;
        ELSIF x =- 4274 THEN
            sigmoid_f := 226;
        ELSIF x =- 4273 THEN
            sigmoid_f := 226;
        ELSIF x =- 4272 THEN
            sigmoid_f := 226;
        ELSIF x =- 4271 THEN
            sigmoid_f := 226;
        ELSIF x =- 4270 THEN
            sigmoid_f := 226;
        ELSIF x =- 4269 THEN
            sigmoid_f := 226;
        ELSIF x =- 4268 THEN
            sigmoid_f := 226;
        ELSIF x =- 4267 THEN
            sigmoid_f := 226;
        ELSIF x =- 4266 THEN
            sigmoid_f := 226;
        ELSIF x =- 4265 THEN
            sigmoid_f := 227;
        ELSIF x =- 4264 THEN
            sigmoid_f := 227;
        ELSIF x =- 4263 THEN
            sigmoid_f := 227;
        ELSIF x =- 4262 THEN
            sigmoid_f := 227;
        ELSIF x =- 4261 THEN
            sigmoid_f := 227;
        ELSIF x =- 4260 THEN
            sigmoid_f := 227;
        ELSIF x =- 4259 THEN
            sigmoid_f := 227;
        ELSIF x =- 4258 THEN
            sigmoid_f := 227;
        ELSIF x =- 4257 THEN
            sigmoid_f := 227;
        ELSIF x =- 4256 THEN
            sigmoid_f := 227;
        ELSIF x =- 4255 THEN
            sigmoid_f := 228;
        ELSIF x =- 4254 THEN
            sigmoid_f := 228;
        ELSIF x =- 4253 THEN
            sigmoid_f := 228;
        ELSIF x =- 4252 THEN
            sigmoid_f := 228;
        ELSIF x =- 4251 THEN
            sigmoid_f := 228;
        ELSIF x =- 4250 THEN
            sigmoid_f := 228;
        ELSIF x =- 4249 THEN
            sigmoid_f := 228;
        ELSIF x =- 4248 THEN
            sigmoid_f := 228;
        ELSIF x =- 4247 THEN
            sigmoid_f := 228;
        ELSIF x =- 4246 THEN
            sigmoid_f := 228;
        ELSIF x =- 4245 THEN
            sigmoid_f := 228;
        ELSIF x =- 4244 THEN
            sigmoid_f := 229;
        ELSIF x =- 4243 THEN
            sigmoid_f := 229;
        ELSIF x =- 4242 THEN
            sigmoid_f := 229;
        ELSIF x =- 4241 THEN
            sigmoid_f := 229;
        ELSIF x =- 4240 THEN
            sigmoid_f := 229;
        ELSIF x =- 4239 THEN
            sigmoid_f := 229;
        ELSIF x =- 4238 THEN
            sigmoid_f := 229;
        ELSIF x =- 4237 THEN
            sigmoid_f := 229;
        ELSIF x =- 4236 THEN
            sigmoid_f := 229;
        ELSIF x =- 4235 THEN
            sigmoid_f := 229;
        ELSIF x =- 4234 THEN
            sigmoid_f := 229;
        ELSIF x =- 4233 THEN
            sigmoid_f := 230;
        ELSIF x =- 4232 THEN
            sigmoid_f := 230;
        ELSIF x =- 4231 THEN
            sigmoid_f := 230;
        ELSIF x =- 4230 THEN
            sigmoid_f := 230;
        ELSIF x =- 4229 THEN
            sigmoid_f := 230;
        ELSIF x =- 4228 THEN
            sigmoid_f := 230;
        ELSIF x =- 4227 THEN
            sigmoid_f := 230;
        ELSIF x =- 4226 THEN
            sigmoid_f := 230;
        ELSIF x =- 4225 THEN
            sigmoid_f := 230;
        ELSIF x =- 4224 THEN
            sigmoid_f := 230;
        ELSIF x =- 4223 THEN
            sigmoid_f := 231;
        ELSIF x =- 4222 THEN
            sigmoid_f := 231;
        ELSIF x =- 4221 THEN
            sigmoid_f := 231;
        ELSIF x =- 4220 THEN
            sigmoid_f := 231;
        ELSIF x =- 4219 THEN
            sigmoid_f := 231;
        ELSIF x =- 4218 THEN
            sigmoid_f := 231;
        ELSIF x =- 4217 THEN
            sigmoid_f := 231;
        ELSIF x =- 4216 THEN
            sigmoid_f := 231;
        ELSIF x =- 4215 THEN
            sigmoid_f := 231;
        ELSIF x =- 4214 THEN
            sigmoid_f := 231;
        ELSIF x =- 4213 THEN
            sigmoid_f := 231;
        ELSIF x =- 4212 THEN
            sigmoid_f := 232;
        ELSIF x =- 4211 THEN
            sigmoid_f := 232;
        ELSIF x =- 4210 THEN
            sigmoid_f := 232;
        ELSIF x =- 4209 THEN
            sigmoid_f := 232;
        ELSIF x =- 4208 THEN
            sigmoid_f := 232;
        ELSIF x =- 4207 THEN
            sigmoid_f := 232;
        ELSIF x =- 4206 THEN
            sigmoid_f := 232;
        ELSIF x =- 4205 THEN
            sigmoid_f := 232;
        ELSIF x =- 4204 THEN
            sigmoid_f := 232;
        ELSIF x =- 4203 THEN
            sigmoid_f := 232;
        ELSIF x =- 4202 THEN
            sigmoid_f := 233;
        ELSIF x =- 4201 THEN
            sigmoid_f := 233;
        ELSIF x =- 4200 THEN
            sigmoid_f := 233;
        ELSIF x =- 4199 THEN
            sigmoid_f := 233;
        ELSIF x =- 4198 THEN
            sigmoid_f := 233;
        ELSIF x =- 4197 THEN
            sigmoid_f := 233;
        ELSIF x =- 4196 THEN
            sigmoid_f := 233;
        ELSIF x =- 4195 THEN
            sigmoid_f := 233;
        ELSIF x =- 4194 THEN
            sigmoid_f := 233;
        ELSIF x =- 4193 THEN
            sigmoid_f := 233;
        ELSIF x =- 4192 THEN
            sigmoid_f := 233;
        ELSIF x =- 4191 THEN
            sigmoid_f := 234;
        ELSIF x =- 4190 THEN
            sigmoid_f := 234;
        ELSIF x =- 4189 THEN
            sigmoid_f := 234;
        ELSIF x =- 4188 THEN
            sigmoid_f := 234;
        ELSIF x =- 4187 THEN
            sigmoid_f := 234;
        ELSIF x =- 4186 THEN
            sigmoid_f := 234;
        ELSIF x =- 4185 THEN
            sigmoid_f := 234;
        ELSIF x =- 4184 THEN
            sigmoid_f := 234;
        ELSIF x =- 4183 THEN
            sigmoid_f := 234;
        ELSIF x =- 4182 THEN
            sigmoid_f := 234;
        ELSIF x =- 4181 THEN
            sigmoid_f := 234;
        ELSIF x =- 4180 THEN
            sigmoid_f := 235;
        ELSIF x =- 4179 THEN
            sigmoid_f := 235;
        ELSIF x =- 4178 THEN
            sigmoid_f := 235;
        ELSIF x =- 4177 THEN
            sigmoid_f := 235;
        ELSIF x =- 4176 THEN
            sigmoid_f := 235;
        ELSIF x =- 4175 THEN
            sigmoid_f := 235;
        ELSIF x =- 4174 THEN
            sigmoid_f := 235;
        ELSIF x =- 4173 THEN
            sigmoid_f := 235;
        ELSIF x =- 4172 THEN
            sigmoid_f := 235;
        ELSIF x =- 4171 THEN
            sigmoid_f := 235;
        ELSIF x =- 4170 THEN
            sigmoid_f := 236;
        ELSIF x =- 4169 THEN
            sigmoid_f := 236;
        ELSIF x =- 4168 THEN
            sigmoid_f := 236;
        ELSIF x =- 4167 THEN
            sigmoid_f := 236;
        ELSIF x =- 4166 THEN
            sigmoid_f := 236;
        ELSIF x =- 4165 THEN
            sigmoid_f := 236;
        ELSIF x =- 4164 THEN
            sigmoid_f := 236;
        ELSIF x =- 4163 THEN
            sigmoid_f := 236;
        ELSIF x =- 4162 THEN
            sigmoid_f := 236;
        ELSIF x =- 4161 THEN
            sigmoid_f := 236;
        ELSIF x =- 4160 THEN
            sigmoid_f := 236;
        ELSIF x =- 4159 THEN
            sigmoid_f := 237;
        ELSIF x =- 4158 THEN
            sigmoid_f := 237;
        ELSIF x =- 4157 THEN
            sigmoid_f := 237;
        ELSIF x =- 4156 THEN
            sigmoid_f := 237;
        ELSIF x =- 4155 THEN
            sigmoid_f := 237;
        ELSIF x =- 4154 THEN
            sigmoid_f := 237;
        ELSIF x =- 4153 THEN
            sigmoid_f := 237;
        ELSIF x =- 4152 THEN
            sigmoid_f := 237;
        ELSIF x =- 4151 THEN
            sigmoid_f := 237;
        ELSIF x =- 4150 THEN
            sigmoid_f := 237;
        ELSIF x =- 4149 THEN
            sigmoid_f := 238;
        ELSIF x =- 4148 THEN
            sigmoid_f := 238;
        ELSIF x =- 4147 THEN
            sigmoid_f := 238;
        ELSIF x =- 4146 THEN
            sigmoid_f := 238;
        ELSIF x =- 4145 THEN
            sigmoid_f := 238;
        ELSIF x =- 4144 THEN
            sigmoid_f := 238;
        ELSIF x =- 4143 THEN
            sigmoid_f := 238;
        ELSIF x =- 4142 THEN
            sigmoid_f := 238;
        ELSIF x =- 4141 THEN
            sigmoid_f := 238;
        ELSIF x =- 4140 THEN
            sigmoid_f := 238;
        ELSIF x =- 4139 THEN
            sigmoid_f := 238;
        ELSIF x =- 4138 THEN
            sigmoid_f := 239;
        ELSIF x =- 4137 THEN
            sigmoid_f := 239;
        ELSIF x =- 4136 THEN
            sigmoid_f := 239;
        ELSIF x =- 4135 THEN
            sigmoid_f := 239;
        ELSIF x =- 4134 THEN
            sigmoid_f := 239;
        ELSIF x =- 4133 THEN
            sigmoid_f := 239;
        ELSIF x =- 4132 THEN
            sigmoid_f := 239;
        ELSIF x =- 4131 THEN
            sigmoid_f := 239;
        ELSIF x =- 4130 THEN
            sigmoid_f := 239;
        ELSIF x =- 4129 THEN
            sigmoid_f := 239;
        ELSIF x =- 4128 THEN
            sigmoid_f := 239;
        ELSIF x =- 4127 THEN
            sigmoid_f := 240;
        ELSIF x =- 4126 THEN
            sigmoid_f := 240;
        ELSIF x =- 4125 THEN
            sigmoid_f := 240;
        ELSIF x =- 4124 THEN
            sigmoid_f := 240;
        ELSIF x =- 4123 THEN
            sigmoid_f := 240;
        ELSIF x =- 4122 THEN
            sigmoid_f := 240;
        ELSIF x =- 4121 THEN
            sigmoid_f := 240;
        ELSIF x =- 4120 THEN
            sigmoid_f := 240;
        ELSIF x =- 4119 THEN
            sigmoid_f := 240;
        ELSIF x =- 4118 THEN
            sigmoid_f := 240;
        ELSIF x =- 4117 THEN
            sigmoid_f := 241;
        ELSIF x =- 4116 THEN
            sigmoid_f := 241;
        ELSIF x =- 4115 THEN
            sigmoid_f := 241;
        ELSIF x =- 4114 THEN
            sigmoid_f := 241;
        ELSIF x =- 4113 THEN
            sigmoid_f := 241;
        ELSIF x =- 4112 THEN
            sigmoid_f := 241;
        ELSIF x =- 4111 THEN
            sigmoid_f := 241;
        ELSIF x =- 4110 THEN
            sigmoid_f := 241;
        ELSIF x =- 4109 THEN
            sigmoid_f := 241;
        ELSIF x =- 4108 THEN
            sigmoid_f := 241;
        ELSIF x =- 4107 THEN
            sigmoid_f := 241;
        ELSIF x =- 4106 THEN
            sigmoid_f := 242;
        ELSIF x =- 4105 THEN
            sigmoid_f := 242;
        ELSIF x =- 4104 THEN
            sigmoid_f := 242;
        ELSIF x =- 4103 THEN
            sigmoid_f := 242;
        ELSIF x =- 4102 THEN
            sigmoid_f := 242;
        ELSIF x =- 4101 THEN
            sigmoid_f := 242;
        ELSIF x =- 4100 THEN
            sigmoid_f := 242;
        ELSIF x =- 4099 THEN
            sigmoid_f := 242;
        ELSIF x =- 4098 THEN
            sigmoid_f := 242;
        ELSIF x =- 4097 THEN
            sigmoid_f := 242;
        ELSIF x =- 4096 THEN
            sigmoid_f := 243;
        ELSIF x =- 4095 THEN
            sigmoid_f := 243;
        ELSIF x =- 4094 THEN
            sigmoid_f := 243;
        ELSIF x =- 4093 THEN
            sigmoid_f := 243;
        ELSIF x =- 4092 THEN
            sigmoid_f := 243;
        ELSIF x =- 4091 THEN
            sigmoid_f := 243;
        ELSIF x =- 4090 THEN
            sigmoid_f := 243;
        ELSIF x =- 4089 THEN
            sigmoid_f := 243;
        ELSIF x =- 4088 THEN
            sigmoid_f := 243;
        ELSIF x =- 4087 THEN
            sigmoid_f := 244;
        ELSIF x =- 4086 THEN
            sigmoid_f := 244;
        ELSIF x =- 4085 THEN
            sigmoid_f := 244;
        ELSIF x =- 4084 THEN
            sigmoid_f := 244;
        ELSIF x =- 4083 THEN
            sigmoid_f := 244;
        ELSIF x =- 4082 THEN
            sigmoid_f := 244;
        ELSIF x =- 4081 THEN
            sigmoid_f := 244;
        ELSIF x =- 4080 THEN
            sigmoid_f := 244;
        ELSIF x =- 4079 THEN
            sigmoid_f := 244;
        ELSIF x =- 4078 THEN
            sigmoid_f := 245;
        ELSIF x =- 4077 THEN
            sigmoid_f := 245;
        ELSIF x =- 4076 THEN
            sigmoid_f := 245;
        ELSIF x =- 4075 THEN
            sigmoid_f := 245;
        ELSIF x =- 4074 THEN
            sigmoid_f := 245;
        ELSIF x =- 4073 THEN
            sigmoid_f := 245;
        ELSIF x =- 4072 THEN
            sigmoid_f := 245;
        ELSIF x =- 4071 THEN
            sigmoid_f := 245;
        ELSIF x =- 4070 THEN
            sigmoid_f := 246;
        ELSIF x =- 4069 THEN
            sigmoid_f := 246;
        ELSIF x =- 4068 THEN
            sigmoid_f := 246;
        ELSIF x =- 4067 THEN
            sigmoid_f := 246;
        ELSIF x =- 4066 THEN
            sigmoid_f := 246;
        ELSIF x =- 4065 THEN
            sigmoid_f := 246;
        ELSIF x =- 4064 THEN
            sigmoid_f := 246;
        ELSIF x =- 4063 THEN
            sigmoid_f := 246;
        ELSIF x =- 4062 THEN
            sigmoid_f := 246;
        ELSIF x =- 4061 THEN
            sigmoid_f := 247;
        ELSIF x =- 4060 THEN
            sigmoid_f := 247;
        ELSIF x =- 4059 THEN
            sigmoid_f := 247;
        ELSIF x =- 4058 THEN
            sigmoid_f := 247;
        ELSIF x =- 4057 THEN
            sigmoid_f := 247;
        ELSIF x =- 4056 THEN
            sigmoid_f := 247;
        ELSIF x =- 4055 THEN
            sigmoid_f := 247;
        ELSIF x =- 4054 THEN
            sigmoid_f := 247;
        ELSIF x =- 4053 THEN
            sigmoid_f := 247;
        ELSIF x =- 4052 THEN
            sigmoid_f := 248;
        ELSIF x =- 4051 THEN
            sigmoid_f := 248;
        ELSIF x =- 4050 THEN
            sigmoid_f := 248;
        ELSIF x =- 4049 THEN
            sigmoid_f := 248;
        ELSIF x =- 4048 THEN
            sigmoid_f := 248;
        ELSIF x =- 4047 THEN
            sigmoid_f := 248;
        ELSIF x =- 4046 THEN
            sigmoid_f := 248;
        ELSIF x =- 4045 THEN
            sigmoid_f := 248;
        ELSIF x =- 4044 THEN
            sigmoid_f := 249;
        ELSIF x =- 4043 THEN
            sigmoid_f := 249;
        ELSIF x =- 4042 THEN
            sigmoid_f := 249;
        ELSIF x =- 4041 THEN
            sigmoid_f := 249;
        ELSIF x =- 4040 THEN
            sigmoid_f := 249;
        ELSIF x =- 4039 THEN
            sigmoid_f := 249;
        ELSIF x =- 4038 THEN
            sigmoid_f := 249;
        ELSIF x =- 4037 THEN
            sigmoid_f := 249;
        ELSIF x =- 4036 THEN
            sigmoid_f := 249;
        ELSIF x =- 4035 THEN
            sigmoid_f := 250;
        ELSIF x =- 4034 THEN
            sigmoid_f := 250;
        ELSIF x =- 4033 THEN
            sigmoid_f := 250;
        ELSIF x =- 4032 THEN
            sigmoid_f := 250;
        ELSIF x =- 4031 THEN
            sigmoid_f := 250;
        ELSIF x =- 4030 THEN
            sigmoid_f := 250;
        ELSIF x =- 4029 THEN
            sigmoid_f := 250;
        ELSIF x =- 4028 THEN
            sigmoid_f := 250;
        ELSIF x =- 4027 THEN
            sigmoid_f := 251;
        ELSIF x =- 4026 THEN
            sigmoid_f := 251;
        ELSIF x =- 4025 THEN
            sigmoid_f := 251;
        ELSIF x =- 4024 THEN
            sigmoid_f := 251;
        ELSIF x =- 4023 THEN
            sigmoid_f := 251;
        ELSIF x =- 4022 THEN
            sigmoid_f := 251;
        ELSIF x =- 4021 THEN
            sigmoid_f := 251;
        ELSIF x =- 4020 THEN
            sigmoid_f := 251;
        ELSIF x =- 4019 THEN
            sigmoid_f := 251;
        ELSIF x =- 4018 THEN
            sigmoid_f := 252;
        ELSIF x =- 4017 THEN
            sigmoid_f := 252;
        ELSIF x =- 4016 THEN
            sigmoid_f := 252;
        ELSIF x =- 4015 THEN
            sigmoid_f := 252;
        ELSIF x =- 4014 THEN
            sigmoid_f := 252;
        ELSIF x =- 4013 THEN
            sigmoid_f := 252;
        ELSIF x =- 4012 THEN
            sigmoid_f := 252;
        ELSIF x =- 4011 THEN
            sigmoid_f := 252;
        ELSIF x =- 4010 THEN
            sigmoid_f := 252;
        ELSIF x =- 4009 THEN
            sigmoid_f := 253;
        ELSIF x =- 4008 THEN
            sigmoid_f := 253;
        ELSIF x =- 4007 THEN
            sigmoid_f := 253;
        ELSIF x =- 4006 THEN
            sigmoid_f := 253;
        ELSIF x =- 4005 THEN
            sigmoid_f := 253;
        ELSIF x =- 4004 THEN
            sigmoid_f := 253;
        ELSIF x =- 4003 THEN
            sigmoid_f := 253;
        ELSIF x =- 4002 THEN
            sigmoid_f := 253;
        ELSIF x =- 4001 THEN
            sigmoid_f := 254;
        ELSIF x =- 4000 THEN
            sigmoid_f := 254;
        ELSIF x =- 3999 THEN
            sigmoid_f := 254;
        ELSIF x =- 3998 THEN
            sigmoid_f := 254;
        ELSIF x =- 3997 THEN
            sigmoid_f := 254;
        ELSIF x =- 3996 THEN
            sigmoid_f := 254;
        ELSIF x =- 3995 THEN
            sigmoid_f := 254;
        ELSIF x =- 3994 THEN
            sigmoid_f := 254;
        ELSIF x =- 3993 THEN
            sigmoid_f := 254;
        ELSIF x =- 3992 THEN
            sigmoid_f := 255;
        ELSIF x =- 3991 THEN
            sigmoid_f := 255;
        ELSIF x =- 3990 THEN
            sigmoid_f := 255;
        ELSIF x =- 3989 THEN
            sigmoid_f := 255;
        ELSIF x =- 3988 THEN
            sigmoid_f := 255;
        ELSIF x =- 3987 THEN
            sigmoid_f := 255;
        ELSIF x =- 3986 THEN
            sigmoid_f := 255;
        ELSIF x =- 3985 THEN
            sigmoid_f := 255;
        ELSIF x =- 3984 THEN
            sigmoid_f := 256;
        ELSIF x =- 3983 THEN
            sigmoid_f := 256;
        ELSIF x =- 3982 THEN
            sigmoid_f := 256;
        ELSIF x =- 3981 THEN
            sigmoid_f := 256;
        ELSIF x =- 3980 THEN
            sigmoid_f := 256;
        ELSIF x =- 3979 THEN
            sigmoid_f := 256;
        ELSIF x =- 3978 THEN
            sigmoid_f := 256;
        ELSIF x =- 3977 THEN
            sigmoid_f := 256;
        ELSIF x =- 3976 THEN
            sigmoid_f := 256;
        ELSIF x =- 3975 THEN
            sigmoid_f := 257;
        ELSIF x =- 3974 THEN
            sigmoid_f := 257;
        ELSIF x =- 3973 THEN
            sigmoid_f := 257;
        ELSIF x =- 3972 THEN
            sigmoid_f := 257;
        ELSIF x =- 3971 THEN
            sigmoid_f := 257;
        ELSIF x =- 3970 THEN
            sigmoid_f := 257;
        ELSIF x =- 3969 THEN
            sigmoid_f := 257;
        ELSIF x =- 3968 THEN
            sigmoid_f := 257;
        ELSIF x =- 3967 THEN
            sigmoid_f := 257;
        ELSIF x =- 3966 THEN
            sigmoid_f := 258;
        ELSIF x =- 3965 THEN
            sigmoid_f := 258;
        ELSIF x =- 3964 THEN
            sigmoid_f := 258;
        ELSIF x =- 3963 THEN
            sigmoid_f := 258;
        ELSIF x =- 3962 THEN
            sigmoid_f := 258;
        ELSIF x =- 3961 THEN
            sigmoid_f := 258;
        ELSIF x =- 3960 THEN
            sigmoid_f := 258;
        ELSIF x =- 3959 THEN
            sigmoid_f := 258;
        ELSIF x =- 3958 THEN
            sigmoid_f := 259;
        ELSIF x =- 3957 THEN
            sigmoid_f := 259;
        ELSIF x =- 3956 THEN
            sigmoid_f := 259;
        ELSIF x =- 3955 THEN
            sigmoid_f := 259;
        ELSIF x =- 3954 THEN
            sigmoid_f := 259;
        ELSIF x =- 3953 THEN
            sigmoid_f := 259;
        ELSIF x =- 3952 THEN
            sigmoid_f := 259;
        ELSIF x =- 3951 THEN
            sigmoid_f := 259;
        ELSIF x =- 3950 THEN
            sigmoid_f := 259;
        ELSIF x =- 3949 THEN
            sigmoid_f := 260;
        ELSIF x =- 3948 THEN
            sigmoid_f := 260;
        ELSIF x =- 3947 THEN
            sigmoid_f := 260;
        ELSIF x =- 3946 THEN
            sigmoid_f := 260;
        ELSIF x =- 3945 THEN
            sigmoid_f := 260;
        ELSIF x =- 3944 THEN
            sigmoid_f := 260;
        ELSIF x =- 3943 THEN
            sigmoid_f := 260;
        ELSIF x =- 3942 THEN
            sigmoid_f := 260;
        ELSIF x =- 3941 THEN
            sigmoid_f := 261;
        ELSIF x =- 3940 THEN
            sigmoid_f := 261;
        ELSIF x =- 3939 THEN
            sigmoid_f := 261;
        ELSIF x =- 3938 THEN
            sigmoid_f := 261;
        ELSIF x =- 3937 THEN
            sigmoid_f := 261;
        ELSIF x =- 3936 THEN
            sigmoid_f := 261;
        ELSIF x =- 3935 THEN
            sigmoid_f := 261;
        ELSIF x =- 3934 THEN
            sigmoid_f := 261;
        ELSIF x =- 3933 THEN
            sigmoid_f := 261;
        ELSIF x =- 3932 THEN
            sigmoid_f := 262;
        ELSIF x =- 3931 THEN
            sigmoid_f := 262;
        ELSIF x =- 3930 THEN
            sigmoid_f := 262;
        ELSIF x =- 3929 THEN
            sigmoid_f := 262;
        ELSIF x =- 3928 THEN
            sigmoid_f := 262;
        ELSIF x =- 3927 THEN
            sigmoid_f := 262;
        ELSIF x =- 3926 THEN
            sigmoid_f := 262;
        ELSIF x =- 3925 THEN
            sigmoid_f := 262;
        ELSIF x =- 3924 THEN
            sigmoid_f := 262;
        ELSIF x =- 3923 THEN
            sigmoid_f := 263;
        ELSIF x =- 3922 THEN
            sigmoid_f := 263;
        ELSIF x =- 3921 THEN
            sigmoid_f := 263;
        ELSIF x =- 3920 THEN
            sigmoid_f := 263;
        ELSIF x =- 3919 THEN
            sigmoid_f := 263;
        ELSIF x =- 3918 THEN
            sigmoid_f := 263;
        ELSIF x =- 3917 THEN
            sigmoid_f := 263;
        ELSIF x =- 3916 THEN
            sigmoid_f := 263;
        ELSIF x =- 3915 THEN
            sigmoid_f := 264;
        ELSIF x =- 3914 THEN
            sigmoid_f := 264;
        ELSIF x =- 3913 THEN
            sigmoid_f := 264;
        ELSIF x =- 3912 THEN
            sigmoid_f := 264;
        ELSIF x =- 3911 THEN
            sigmoid_f := 264;
        ELSIF x =- 3910 THEN
            sigmoid_f := 264;
        ELSIF x =- 3909 THEN
            sigmoid_f := 264;
        ELSIF x =- 3908 THEN
            sigmoid_f := 264;
        ELSIF x =- 3907 THEN
            sigmoid_f := 264;
        ELSIF x =- 3906 THEN
            sigmoid_f := 265;
        ELSIF x =- 3905 THEN
            sigmoid_f := 265;
        ELSIF x =- 3904 THEN
            sigmoid_f := 265;
        ELSIF x =- 3903 THEN
            sigmoid_f := 265;
        ELSIF x =- 3902 THEN
            sigmoid_f := 265;
        ELSIF x =- 3901 THEN
            sigmoid_f := 265;
        ELSIF x =- 3900 THEN
            sigmoid_f := 265;
        ELSIF x =- 3899 THEN
            sigmoid_f := 265;
        ELSIF x =- 3898 THEN
            sigmoid_f := 266;
        ELSIF x =- 3897 THEN
            sigmoid_f := 266;
        ELSIF x =- 3896 THEN
            sigmoid_f := 266;
        ELSIF x =- 3895 THEN
            sigmoid_f := 266;
        ELSIF x =- 3894 THEN
            sigmoid_f := 266;
        ELSIF x =- 3893 THEN
            sigmoid_f := 266;
        ELSIF x =- 3892 THEN
            sigmoid_f := 266;
        ELSIF x =- 3891 THEN
            sigmoid_f := 266;
        ELSIF x =- 3890 THEN
            sigmoid_f := 266;
        ELSIF x =- 3889 THEN
            sigmoid_f := 267;
        ELSIF x =- 3888 THEN
            sigmoid_f := 267;
        ELSIF x =- 3887 THEN
            sigmoid_f := 267;
        ELSIF x =- 3886 THEN
            sigmoid_f := 267;
        ELSIF x =- 3885 THEN
            sigmoid_f := 267;
        ELSIF x =- 3884 THEN
            sigmoid_f := 267;
        ELSIF x =- 3883 THEN
            sigmoid_f := 267;
        ELSIF x =- 3882 THEN
            sigmoid_f := 267;
        ELSIF x =- 3881 THEN
            sigmoid_f := 267;
        ELSIF x =- 3880 THEN
            sigmoid_f := 268;
        ELSIF x =- 3879 THEN
            sigmoid_f := 268;
        ELSIF x =- 3878 THEN
            sigmoid_f := 268;
        ELSIF x =- 3877 THEN
            sigmoid_f := 268;
        ELSIF x =- 3876 THEN
            sigmoid_f := 268;
        ELSIF x =- 3875 THEN
            sigmoid_f := 268;
        ELSIF x =- 3874 THEN
            sigmoid_f := 268;
        ELSIF x =- 3873 THEN
            sigmoid_f := 268;
        ELSIF x =- 3872 THEN
            sigmoid_f := 269;
        ELSIF x =- 3871 THEN
            sigmoid_f := 269;
        ELSIF x =- 3870 THEN
            sigmoid_f := 269;
        ELSIF x =- 3869 THEN
            sigmoid_f := 269;
        ELSIF x =- 3868 THEN
            sigmoid_f := 269;
        ELSIF x =- 3867 THEN
            sigmoid_f := 269;
        ELSIF x =- 3866 THEN
            sigmoid_f := 269;
        ELSIF x =- 3865 THEN
            sigmoid_f := 269;
        ELSIF x =- 3864 THEN
            sigmoid_f := 269;
        ELSIF x =- 3863 THEN
            sigmoid_f := 270;
        ELSIF x =- 3862 THEN
            sigmoid_f := 270;
        ELSIF x =- 3861 THEN
            sigmoid_f := 270;
        ELSIF x =- 3860 THEN
            sigmoid_f := 270;
        ELSIF x =- 3859 THEN
            sigmoid_f := 270;
        ELSIF x =- 3858 THEN
            sigmoid_f := 270;
        ELSIF x =- 3857 THEN
            sigmoid_f := 270;
        ELSIF x =- 3856 THEN
            sigmoid_f := 270;
        ELSIF x =- 3855 THEN
            sigmoid_f := 271;
        ELSIF x =- 3854 THEN
            sigmoid_f := 271;
        ELSIF x =- 3853 THEN
            sigmoid_f := 271;
        ELSIF x =- 3852 THEN
            sigmoid_f := 271;
        ELSIF x =- 3851 THEN
            sigmoid_f := 271;
        ELSIF x =- 3850 THEN
            sigmoid_f := 271;
        ELSIF x =- 3849 THEN
            sigmoid_f := 271;
        ELSIF x =- 3848 THEN
            sigmoid_f := 271;
        ELSIF x =- 3847 THEN
            sigmoid_f := 271;
        ELSIF x =- 3846 THEN
            sigmoid_f := 272;
        ELSIF x =- 3845 THEN
            sigmoid_f := 272;
        ELSIF x =- 3844 THEN
            sigmoid_f := 272;
        ELSIF x =- 3843 THEN
            sigmoid_f := 272;
        ELSIF x =- 3842 THEN
            sigmoid_f := 272;
        ELSIF x =- 3841 THEN
            sigmoid_f := 272;
        ELSIF x =- 3840 THEN
            sigmoid_f := 272;
        ELSIF x =- 3839 THEN
            sigmoid_f := 272;
        ELSIF x =- 3838 THEN
            sigmoid_f := 272;
        ELSIF x =- 3837 THEN
            sigmoid_f := 273;
        ELSIF x =- 3836 THEN
            sigmoid_f := 273;
        ELSIF x =- 3835 THEN
            sigmoid_f := 273;
        ELSIF x =- 3834 THEN
            sigmoid_f := 273;
        ELSIF x =- 3833 THEN
            sigmoid_f := 273;
        ELSIF x =- 3832 THEN
            sigmoid_f := 273;
        ELSIF x =- 3831 THEN
            sigmoid_f := 273;
        ELSIF x =- 3830 THEN
            sigmoid_f := 273;
        ELSIF x =- 3829 THEN
            sigmoid_f := 274;
        ELSIF x =- 3828 THEN
            sigmoid_f := 274;
        ELSIF x =- 3827 THEN
            sigmoid_f := 274;
        ELSIF x =- 3826 THEN
            sigmoid_f := 274;
        ELSIF x =- 3825 THEN
            sigmoid_f := 274;
        ELSIF x =- 3824 THEN
            sigmoid_f := 274;
        ELSIF x =- 3823 THEN
            sigmoid_f := 274;
        ELSIF x =- 3822 THEN
            sigmoid_f := 274;
        ELSIF x =- 3821 THEN
            sigmoid_f := 274;
        ELSIF x =- 3820 THEN
            sigmoid_f := 275;
        ELSIF x =- 3819 THEN
            sigmoid_f := 275;
        ELSIF x =- 3818 THEN
            sigmoid_f := 275;
        ELSIF x =- 3817 THEN
            sigmoid_f := 275;
        ELSIF x =- 3816 THEN
            sigmoid_f := 275;
        ELSIF x =- 3815 THEN
            sigmoid_f := 275;
        ELSIF x =- 3814 THEN
            sigmoid_f := 275;
        ELSIF x =- 3813 THEN
            sigmoid_f := 275;
        ELSIF x =- 3812 THEN
            sigmoid_f := 276;
        ELSIF x =- 3811 THEN
            sigmoid_f := 276;
        ELSIF x =- 3810 THEN
            sigmoid_f := 276;
        ELSIF x =- 3809 THEN
            sigmoid_f := 276;
        ELSIF x =- 3808 THEN
            sigmoid_f := 276;
        ELSIF x =- 3807 THEN
            sigmoid_f := 276;
        ELSIF x =- 3806 THEN
            sigmoid_f := 276;
        ELSIF x =- 3805 THEN
            sigmoid_f := 276;
        ELSIF x =- 3804 THEN
            sigmoid_f := 276;
        ELSIF x =- 3803 THEN
            sigmoid_f := 277;
        ELSIF x =- 3802 THEN
            sigmoid_f := 277;
        ELSIF x =- 3801 THEN
            sigmoid_f := 277;
        ELSIF x =- 3800 THEN
            sigmoid_f := 277;
        ELSIF x =- 3799 THEN
            sigmoid_f := 277;
        ELSIF x =- 3798 THEN
            sigmoid_f := 277;
        ELSIF x =- 3797 THEN
            sigmoid_f := 277;
        ELSIF x =- 3796 THEN
            sigmoid_f := 277;
        ELSIF x =- 3795 THEN
            sigmoid_f := 277;
        ELSIF x =- 3794 THEN
            sigmoid_f := 278;
        ELSIF x =- 3793 THEN
            sigmoid_f := 278;
        ELSIF x =- 3792 THEN
            sigmoid_f := 278;
        ELSIF x =- 3791 THEN
            sigmoid_f := 278;
        ELSIF x =- 3790 THEN
            sigmoid_f := 278;
        ELSIF x =- 3789 THEN
            sigmoid_f := 278;
        ELSIF x =- 3788 THEN
            sigmoid_f := 278;
        ELSIF x =- 3787 THEN
            sigmoid_f := 278;
        ELSIF x =- 3786 THEN
            sigmoid_f := 279;
        ELSIF x =- 3785 THEN
            sigmoid_f := 279;
        ELSIF x =- 3784 THEN
            sigmoid_f := 279;
        ELSIF x =- 3783 THEN
            sigmoid_f := 279;
        ELSIF x =- 3782 THEN
            sigmoid_f := 279;
        ELSIF x =- 3781 THEN
            sigmoid_f := 279;
        ELSIF x =- 3780 THEN
            sigmoid_f := 279;
        ELSIF x =- 3779 THEN
            sigmoid_f := 279;
        ELSIF x =- 3778 THEN
            sigmoid_f := 279;
        ELSIF x =- 3777 THEN
            sigmoid_f := 280;
        ELSIF x =- 3776 THEN
            sigmoid_f := 280;
        ELSIF x =- 3775 THEN
            sigmoid_f := 280;
        ELSIF x =- 3774 THEN
            sigmoid_f := 280;
        ELSIF x =- 3773 THEN
            sigmoid_f := 280;
        ELSIF x =- 3772 THEN
            sigmoid_f := 280;
        ELSIF x =- 3771 THEN
            sigmoid_f := 280;
        ELSIF x =- 3770 THEN
            sigmoid_f := 280;
        ELSIF x =- 3769 THEN
            sigmoid_f := 281;
        ELSIF x =- 3768 THEN
            sigmoid_f := 281;
        ELSIF x =- 3767 THEN
            sigmoid_f := 281;
        ELSIF x =- 3766 THEN
            sigmoid_f := 281;
        ELSIF x =- 3765 THEN
            sigmoid_f := 281;
        ELSIF x =- 3764 THEN
            sigmoid_f := 281;
        ELSIF x =- 3763 THEN
            sigmoid_f := 281;
        ELSIF x =- 3762 THEN
            sigmoid_f := 281;
        ELSIF x =- 3761 THEN
            sigmoid_f := 281;
        ELSIF x =- 3760 THEN
            sigmoid_f := 282;
        ELSIF x =- 3759 THEN
            sigmoid_f := 282;
        ELSIF x =- 3758 THEN
            sigmoid_f := 282;
        ELSIF x =- 3757 THEN
            sigmoid_f := 282;
        ELSIF x =- 3756 THEN
            sigmoid_f := 282;
        ELSIF x =- 3755 THEN
            sigmoid_f := 282;
        ELSIF x =- 3754 THEN
            sigmoid_f := 282;
        ELSIF x =- 3753 THEN
            sigmoid_f := 282;
        ELSIF x =- 3752 THEN
            sigmoid_f := 282;
        ELSIF x =- 3751 THEN
            sigmoid_f := 283;
        ELSIF x =- 3750 THEN
            sigmoid_f := 283;
        ELSIF x =- 3749 THEN
            sigmoid_f := 283;
        ELSIF x =- 3748 THEN
            sigmoid_f := 283;
        ELSIF x =- 3747 THEN
            sigmoid_f := 283;
        ELSIF x =- 3746 THEN
            sigmoid_f := 283;
        ELSIF x =- 3745 THEN
            sigmoid_f := 283;
        ELSIF x =- 3744 THEN
            sigmoid_f := 283;
        ELSIF x =- 3743 THEN
            sigmoid_f := 284;
        ELSIF x =- 3742 THEN
            sigmoid_f := 284;
        ELSIF x =- 3741 THEN
            sigmoid_f := 284;
        ELSIF x =- 3740 THEN
            sigmoid_f := 284;
        ELSIF x =- 3739 THEN
            sigmoid_f := 284;
        ELSIF x =- 3738 THEN
            sigmoid_f := 284;
        ELSIF x =- 3737 THEN
            sigmoid_f := 284;
        ELSIF x =- 3736 THEN
            sigmoid_f := 284;
        ELSIF x =- 3735 THEN
            sigmoid_f := 284;
        ELSIF x =- 3734 THEN
            sigmoid_f := 285;
        ELSIF x =- 3733 THEN
            sigmoid_f := 285;
        ELSIF x =- 3732 THEN
            sigmoid_f := 285;
        ELSIF x =- 3731 THEN
            sigmoid_f := 285;
        ELSIF x =- 3730 THEN
            sigmoid_f := 285;
        ELSIF x =- 3729 THEN
            sigmoid_f := 285;
        ELSIF x =- 3728 THEN
            sigmoid_f := 285;
        ELSIF x =- 3727 THEN
            sigmoid_f := 285;
        ELSIF x =- 3726 THEN
            sigmoid_f := 285;
        ELSIF x =- 3725 THEN
            sigmoid_f := 286;
        ELSIF x =- 3724 THEN
            sigmoid_f := 286;
        ELSIF x =- 3723 THEN
            sigmoid_f := 286;
        ELSIF x =- 3722 THEN
            sigmoid_f := 286;
        ELSIF x =- 3721 THEN
            sigmoid_f := 286;
        ELSIF x =- 3720 THEN
            sigmoid_f := 286;
        ELSIF x =- 3719 THEN
            sigmoid_f := 286;
        ELSIF x =- 3718 THEN
            sigmoid_f := 286;
        ELSIF x =- 3717 THEN
            sigmoid_f := 287;
        ELSIF x =- 3716 THEN
            sigmoid_f := 287;
        ELSIF x =- 3715 THEN
            sigmoid_f := 287;
        ELSIF x =- 3714 THEN
            sigmoid_f := 287;
        ELSIF x =- 3713 THEN
            sigmoid_f := 287;
        ELSIF x =- 3712 THEN
            sigmoid_f := 287;
        ELSIF x =- 3711 THEN
            sigmoid_f := 287;
        ELSIF x =- 3710 THEN
            sigmoid_f := 287;
        ELSIF x =- 3709 THEN
            sigmoid_f := 287;
        ELSIF x =- 3708 THEN
            sigmoid_f := 288;
        ELSIF x =- 3707 THEN
            sigmoid_f := 288;
        ELSIF x =- 3706 THEN
            sigmoid_f := 288;
        ELSIF x =- 3705 THEN
            sigmoid_f := 288;
        ELSIF x =- 3704 THEN
            sigmoid_f := 288;
        ELSIF x =- 3703 THEN
            sigmoid_f := 288;
        ELSIF x =- 3702 THEN
            sigmoid_f := 288;
        ELSIF x =- 3701 THEN
            sigmoid_f := 288;
        ELSIF x =- 3700 THEN
            sigmoid_f := 289;
        ELSIF x =- 3699 THEN
            sigmoid_f := 289;
        ELSIF x =- 3698 THEN
            sigmoid_f := 289;
        ELSIF x =- 3697 THEN
            sigmoid_f := 289;
        ELSIF x =- 3696 THEN
            sigmoid_f := 289;
        ELSIF x =- 3695 THEN
            sigmoid_f := 289;
        ELSIF x =- 3694 THEN
            sigmoid_f := 289;
        ELSIF x =- 3693 THEN
            sigmoid_f := 289;
        ELSIF x =- 3692 THEN
            sigmoid_f := 289;
        ELSIF x =- 3691 THEN
            sigmoid_f := 290;
        ELSIF x =- 3690 THEN
            sigmoid_f := 290;
        ELSIF x =- 3689 THEN
            sigmoid_f := 290;
        ELSIF x =- 3688 THEN
            sigmoid_f := 290;
        ELSIF x =- 3687 THEN
            sigmoid_f := 290;
        ELSIF x =- 3686 THEN
            sigmoid_f := 290;
        ELSIF x =- 3685 THEN
            sigmoid_f := 290;
        ELSIF x =- 3684 THEN
            sigmoid_f := 290;
        ELSIF x =- 3683 THEN
            sigmoid_f := 290;
        ELSIF x =- 3682 THEN
            sigmoid_f := 291;
        ELSIF x =- 3681 THEN
            sigmoid_f := 291;
        ELSIF x =- 3680 THEN
            sigmoid_f := 291;
        ELSIF x =- 3679 THEN
            sigmoid_f := 291;
        ELSIF x =- 3678 THEN
            sigmoid_f := 291;
        ELSIF x =- 3677 THEN
            sigmoid_f := 291;
        ELSIF x =- 3676 THEN
            sigmoid_f := 291;
        ELSIF x =- 3675 THEN
            sigmoid_f := 291;
        ELSIF x =- 3674 THEN
            sigmoid_f := 292;
        ELSIF x =- 3673 THEN
            sigmoid_f := 292;
        ELSIF x =- 3672 THEN
            sigmoid_f := 292;
        ELSIF x =- 3671 THEN
            sigmoid_f := 292;
        ELSIF x =- 3670 THEN
            sigmoid_f := 292;
        ELSIF x =- 3669 THEN
            sigmoid_f := 292;
        ELSIF x =- 3668 THEN
            sigmoid_f := 292;
        ELSIF x =- 3667 THEN
            sigmoid_f := 292;
        ELSIF x =- 3666 THEN
            sigmoid_f := 292;
        ELSIF x =- 3665 THEN
            sigmoid_f := 293;
        ELSIF x =- 3664 THEN
            sigmoid_f := 293;
        ELSIF x =- 3663 THEN
            sigmoid_f := 293;
        ELSIF x =- 3662 THEN
            sigmoid_f := 293;
        ELSIF x =- 3661 THEN
            sigmoid_f := 293;
        ELSIF x =- 3660 THEN
            sigmoid_f := 293;
        ELSIF x =- 3659 THEN
            sigmoid_f := 293;
        ELSIF x =- 3658 THEN
            sigmoid_f := 293;
        ELSIF x =- 3657 THEN
            sigmoid_f := 294;
        ELSIF x =- 3656 THEN
            sigmoid_f := 294;
        ELSIF x =- 3655 THEN
            sigmoid_f := 294;
        ELSIF x =- 3654 THEN
            sigmoid_f := 294;
        ELSIF x =- 3653 THEN
            sigmoid_f := 294;
        ELSIF x =- 3652 THEN
            sigmoid_f := 294;
        ELSIF x =- 3651 THEN
            sigmoid_f := 294;
        ELSIF x =- 3650 THEN
            sigmoid_f := 294;
        ELSIF x =- 3649 THEN
            sigmoid_f := 294;
        ELSIF x =- 3648 THEN
            sigmoid_f := 295;
        ELSIF x =- 3647 THEN
            sigmoid_f := 295;
        ELSIF x =- 3646 THEN
            sigmoid_f := 295;
        ELSIF x =- 3645 THEN
            sigmoid_f := 295;
        ELSIF x =- 3644 THEN
            sigmoid_f := 295;
        ELSIF x =- 3643 THEN
            sigmoid_f := 295;
        ELSIF x =- 3642 THEN
            sigmoid_f := 295;
        ELSIF x =- 3641 THEN
            sigmoid_f := 295;
        ELSIF x =- 3640 THEN
            sigmoid_f := 295;
        ELSIF x =- 3639 THEN
            sigmoid_f := 296;
        ELSIF x =- 3638 THEN
            sigmoid_f := 296;
        ELSIF x =- 3637 THEN
            sigmoid_f := 296;
        ELSIF x =- 3636 THEN
            sigmoid_f := 296;
        ELSIF x =- 3635 THEN
            sigmoid_f := 296;
        ELSIF x =- 3634 THEN
            sigmoid_f := 296;
        ELSIF x =- 3633 THEN
            sigmoid_f := 296;
        ELSIF x =- 3632 THEN
            sigmoid_f := 296;
        ELSIF x =- 3631 THEN
            sigmoid_f := 297;
        ELSIF x =- 3630 THEN
            sigmoid_f := 297;
        ELSIF x =- 3629 THEN
            sigmoid_f := 297;
        ELSIF x =- 3628 THEN
            sigmoid_f := 297;
        ELSIF x =- 3627 THEN
            sigmoid_f := 297;
        ELSIF x =- 3626 THEN
            sigmoid_f := 297;
        ELSIF x =- 3625 THEN
            sigmoid_f := 297;
        ELSIF x =- 3624 THEN
            sigmoid_f := 297;
        ELSIF x =- 3623 THEN
            sigmoid_f := 297;
        ELSIF x =- 3622 THEN
            sigmoid_f := 298;
        ELSIF x =- 3621 THEN
            sigmoid_f := 298;
        ELSIF x =- 3620 THEN
            sigmoid_f := 298;
        ELSIF x =- 3619 THEN
            sigmoid_f := 298;
        ELSIF x =- 3618 THEN
            sigmoid_f := 298;
        ELSIF x =- 3617 THEN
            sigmoid_f := 298;
        ELSIF x =- 3616 THEN
            sigmoid_f := 298;
        ELSIF x =- 3615 THEN
            sigmoid_f := 298;
        ELSIF x =- 3614 THEN
            sigmoid_f := 299;
        ELSIF x =- 3613 THEN
            sigmoid_f := 299;
        ELSIF x =- 3612 THEN
            sigmoid_f := 299;
        ELSIF x =- 3611 THEN
            sigmoid_f := 299;
        ELSIF x =- 3610 THEN
            sigmoid_f := 299;
        ELSIF x =- 3609 THEN
            sigmoid_f := 299;
        ELSIF x =- 3608 THEN
            sigmoid_f := 299;
        ELSIF x =- 3607 THEN
            sigmoid_f := 299;
        ELSIF x =- 3606 THEN
            sigmoid_f := 299;
        ELSIF x =- 3605 THEN
            sigmoid_f := 300;
        ELSIF x =- 3604 THEN
            sigmoid_f := 300;
        ELSIF x =- 3603 THEN
            sigmoid_f := 300;
        ELSIF x =- 3602 THEN
            sigmoid_f := 300;
        ELSIF x =- 3601 THEN
            sigmoid_f := 300;
        ELSIF x =- 3600 THEN
            sigmoid_f := 300;
        ELSIF x =- 3599 THEN
            sigmoid_f := 300;
        ELSIF x =- 3598 THEN
            sigmoid_f := 300;
        ELSIF x =- 3597 THEN
            sigmoid_f := 300;
        ELSIF x =- 3596 THEN
            sigmoid_f := 301;
        ELSIF x =- 3595 THEN
            sigmoid_f := 301;
        ELSIF x =- 3594 THEN
            sigmoid_f := 301;
        ELSIF x =- 3593 THEN
            sigmoid_f := 301;
        ELSIF x =- 3592 THEN
            sigmoid_f := 301;
        ELSIF x =- 3591 THEN
            sigmoid_f := 301;
        ELSIF x =- 3590 THEN
            sigmoid_f := 301;
        ELSIF x =- 3589 THEN
            sigmoid_f := 301;
        ELSIF x =- 3588 THEN
            sigmoid_f := 302;
        ELSIF x =- 3587 THEN
            sigmoid_f := 302;
        ELSIF x =- 3586 THEN
            sigmoid_f := 302;
        ELSIF x =- 3585 THEN
            sigmoid_f := 302;
        ELSIF x =- 3584 THEN
            sigmoid_f := 302;
        ELSIF x =- 3583 THEN
            sigmoid_f := 302;
        ELSIF x =- 3582 THEN
            sigmoid_f := 302;
        ELSIF x =- 3581 THEN
            sigmoid_f := 302;
        ELSIF x =- 3580 THEN
            sigmoid_f := 302;
        ELSIF x =- 3579 THEN
            sigmoid_f := 302;
        ELSIF x =- 3578 THEN
            sigmoid_f := 303;
        ELSIF x =- 3577 THEN
            sigmoid_f := 303;
        ELSIF x =- 3576 THEN
            sigmoid_f := 303;
        ELSIF x =- 3575 THEN
            sigmoid_f := 303;
        ELSIF x =- 3574 THEN
            sigmoid_f := 303;
        ELSIF x =- 3573 THEN
            sigmoid_f := 303;
        ELSIF x =- 3572 THEN
            sigmoid_f := 303;
        ELSIF x =- 3571 THEN
            sigmoid_f := 304;
        ELSIF x =- 3570 THEN
            sigmoid_f := 304;
        ELSIF x =- 3569 THEN
            sigmoid_f := 304;
        ELSIF x =- 3568 THEN
            sigmoid_f := 304;
        ELSIF x =- 3567 THEN
            sigmoid_f := 304;
        ELSIF x =- 3566 THEN
            sigmoid_f := 304;
        ELSIF x =- 3565 THEN
            sigmoid_f := 304;
        ELSIF x =- 3564 THEN
            sigmoid_f := 304;
        ELSIF x =- 3563 THEN
            sigmoid_f := 305;
        ELSIF x =- 3562 THEN
            sigmoid_f := 305;
        ELSIF x =- 3561 THEN
            sigmoid_f := 305;
        ELSIF x =- 3560 THEN
            sigmoid_f := 305;
        ELSIF x =- 3559 THEN
            sigmoid_f := 305;
        ELSIF x =- 3558 THEN
            sigmoid_f := 305;
        ELSIF x =- 3557 THEN
            sigmoid_f := 305;
        ELSIF x =- 3556 THEN
            sigmoid_f := 306;
        ELSIF x =- 3555 THEN
            sigmoid_f := 306;
        ELSIF x =- 3554 THEN
            sigmoid_f := 306;
        ELSIF x =- 3553 THEN
            sigmoid_f := 306;
        ELSIF x =- 3552 THEN
            sigmoid_f := 306;
        ELSIF x =- 3551 THEN
            sigmoid_f := 306;
        ELSIF x =- 3550 THEN
            sigmoid_f := 306;
        ELSIF x =- 3549 THEN
            sigmoid_f := 307;
        ELSIF x =- 3548 THEN
            sigmoid_f := 307;
        ELSIF x =- 3547 THEN
            sigmoid_f := 307;
        ELSIF x =- 3546 THEN
            sigmoid_f := 307;
        ELSIF x =- 3545 THEN
            sigmoid_f := 307;
        ELSIF x =- 3544 THEN
            sigmoid_f := 307;
        ELSIF x =- 3543 THEN
            sigmoid_f := 307;
        ELSIF x =- 3542 THEN
            sigmoid_f := 308;
        ELSIF x =- 3541 THEN
            sigmoid_f := 308;
        ELSIF x =- 3540 THEN
            sigmoid_f := 308;
        ELSIF x =- 3539 THEN
            sigmoid_f := 308;
        ELSIF x =- 3538 THEN
            sigmoid_f := 308;
        ELSIF x =- 3537 THEN
            sigmoid_f := 308;
        ELSIF x =- 3536 THEN
            sigmoid_f := 308;
        ELSIF x =- 3535 THEN
            sigmoid_f := 308;
        ELSIF x =- 3534 THEN
            sigmoid_f := 309;
        ELSIF x =- 3533 THEN
            sigmoid_f := 309;
        ELSIF x =- 3532 THEN
            sigmoid_f := 309;
        ELSIF x =- 3531 THEN
            sigmoid_f := 309;
        ELSIF x =- 3530 THEN
            sigmoid_f := 309;
        ELSIF x =- 3529 THEN
            sigmoid_f := 309;
        ELSIF x =- 3528 THEN
            sigmoid_f := 309;
        ELSIF x =- 3527 THEN
            sigmoid_f := 310;
        ELSIF x =- 3526 THEN
            sigmoid_f := 310;
        ELSIF x =- 3525 THEN
            sigmoid_f := 310;
        ELSIF x =- 3524 THEN
            sigmoid_f := 310;
        ELSIF x =- 3523 THEN
            sigmoid_f := 310;
        ELSIF x =- 3522 THEN
            sigmoid_f := 310;
        ELSIF x =- 3521 THEN
            sigmoid_f := 310;
        ELSIF x =- 3520 THEN
            sigmoid_f := 311;
        ELSIF x =- 3519 THEN
            sigmoid_f := 311;
        ELSIF x =- 3518 THEN
            sigmoid_f := 311;
        ELSIF x =- 3517 THEN
            sigmoid_f := 311;
        ELSIF x =- 3516 THEN
            sigmoid_f := 311;
        ELSIF x =- 3515 THEN
            sigmoid_f := 311;
        ELSIF x =- 3514 THEN
            sigmoid_f := 311;
        ELSIF x =- 3513 THEN
            sigmoid_f := 311;
        ELSIF x =- 3512 THEN
            sigmoid_f := 312;
        ELSIF x =- 3511 THEN
            sigmoid_f := 312;
        ELSIF x =- 3510 THEN
            sigmoid_f := 312;
        ELSIF x =- 3509 THEN
            sigmoid_f := 312;
        ELSIF x =- 3508 THEN
            sigmoid_f := 312;
        ELSIF x =- 3507 THEN
            sigmoid_f := 312;
        ELSIF x =- 3506 THEN
            sigmoid_f := 312;
        ELSIF x =- 3505 THEN
            sigmoid_f := 313;
        ELSIF x =- 3504 THEN
            sigmoid_f := 313;
        ELSIF x =- 3503 THEN
            sigmoid_f := 313;
        ELSIF x =- 3502 THEN
            sigmoid_f := 313;
        ELSIF x =- 3501 THEN
            sigmoid_f := 313;
        ELSIF x =- 3500 THEN
            sigmoid_f := 313;
        ELSIF x =- 3499 THEN
            sigmoid_f := 313;
        ELSIF x =- 3498 THEN
            sigmoid_f := 314;
        ELSIF x =- 3497 THEN
            sigmoid_f := 314;
        ELSIF x =- 3496 THEN
            sigmoid_f := 314;
        ELSIF x =- 3495 THEN
            sigmoid_f := 314;
        ELSIF x =- 3494 THEN
            sigmoid_f := 314;
        ELSIF x =- 3493 THEN
            sigmoid_f := 314;
        ELSIF x =- 3492 THEN
            sigmoid_f := 314;
        ELSIF x =- 3491 THEN
            sigmoid_f := 315;
        ELSIF x =- 3490 THEN
            sigmoid_f := 315;
        ELSIF x =- 3489 THEN
            sigmoid_f := 315;
        ELSIF x =- 3488 THEN
            sigmoid_f := 315;
        ELSIF x =- 3487 THEN
            sigmoid_f := 315;
        ELSIF x =- 3486 THEN
            sigmoid_f := 315;
        ELSIF x =- 3485 THEN
            sigmoid_f := 315;
        ELSIF x =- 3484 THEN
            sigmoid_f := 315;
        ELSIF x =- 3483 THEN
            sigmoid_f := 316;
        ELSIF x =- 3482 THEN
            sigmoid_f := 316;
        ELSIF x =- 3481 THEN
            sigmoid_f := 316;
        ELSIF x =- 3480 THEN
            sigmoid_f := 316;
        ELSIF x =- 3479 THEN
            sigmoid_f := 316;
        ELSIF x =- 3478 THEN
            sigmoid_f := 316;
        ELSIF x =- 3477 THEN
            sigmoid_f := 316;
        ELSIF x =- 3476 THEN
            sigmoid_f := 317;
        ELSIF x =- 3475 THEN
            sigmoid_f := 317;
        ELSIF x =- 3474 THEN
            sigmoid_f := 317;
        ELSIF x =- 3473 THEN
            sigmoid_f := 317;
        ELSIF x =- 3472 THEN
            sigmoid_f := 317;
        ELSIF x =- 3471 THEN
            sigmoid_f := 317;
        ELSIF x =- 3470 THEN
            sigmoid_f := 317;
        ELSIF x =- 3469 THEN
            sigmoid_f := 318;
        ELSIF x =- 3468 THEN
            sigmoid_f := 318;
        ELSIF x =- 3467 THEN
            sigmoid_f := 318;
        ELSIF x =- 3466 THEN
            sigmoid_f := 318;
        ELSIF x =- 3465 THEN
            sigmoid_f := 318;
        ELSIF x =- 3464 THEN
            sigmoid_f := 318;
        ELSIF x =- 3463 THEN
            sigmoid_f := 318;
        ELSIF x =- 3462 THEN
            sigmoid_f := 318;
        ELSIF x =- 3461 THEN
            sigmoid_f := 319;
        ELSIF x =- 3460 THEN
            sigmoid_f := 319;
        ELSIF x =- 3459 THEN
            sigmoid_f := 319;
        ELSIF x =- 3458 THEN
            sigmoid_f := 319;
        ELSIF x =- 3457 THEN
            sigmoid_f := 319;
        ELSIF x =- 3456 THEN
            sigmoid_f := 319;
        ELSIF x =- 3455 THEN
            sigmoid_f := 319;
        ELSIF x =- 3454 THEN
            sigmoid_f := 320;
        ELSIF x =- 3453 THEN
            sigmoid_f := 320;
        ELSIF x =- 3452 THEN
            sigmoid_f := 320;
        ELSIF x =- 3451 THEN
            sigmoid_f := 320;
        ELSIF x =- 3450 THEN
            sigmoid_f := 320;
        ELSIF x =- 3449 THEN
            sigmoid_f := 320;
        ELSIF x =- 3448 THEN
            sigmoid_f := 320;
        ELSIF x =- 3447 THEN
            sigmoid_f := 321;
        ELSIF x =- 3446 THEN
            sigmoid_f := 321;
        ELSIF x =- 3445 THEN
            sigmoid_f := 321;
        ELSIF x =- 3444 THEN
            sigmoid_f := 321;
        ELSIF x =- 3443 THEN
            sigmoid_f := 321;
        ELSIF x =- 3442 THEN
            sigmoid_f := 321;
        ELSIF x =- 3441 THEN
            sigmoid_f := 321;
        ELSIF x =- 3440 THEN
            sigmoid_f := 322;
        ELSIF x =- 3439 THEN
            sigmoid_f := 322;
        ELSIF x =- 3438 THEN
            sigmoid_f := 322;
        ELSIF x =- 3437 THEN
            sigmoid_f := 322;
        ELSIF x =- 3436 THEN
            sigmoid_f := 322;
        ELSIF x =- 3435 THEN
            sigmoid_f := 322;
        ELSIF x =- 3434 THEN
            sigmoid_f := 322;
        ELSIF x =- 3433 THEN
            sigmoid_f := 322;
        ELSIF x =- 3432 THEN
            sigmoid_f := 323;
        ELSIF x =- 3431 THEN
            sigmoid_f := 323;
        ELSIF x =- 3430 THEN
            sigmoid_f := 323;
        ELSIF x =- 3429 THEN
            sigmoid_f := 323;
        ELSIF x =- 3428 THEN
            sigmoid_f := 323;
        ELSIF x =- 3427 THEN
            sigmoid_f := 323;
        ELSIF x =- 3426 THEN
            sigmoid_f := 323;
        ELSIF x =- 3425 THEN
            sigmoid_f := 324;
        ELSIF x =- 3424 THEN
            sigmoid_f := 324;
        ELSIF x =- 3423 THEN
            sigmoid_f := 324;
        ELSIF x =- 3422 THEN
            sigmoid_f := 324;
        ELSIF x =- 3421 THEN
            sigmoid_f := 324;
        ELSIF x =- 3420 THEN
            sigmoid_f := 324;
        ELSIF x =- 3419 THEN
            sigmoid_f := 324;
        ELSIF x =- 3418 THEN
            sigmoid_f := 325;
        ELSIF x =- 3417 THEN
            sigmoid_f := 325;
        ELSIF x =- 3416 THEN
            sigmoid_f := 325;
        ELSIF x =- 3415 THEN
            sigmoid_f := 325;
        ELSIF x =- 3414 THEN
            sigmoid_f := 325;
        ELSIF x =- 3413 THEN
            sigmoid_f := 325;
        ELSIF x =- 3412 THEN
            sigmoid_f := 325;
        ELSIF x =- 3411 THEN
            sigmoid_f := 325;
        ELSIF x =- 3410 THEN
            sigmoid_f := 326;
        ELSIF x =- 3409 THEN
            sigmoid_f := 326;
        ELSIF x =- 3408 THEN
            sigmoid_f := 326;
        ELSIF x =- 3407 THEN
            sigmoid_f := 326;
        ELSIF x =- 3406 THEN
            sigmoid_f := 326;
        ELSIF x =- 3405 THEN
            sigmoid_f := 326;
        ELSIF x =- 3404 THEN
            sigmoid_f := 326;
        ELSIF x =- 3403 THEN
            sigmoid_f := 327;
        ELSIF x =- 3402 THEN
            sigmoid_f := 327;
        ELSIF x =- 3401 THEN
            sigmoid_f := 327;
        ELSIF x =- 3400 THEN
            sigmoid_f := 327;
        ELSIF x =- 3399 THEN
            sigmoid_f := 327;
        ELSIF x =- 3398 THEN
            sigmoid_f := 327;
        ELSIF x =- 3397 THEN
            sigmoid_f := 327;
        ELSIF x =- 3396 THEN
            sigmoid_f := 328;
        ELSIF x =- 3395 THEN
            sigmoid_f := 328;
        ELSIF x =- 3394 THEN
            sigmoid_f := 328;
        ELSIF x =- 3393 THEN
            sigmoid_f := 328;
        ELSIF x =- 3392 THEN
            sigmoid_f := 328;
        ELSIF x =- 3391 THEN
            sigmoid_f := 328;
        ELSIF x =- 3390 THEN
            sigmoid_f := 328;
        ELSIF x =- 3389 THEN
            sigmoid_f := 329;
        ELSIF x =- 3388 THEN
            sigmoid_f := 329;
        ELSIF x =- 3387 THEN
            sigmoid_f := 329;
        ELSIF x =- 3386 THEN
            sigmoid_f := 329;
        ELSIF x =- 3385 THEN
            sigmoid_f := 329;
        ELSIF x =- 3384 THEN
            sigmoid_f := 329;
        ELSIF x =- 3383 THEN
            sigmoid_f := 329;
        ELSIF x =- 3382 THEN
            sigmoid_f := 329;
        ELSIF x =- 3381 THEN
            sigmoid_f := 330;
        ELSIF x =- 3380 THEN
            sigmoid_f := 330;
        ELSIF x =- 3379 THEN
            sigmoid_f := 330;
        ELSIF x =- 3378 THEN
            sigmoid_f := 330;
        ELSIF x =- 3377 THEN
            sigmoid_f := 330;
        ELSIF x =- 3376 THEN
            sigmoid_f := 330;
        ELSIF x =- 3375 THEN
            sigmoid_f := 330;
        ELSIF x =- 3374 THEN
            sigmoid_f := 331;
        ELSIF x =- 3373 THEN
            sigmoid_f := 331;
        ELSIF x =- 3372 THEN
            sigmoid_f := 331;
        ELSIF x =- 3371 THEN
            sigmoid_f := 331;
        ELSIF x =- 3370 THEN
            sigmoid_f := 331;
        ELSIF x =- 3369 THEN
            sigmoid_f := 331;
        ELSIF x =- 3368 THEN
            sigmoid_f := 331;
        ELSIF x =- 3367 THEN
            sigmoid_f := 332;
        ELSIF x =- 3366 THEN
            sigmoid_f := 332;
        ELSIF x =- 3365 THEN
            sigmoid_f := 332;
        ELSIF x =- 3364 THEN
            sigmoid_f := 332;
        ELSIF x =- 3363 THEN
            sigmoid_f := 332;
        ELSIF x =- 3362 THEN
            sigmoid_f := 332;
        ELSIF x =- 3361 THEN
            sigmoid_f := 332;
        ELSIF x =- 3360 THEN
            sigmoid_f := 332;
        ELSIF x =- 3359 THEN
            sigmoid_f := 333;
        ELSIF x =- 3358 THEN
            sigmoid_f := 333;
        ELSIF x =- 3357 THEN
            sigmoid_f := 333;
        ELSIF x =- 3356 THEN
            sigmoid_f := 333;
        ELSIF x =- 3355 THEN
            sigmoid_f := 333;
        ELSIF x =- 3354 THEN
            sigmoid_f := 333;
        ELSIF x =- 3353 THEN
            sigmoid_f := 333;
        ELSIF x =- 3352 THEN
            sigmoid_f := 334;
        ELSIF x =- 3351 THEN
            sigmoid_f := 334;
        ELSIF x =- 3350 THEN
            sigmoid_f := 334;
        ELSIF x =- 3349 THEN
            sigmoid_f := 334;
        ELSIF x =- 3348 THEN
            sigmoid_f := 334;
        ELSIF x =- 3347 THEN
            sigmoid_f := 334;
        ELSIF x =- 3346 THEN
            sigmoid_f := 334;
        ELSIF x =- 3345 THEN
            sigmoid_f := 335;
        ELSIF x =- 3344 THEN
            sigmoid_f := 335;
        ELSIF x =- 3343 THEN
            sigmoid_f := 335;
        ELSIF x =- 3342 THEN
            sigmoid_f := 335;
        ELSIF x =- 3341 THEN
            sigmoid_f := 335;
        ELSIF x =- 3340 THEN
            sigmoid_f := 335;
        ELSIF x =- 3339 THEN
            sigmoid_f := 335;
        ELSIF x =- 3338 THEN
            sigmoid_f := 336;
        ELSIF x =- 3337 THEN
            sigmoid_f := 336;
        ELSIF x =- 3336 THEN
            sigmoid_f := 336;
        ELSIF x =- 3335 THEN
            sigmoid_f := 336;
        ELSIF x =- 3334 THEN
            sigmoid_f := 336;
        ELSIF x =- 3333 THEN
            sigmoid_f := 336;
        ELSIF x =- 3332 THEN
            sigmoid_f := 336;
        ELSIF x =- 3331 THEN
            sigmoid_f := 336;
        ELSIF x =- 3330 THEN
            sigmoid_f := 337;
        ELSIF x =- 3329 THEN
            sigmoid_f := 337;
        ELSIF x =- 3328 THEN
            sigmoid_f := 337;
        ELSIF x =- 3327 THEN
            sigmoid_f := 337;
        ELSIF x =- 3326 THEN
            sigmoid_f := 337;
        ELSIF x =- 3325 THEN
            sigmoid_f := 337;
        ELSIF x =- 3324 THEN
            sigmoid_f := 337;
        ELSIF x =- 3323 THEN
            sigmoid_f := 338;
        ELSIF x =- 3322 THEN
            sigmoid_f := 338;
        ELSIF x =- 3321 THEN
            sigmoid_f := 338;
        ELSIF x =- 3320 THEN
            sigmoid_f := 338;
        ELSIF x =- 3319 THEN
            sigmoid_f := 338;
        ELSIF x =- 3318 THEN
            sigmoid_f := 338;
        ELSIF x =- 3317 THEN
            sigmoid_f := 338;
        ELSIF x =- 3316 THEN
            sigmoid_f := 339;
        ELSIF x =- 3315 THEN
            sigmoid_f := 339;
        ELSIF x =- 3314 THEN
            sigmoid_f := 339;
        ELSIF x =- 3313 THEN
            sigmoid_f := 339;
        ELSIF x =- 3312 THEN
            sigmoid_f := 339;
        ELSIF x =- 3311 THEN
            sigmoid_f := 339;
        ELSIF x =- 3310 THEN
            sigmoid_f := 339;
        ELSIF x =- 3309 THEN
            sigmoid_f := 339;
        ELSIF x =- 3308 THEN
            sigmoid_f := 340;
        ELSIF x =- 3307 THEN
            sigmoid_f := 340;
        ELSIF x =- 3306 THEN
            sigmoid_f := 340;
        ELSIF x =- 3305 THEN
            sigmoid_f := 340;
        ELSIF x =- 3304 THEN
            sigmoid_f := 340;
        ELSIF x =- 3303 THEN
            sigmoid_f := 340;
        ELSIF x =- 3302 THEN
            sigmoid_f := 340;
        ELSIF x =- 3301 THEN
            sigmoid_f := 341;
        ELSIF x =- 3300 THEN
            sigmoid_f := 341;
        ELSIF x =- 3299 THEN
            sigmoid_f := 341;
        ELSIF x =- 3298 THEN
            sigmoid_f := 341;
        ELSIF x =- 3297 THEN
            sigmoid_f := 341;
        ELSIF x =- 3296 THEN
            sigmoid_f := 341;
        ELSIF x =- 3295 THEN
            sigmoid_f := 341;
        ELSIF x =- 3294 THEN
            sigmoid_f := 342;
        ELSIF x =- 3293 THEN
            sigmoid_f := 342;
        ELSIF x =- 3292 THEN
            sigmoid_f := 342;
        ELSIF x =- 3291 THEN
            sigmoid_f := 342;
        ELSIF x =- 3290 THEN
            sigmoid_f := 342;
        ELSIF x =- 3289 THEN
            sigmoid_f := 342;
        ELSIF x =- 3288 THEN
            sigmoid_f := 342;
        ELSIF x =- 3287 THEN
            sigmoid_f := 343;
        ELSIF x =- 3286 THEN
            sigmoid_f := 343;
        ELSIF x =- 3285 THEN
            sigmoid_f := 343;
        ELSIF x =- 3284 THEN
            sigmoid_f := 343;
        ELSIF x =- 3283 THEN
            sigmoid_f := 343;
        ELSIF x =- 3282 THEN
            sigmoid_f := 343;
        ELSIF x =- 3281 THEN
            sigmoid_f := 343;
        ELSIF x =- 3280 THEN
            sigmoid_f := 343;
        ELSIF x =- 3279 THEN
            sigmoid_f := 344;
        ELSIF x =- 3278 THEN
            sigmoid_f := 344;
        ELSIF x =- 3277 THEN
            sigmoid_f := 344;
        ELSIF x =- 3276 THEN
            sigmoid_f := 344;
        ELSIF x =- 3275 THEN
            sigmoid_f := 344;
        ELSIF x =- 3274 THEN
            sigmoid_f := 344;
        ELSIF x =- 3273 THEN
            sigmoid_f := 344;
        ELSIF x =- 3272 THEN
            sigmoid_f := 345;
        ELSIF x =- 3271 THEN
            sigmoid_f := 345;
        ELSIF x =- 3270 THEN
            sigmoid_f := 345;
        ELSIF x =- 3269 THEN
            sigmoid_f := 345;
        ELSIF x =- 3268 THEN
            sigmoid_f := 345;
        ELSIF x =- 3267 THEN
            sigmoid_f := 345;
        ELSIF x =- 3266 THEN
            sigmoid_f := 345;
        ELSIF x =- 3265 THEN
            sigmoid_f := 346;
        ELSIF x =- 3264 THEN
            sigmoid_f := 346;
        ELSIF x =- 3263 THEN
            sigmoid_f := 346;
        ELSIF x =- 3262 THEN
            sigmoid_f := 346;
        ELSIF x =- 3261 THEN
            sigmoid_f := 346;
        ELSIF x =- 3260 THEN
            sigmoid_f := 346;
        ELSIF x =- 3259 THEN
            sigmoid_f := 346;
        ELSIF x =- 3258 THEN
            sigmoid_f := 346;
        ELSIF x =- 3257 THEN
            sigmoid_f := 347;
        ELSIF x =- 3256 THEN
            sigmoid_f := 347;
        ELSIF x =- 3255 THEN
            sigmoid_f := 347;
        ELSIF x =- 3254 THEN
            sigmoid_f := 347;
        ELSIF x =- 3253 THEN
            sigmoid_f := 347;
        ELSIF x =- 3252 THEN
            sigmoid_f := 347;
        ELSIF x =- 3251 THEN
            sigmoid_f := 347;
        ELSIF x =- 3250 THEN
            sigmoid_f := 348;
        ELSIF x =- 3249 THEN
            sigmoid_f := 348;
        ELSIF x =- 3248 THEN
            sigmoid_f := 348;
        ELSIF x =- 3247 THEN
            sigmoid_f := 348;
        ELSIF x =- 3246 THEN
            sigmoid_f := 348;
        ELSIF x =- 3245 THEN
            sigmoid_f := 348;
        ELSIF x =- 3244 THEN
            sigmoid_f := 348;
        ELSIF x =- 3243 THEN
            sigmoid_f := 349;
        ELSIF x =- 3242 THEN
            sigmoid_f := 349;
        ELSIF x =- 3241 THEN
            sigmoid_f := 349;
        ELSIF x =- 3240 THEN
            sigmoid_f := 349;
        ELSIF x =- 3239 THEN
            sigmoid_f := 349;
        ELSIF x =- 3238 THEN
            sigmoid_f := 349;
        ELSIF x =- 3237 THEN
            sigmoid_f := 349;
        ELSIF x =- 3236 THEN
            sigmoid_f := 349;
        ELSIF x =- 3235 THEN
            sigmoid_f := 350;
        ELSIF x =- 3234 THEN
            sigmoid_f := 350;
        ELSIF x =- 3233 THEN
            sigmoid_f := 350;
        ELSIF x =- 3232 THEN
            sigmoid_f := 350;
        ELSIF x =- 3231 THEN
            sigmoid_f := 350;
        ELSIF x =- 3230 THEN
            sigmoid_f := 350;
        ELSIF x =- 3229 THEN
            sigmoid_f := 350;
        ELSIF x =- 3228 THEN
            sigmoid_f := 351;
        ELSIF x =- 3227 THEN
            sigmoid_f := 351;
        ELSIF x =- 3226 THEN
            sigmoid_f := 351;
        ELSIF x =- 3225 THEN
            sigmoid_f := 351;
        ELSIF x =- 3224 THEN
            sigmoid_f := 351;
        ELSIF x =- 3223 THEN
            sigmoid_f := 351;
        ELSIF x =- 3222 THEN
            sigmoid_f := 351;
        ELSIF x =- 3221 THEN
            sigmoid_f := 352;
        ELSIF x =- 3220 THEN
            sigmoid_f := 352;
        ELSIF x =- 3219 THEN
            sigmoid_f := 352;
        ELSIF x =- 3218 THEN
            sigmoid_f := 352;
        ELSIF x =- 3217 THEN
            sigmoid_f := 352;
        ELSIF x =- 3216 THEN
            sigmoid_f := 352;
        ELSIF x =- 3215 THEN
            sigmoid_f := 352;
        ELSIF x =- 3214 THEN
            sigmoid_f := 353;
        ELSIF x =- 3213 THEN
            sigmoid_f := 353;
        ELSIF x =- 3212 THEN
            sigmoid_f := 353;
        ELSIF x =- 3211 THEN
            sigmoid_f := 353;
        ELSIF x =- 3210 THEN
            sigmoid_f := 353;
        ELSIF x =- 3209 THEN
            sigmoid_f := 353;
        ELSIF x =- 3208 THEN
            sigmoid_f := 353;
        ELSIF x =- 3207 THEN
            sigmoid_f := 353;
        ELSIF x =- 3206 THEN
            sigmoid_f := 354;
        ELSIF x =- 3205 THEN
            sigmoid_f := 354;
        ELSIF x =- 3204 THEN
            sigmoid_f := 354;
        ELSIF x =- 3203 THEN
            sigmoid_f := 354;
        ELSIF x =- 3202 THEN
            sigmoid_f := 354;
        ELSIF x =- 3201 THEN
            sigmoid_f := 354;
        ELSIF x =- 3200 THEN
            sigmoid_f := 354;
        ELSIF x =- 3199 THEN
            sigmoid_f := 355;
        ELSIF x =- 3198 THEN
            sigmoid_f := 355;
        ELSIF x =- 3197 THEN
            sigmoid_f := 355;
        ELSIF x =- 3196 THEN
            sigmoid_f := 355;
        ELSIF x =- 3195 THEN
            sigmoid_f := 355;
        ELSIF x =- 3194 THEN
            sigmoid_f := 355;
        ELSIF x =- 3193 THEN
            sigmoid_f := 355;
        ELSIF x =- 3192 THEN
            sigmoid_f := 356;
        ELSIF x =- 3191 THEN
            sigmoid_f := 356;
        ELSIF x =- 3190 THEN
            sigmoid_f := 356;
        ELSIF x =- 3189 THEN
            sigmoid_f := 356;
        ELSIF x =- 3188 THEN
            sigmoid_f := 356;
        ELSIF x =- 3187 THEN
            sigmoid_f := 356;
        ELSIF x =- 3186 THEN
            sigmoid_f := 356;
        ELSIF x =- 3185 THEN
            sigmoid_f := 356;
        ELSIF x =- 3184 THEN
            sigmoid_f := 357;
        ELSIF x =- 3183 THEN
            sigmoid_f := 357;
        ELSIF x =- 3182 THEN
            sigmoid_f := 357;
        ELSIF x =- 3181 THEN
            sigmoid_f := 357;
        ELSIF x =- 3180 THEN
            sigmoid_f := 357;
        ELSIF x =- 3179 THEN
            sigmoid_f := 357;
        ELSIF x =- 3178 THEN
            sigmoid_f := 357;
        ELSIF x =- 3177 THEN
            sigmoid_f := 358;
        ELSIF x =- 3176 THEN
            sigmoid_f := 358;
        ELSIF x =- 3175 THEN
            sigmoid_f := 358;
        ELSIF x =- 3174 THEN
            sigmoid_f := 358;
        ELSIF x =- 3173 THEN
            sigmoid_f := 358;
        ELSIF x =- 3172 THEN
            sigmoid_f := 358;
        ELSIF x =- 3171 THEN
            sigmoid_f := 358;
        ELSIF x =- 3170 THEN
            sigmoid_f := 359;
        ELSIF x =- 3169 THEN
            sigmoid_f := 359;
        ELSIF x =- 3168 THEN
            sigmoid_f := 359;
        ELSIF x =- 3167 THEN
            sigmoid_f := 359;
        ELSIF x =- 3166 THEN
            sigmoid_f := 359;
        ELSIF x =- 3165 THEN
            sigmoid_f := 359;
        ELSIF x =- 3164 THEN
            sigmoid_f := 359;
        ELSIF x =- 3163 THEN
            sigmoid_f := 360;
        ELSIF x =- 3162 THEN
            sigmoid_f := 360;
        ELSIF x =- 3161 THEN
            sigmoid_f := 360;
        ELSIF x =- 3160 THEN
            sigmoid_f := 360;
        ELSIF x =- 3159 THEN
            sigmoid_f := 360;
        ELSIF x =- 3158 THEN
            sigmoid_f := 360;
        ELSIF x =- 3157 THEN
            sigmoid_f := 360;
        ELSIF x =- 3156 THEN
            sigmoid_f := 360;
        ELSIF x =- 3155 THEN
            sigmoid_f := 361;
        ELSIF x =- 3154 THEN
            sigmoid_f := 361;
        ELSIF x =- 3153 THEN
            sigmoid_f := 361;
        ELSIF x =- 3152 THEN
            sigmoid_f := 361;
        ELSIF x =- 3151 THEN
            sigmoid_f := 361;
        ELSIF x =- 3150 THEN
            sigmoid_f := 361;
        ELSIF x =- 3149 THEN
            sigmoid_f := 361;
        ELSIF x =- 3148 THEN
            sigmoid_f := 362;
        ELSIF x =- 3147 THEN
            sigmoid_f := 362;
        ELSIF x =- 3146 THEN
            sigmoid_f := 362;
        ELSIF x =- 3145 THEN
            sigmoid_f := 362;
        ELSIF x =- 3144 THEN
            sigmoid_f := 362;
        ELSIF x =- 3143 THEN
            sigmoid_f := 362;
        ELSIF x =- 3142 THEN
            sigmoid_f := 362;
        ELSIF x =- 3141 THEN
            sigmoid_f := 363;
        ELSIF x =- 3140 THEN
            sigmoid_f := 363;
        ELSIF x =- 3139 THEN
            sigmoid_f := 363;
        ELSIF x =- 3138 THEN
            sigmoid_f := 363;
        ELSIF x =- 3137 THEN
            sigmoid_f := 363;
        ELSIF x =- 3136 THEN
            sigmoid_f := 363;
        ELSIF x =- 3135 THEN
            sigmoid_f := 363;
        ELSIF x =- 3134 THEN
            sigmoid_f := 363;
        ELSIF x =- 3133 THEN
            sigmoid_f := 364;
        ELSIF x =- 3132 THEN
            sigmoid_f := 364;
        ELSIF x =- 3131 THEN
            sigmoid_f := 364;
        ELSIF x =- 3130 THEN
            sigmoid_f := 364;
        ELSIF x =- 3129 THEN
            sigmoid_f := 364;
        ELSIF x =- 3128 THEN
            sigmoid_f := 364;
        ELSIF x =- 3127 THEN
            sigmoid_f := 364;
        ELSIF x =- 3126 THEN
            sigmoid_f := 365;
        ELSIF x =- 3125 THEN
            sigmoid_f := 365;
        ELSIF x =- 3124 THEN
            sigmoid_f := 365;
        ELSIF x =- 3123 THEN
            sigmoid_f := 365;
        ELSIF x =- 3122 THEN
            sigmoid_f := 365;
        ELSIF x =- 3121 THEN
            sigmoid_f := 365;
        ELSIF x =- 3120 THEN
            sigmoid_f := 365;
        ELSIF x =- 3119 THEN
            sigmoid_f := 366;
        ELSIF x =- 3118 THEN
            sigmoid_f := 366;
        ELSIF x =- 3117 THEN
            sigmoid_f := 366;
        ELSIF x =- 3116 THEN
            sigmoid_f := 366;
        ELSIF x =- 3115 THEN
            sigmoid_f := 366;
        ELSIF x =- 3114 THEN
            sigmoid_f := 366;
        ELSIF x =- 3113 THEN
            sigmoid_f := 366;
        ELSIF x =- 3112 THEN
            sigmoid_f := 367;
        ELSIF x =- 3111 THEN
            sigmoid_f := 367;
        ELSIF x =- 3110 THEN
            sigmoid_f := 367;
        ELSIF x =- 3109 THEN
            sigmoid_f := 367;
        ELSIF x =- 3108 THEN
            sigmoid_f := 367;
        ELSIF x =- 3107 THEN
            sigmoid_f := 367;
        ELSIF x =- 3106 THEN
            sigmoid_f := 367;
        ELSIF x =- 3105 THEN
            sigmoid_f := 367;
        ELSIF x =- 3104 THEN
            sigmoid_f := 368;
        ELSIF x =- 3103 THEN
            sigmoid_f := 368;
        ELSIF x =- 3102 THEN
            sigmoid_f := 368;
        ELSIF x =- 3101 THEN
            sigmoid_f := 368;
        ELSIF x =- 3100 THEN
            sigmoid_f := 368;
        ELSIF x =- 3099 THEN
            sigmoid_f := 368;
        ELSIF x =- 3098 THEN
            sigmoid_f := 368;
        ELSIF x =- 3097 THEN
            sigmoid_f := 369;
        ELSIF x =- 3096 THEN
            sigmoid_f := 369;
        ELSIF x =- 3095 THEN
            sigmoid_f := 369;
        ELSIF x =- 3094 THEN
            sigmoid_f := 369;
        ELSIF x =- 3093 THEN
            sigmoid_f := 369;
        ELSIF x =- 3092 THEN
            sigmoid_f := 369;
        ELSIF x =- 3091 THEN
            sigmoid_f := 369;
        ELSIF x =- 3090 THEN
            sigmoid_f := 370;
        ELSIF x =- 3089 THEN
            sigmoid_f := 370;
        ELSIF x =- 3088 THEN
            sigmoid_f := 370;
        ELSIF x =- 3087 THEN
            sigmoid_f := 370;
        ELSIF x =- 3086 THEN
            sigmoid_f := 370;
        ELSIF x =- 3085 THEN
            sigmoid_f := 370;
        ELSIF x =- 3084 THEN
            sigmoid_f := 370;
        ELSIF x =- 3083 THEN
            sigmoid_f := 370;
        ELSIF x =- 3082 THEN
            sigmoid_f := 371;
        ELSIF x =- 3081 THEN
            sigmoid_f := 371;
        ELSIF x =- 3080 THEN
            sigmoid_f := 371;
        ELSIF x =- 3079 THEN
            sigmoid_f := 371;
        ELSIF x =- 3078 THEN
            sigmoid_f := 371;
        ELSIF x =- 3077 THEN
            sigmoid_f := 371;
        ELSIF x =- 3076 THEN
            sigmoid_f := 371;
        ELSIF x =- 3075 THEN
            sigmoid_f := 372;
        ELSIF x =- 3074 THEN
            sigmoid_f := 372;
        ELSIF x =- 3073 THEN
            sigmoid_f := 372;
        ELSIF x =- 3072 THEN
            sigmoid_f := 372;
        ELSIF x =- 3071 THEN
            sigmoid_f := 372;
        ELSIF x =- 3070 THEN
            sigmoid_f := 372;
        ELSIF x =- 3069 THEN
            sigmoid_f := 372;
        ELSIF x =- 3068 THEN
            sigmoid_f := 373;
        ELSIF x =- 3067 THEN
            sigmoid_f := 373;
        ELSIF x =- 3066 THEN
            sigmoid_f := 373;
        ELSIF x =- 3065 THEN
            sigmoid_f := 373;
        ELSIF x =- 3064 THEN
            sigmoid_f := 373;
        ELSIF x =- 3063 THEN
            sigmoid_f := 373;
        ELSIF x =- 3062 THEN
            sigmoid_f := 374;
        ELSIF x =- 3061 THEN
            sigmoid_f := 374;
        ELSIF x =- 3060 THEN
            sigmoid_f := 374;
        ELSIF x =- 3059 THEN
            sigmoid_f := 374;
        ELSIF x =- 3058 THEN
            sigmoid_f := 374;
        ELSIF x =- 3057 THEN
            sigmoid_f := 374;
        ELSIF x =- 3056 THEN
            sigmoid_f := 375;
        ELSIF x =- 3055 THEN
            sigmoid_f := 375;
        ELSIF x =- 3054 THEN
            sigmoid_f := 375;
        ELSIF x =- 3053 THEN
            sigmoid_f := 375;
        ELSIF x =- 3052 THEN
            sigmoid_f := 375;
        ELSIF x =- 3051 THEN
            sigmoid_f := 375;
        ELSIF x =- 3050 THEN
            sigmoid_f := 376;
        ELSIF x =- 3049 THEN
            sigmoid_f := 376;
        ELSIF x =- 3048 THEN
            sigmoid_f := 376;
        ELSIF x =- 3047 THEN
            sigmoid_f := 376;
        ELSIF x =- 3046 THEN
            sigmoid_f := 376;
        ELSIF x =- 3045 THEN
            sigmoid_f := 376;
        ELSIF x =- 3044 THEN
            sigmoid_f := 376;
        ELSIF x =- 3043 THEN
            sigmoid_f := 377;
        ELSIF x =- 3042 THEN
            sigmoid_f := 377;
        ELSIF x =- 3041 THEN
            sigmoid_f := 377;
        ELSIF x =- 3040 THEN
            sigmoid_f := 377;
        ELSIF x =- 3039 THEN
            sigmoid_f := 377;
        ELSIF x =- 3038 THEN
            sigmoid_f := 377;
        ELSIF x =- 3037 THEN
            sigmoid_f := 378;
        ELSIF x =- 3036 THEN
            sigmoid_f := 378;
        ELSIF x =- 3035 THEN
            sigmoid_f := 378;
        ELSIF x =- 3034 THEN
            sigmoid_f := 378;
        ELSIF x =- 3033 THEN
            sigmoid_f := 378;
        ELSIF x =- 3032 THEN
            sigmoid_f := 378;
        ELSIF x =- 3031 THEN
            sigmoid_f := 379;
        ELSIF x =- 3030 THEN
            sigmoid_f := 379;
        ELSIF x =- 3029 THEN
            sigmoid_f := 379;
        ELSIF x =- 3028 THEN
            sigmoid_f := 379;
        ELSIF x =- 3027 THEN
            sigmoid_f := 379;
        ELSIF x =- 3026 THEN
            sigmoid_f := 379;
        ELSIF x =- 3025 THEN
            sigmoid_f := 380;
        ELSIF x =- 3024 THEN
            sigmoid_f := 380;
        ELSIF x =- 3023 THEN
            sigmoid_f := 380;
        ELSIF x =- 3022 THEN
            sigmoid_f := 380;
        ELSIF x =- 3021 THEN
            sigmoid_f := 380;
        ELSIF x =- 3020 THEN
            sigmoid_f := 380;
        ELSIF x =- 3019 THEN
            sigmoid_f := 381;
        ELSIF x =- 3018 THEN
            sigmoid_f := 381;
        ELSIF x =- 3017 THEN
            sigmoid_f := 381;
        ELSIF x =- 3016 THEN
            sigmoid_f := 381;
        ELSIF x =- 3015 THEN
            sigmoid_f := 381;
        ELSIF x =- 3014 THEN
            sigmoid_f := 381;
        ELSIF x =- 3013 THEN
            sigmoid_f := 381;
        ELSIF x =- 3012 THEN
            sigmoid_f := 382;
        ELSIF x =- 3011 THEN
            sigmoid_f := 382;
        ELSIF x =- 3010 THEN
            sigmoid_f := 382;
        ELSIF x =- 3009 THEN
            sigmoid_f := 382;
        ELSIF x =- 3008 THEN
            sigmoid_f := 382;
        ELSIF x =- 3007 THEN
            sigmoid_f := 382;
        ELSIF x =- 3006 THEN
            sigmoid_f := 383;
        ELSIF x =- 3005 THEN
            sigmoid_f := 383;
        ELSIF x =- 3004 THEN
            sigmoid_f := 383;
        ELSIF x =- 3003 THEN
            sigmoid_f := 383;
        ELSIF x =- 3002 THEN
            sigmoid_f := 383;
        ELSIF x =- 3001 THEN
            sigmoid_f := 383;
        ELSIF x =- 3000 THEN
            sigmoid_f := 384;
        ELSIF x =- 2999 THEN
            sigmoid_f := 384;
        ELSIF x =- 2998 THEN
            sigmoid_f := 384;
        ELSIF x =- 2997 THEN
            sigmoid_f := 384;
        ELSIF x =- 2996 THEN
            sigmoid_f := 384;
        ELSIF x =- 2995 THEN
            sigmoid_f := 384;
        ELSIF x =- 2994 THEN
            sigmoid_f := 385;
        ELSIF x =- 2993 THEN
            sigmoid_f := 385;
        ELSIF x =- 2992 THEN
            sigmoid_f := 385;
        ELSIF x =- 2991 THEN
            sigmoid_f := 385;
        ELSIF x =- 2990 THEN
            sigmoid_f := 385;
        ELSIF x =- 2989 THEN
            sigmoid_f := 385;
        ELSIF x =- 2988 THEN
            sigmoid_f := 385;
        ELSIF x =- 2987 THEN
            sigmoid_f := 386;
        ELSIF x =- 2986 THEN
            sigmoid_f := 386;
        ELSIF x =- 2985 THEN
            sigmoid_f := 386;
        ELSIF x =- 2984 THEN
            sigmoid_f := 386;
        ELSIF x =- 2983 THEN
            sigmoid_f := 386;
        ELSIF x =- 2982 THEN
            sigmoid_f := 386;
        ELSIF x =- 2981 THEN
            sigmoid_f := 387;
        ELSIF x =- 2980 THEN
            sigmoid_f := 387;
        ELSIF x =- 2979 THEN
            sigmoid_f := 387;
        ELSIF x =- 2978 THEN
            sigmoid_f := 387;
        ELSIF x =- 2977 THEN
            sigmoid_f := 387;
        ELSIF x =- 2976 THEN
            sigmoid_f := 387;
        ELSIF x =- 2975 THEN
            sigmoid_f := 388;
        ELSIF x =- 2974 THEN
            sigmoid_f := 388;
        ELSIF x =- 2973 THEN
            sigmoid_f := 388;
        ELSIF x =- 2972 THEN
            sigmoid_f := 388;
        ELSIF x =- 2971 THEN
            sigmoid_f := 388;
        ELSIF x =- 2970 THEN
            sigmoid_f := 388;
        ELSIF x =- 2969 THEN
            sigmoid_f := 389;
        ELSIF x =- 2968 THEN
            sigmoid_f := 389;
        ELSIF x =- 2967 THEN
            sigmoid_f := 389;
        ELSIF x =- 2966 THEN
            sigmoid_f := 389;
        ELSIF x =- 2965 THEN
            sigmoid_f := 389;
        ELSIF x =- 2964 THEN
            sigmoid_f := 389;
        ELSIF x =- 2963 THEN
            sigmoid_f := 390;
        ELSIF x =- 2962 THEN
            sigmoid_f := 390;
        ELSIF x =- 2961 THEN
            sigmoid_f := 390;
        ELSIF x =- 2960 THEN
            sigmoid_f := 390;
        ELSIF x =- 2959 THEN
            sigmoid_f := 390;
        ELSIF x =- 2958 THEN
            sigmoid_f := 390;
        ELSIF x =- 2957 THEN
            sigmoid_f := 390;
        ELSIF x =- 2956 THEN
            sigmoid_f := 391;
        ELSIF x =- 2955 THEN
            sigmoid_f := 391;
        ELSIF x =- 2954 THEN
            sigmoid_f := 391;
        ELSIF x =- 2953 THEN
            sigmoid_f := 391;
        ELSIF x =- 2952 THEN
            sigmoid_f := 391;
        ELSIF x =- 2951 THEN
            sigmoid_f := 391;
        ELSIF x =- 2950 THEN
            sigmoid_f := 392;
        ELSIF x =- 2949 THEN
            sigmoid_f := 392;
        ELSIF x =- 2948 THEN
            sigmoid_f := 392;
        ELSIF x =- 2947 THEN
            sigmoid_f := 392;
        ELSIF x =- 2946 THEN
            sigmoid_f := 392;
        ELSIF x =- 2945 THEN
            sigmoid_f := 392;
        ELSIF x =- 2944 THEN
            sigmoid_f := 393;
        ELSIF x =- 2943 THEN
            sigmoid_f := 393;
        ELSIF x =- 2942 THEN
            sigmoid_f := 393;
        ELSIF x =- 2941 THEN
            sigmoid_f := 393;
        ELSIF x =- 2940 THEN
            sigmoid_f := 393;
        ELSIF x =- 2939 THEN
            sigmoid_f := 393;
        ELSIF x =- 2938 THEN
            sigmoid_f := 394;
        ELSIF x =- 2937 THEN
            sigmoid_f := 394;
        ELSIF x =- 2936 THEN
            sigmoid_f := 394;
        ELSIF x =- 2935 THEN
            sigmoid_f := 394;
        ELSIF x =- 2934 THEN
            sigmoid_f := 394;
        ELSIF x =- 2933 THEN
            sigmoid_f := 394;
        ELSIF x =- 2932 THEN
            sigmoid_f := 394;
        ELSIF x =- 2931 THEN
            sigmoid_f := 395;
        ELSIF x =- 2930 THEN
            sigmoid_f := 395;
        ELSIF x =- 2929 THEN
            sigmoid_f := 395;
        ELSIF x =- 2928 THEN
            sigmoid_f := 395;
        ELSIF x =- 2927 THEN
            sigmoid_f := 395;
        ELSIF x =- 2926 THEN
            sigmoid_f := 395;
        ELSIF x =- 2925 THEN
            sigmoid_f := 396;
        ELSIF x =- 2924 THEN
            sigmoid_f := 396;
        ELSIF x =- 2923 THEN
            sigmoid_f := 396;
        ELSIF x =- 2922 THEN
            sigmoid_f := 396;
        ELSIF x =- 2921 THEN
            sigmoid_f := 396;
        ELSIF x =- 2920 THEN
            sigmoid_f := 396;
        ELSIF x =- 2919 THEN
            sigmoid_f := 397;
        ELSIF x =- 2918 THEN
            sigmoid_f := 397;
        ELSIF x =- 2917 THEN
            sigmoid_f := 397;
        ELSIF x =- 2916 THEN
            sigmoid_f := 397;
        ELSIF x =- 2915 THEN
            sigmoid_f := 397;
        ELSIF x =- 2914 THEN
            sigmoid_f := 397;
        ELSIF x =- 2913 THEN
            sigmoid_f := 398;
        ELSIF x =- 2912 THEN
            sigmoid_f := 398;
        ELSIF x =- 2911 THEN
            sigmoid_f := 398;
        ELSIF x =- 2910 THEN
            sigmoid_f := 398;
        ELSIF x =- 2909 THEN
            sigmoid_f := 398;
        ELSIF x =- 2908 THEN
            sigmoid_f := 398;
        ELSIF x =- 2907 THEN
            sigmoid_f := 399;
        ELSIF x =- 2906 THEN
            sigmoid_f := 399;
        ELSIF x =- 2905 THEN
            sigmoid_f := 399;
        ELSIF x =- 2904 THEN
            sigmoid_f := 399;
        ELSIF x =- 2903 THEN
            sigmoid_f := 399;
        ELSIF x =- 2902 THEN
            sigmoid_f := 399;
        ELSIF x =- 2901 THEN
            sigmoid_f := 399;
        ELSIF x =- 2900 THEN
            sigmoid_f := 400;
        ELSIF x =- 2899 THEN
            sigmoid_f := 400;
        ELSIF x =- 2898 THEN
            sigmoid_f := 400;
        ELSIF x =- 2897 THEN
            sigmoid_f := 400;
        ELSIF x =- 2896 THEN
            sigmoid_f := 400;
        ELSIF x =- 2895 THEN
            sigmoid_f := 400;
        ELSIF x =- 2894 THEN
            sigmoid_f := 401;
        ELSIF x =- 2893 THEN
            sigmoid_f := 401;
        ELSIF x =- 2892 THEN
            sigmoid_f := 401;
        ELSIF x =- 2891 THEN
            sigmoid_f := 401;
        ELSIF x =- 2890 THEN
            sigmoid_f := 401;
        ELSIF x =- 2889 THEN
            sigmoid_f := 401;
        ELSIF x =- 2888 THEN
            sigmoid_f := 402;
        ELSIF x =- 2887 THEN
            sigmoid_f := 402;
        ELSIF x =- 2886 THEN
            sigmoid_f := 402;
        ELSIF x =- 2885 THEN
            sigmoid_f := 402;
        ELSIF x =- 2884 THEN
            sigmoid_f := 402;
        ELSIF x =- 2883 THEN
            sigmoid_f := 402;
        ELSIF x =- 2882 THEN
            sigmoid_f := 403;
        ELSIF x =- 2881 THEN
            sigmoid_f := 403;
        ELSIF x =- 2880 THEN
            sigmoid_f := 403;
        ELSIF x =- 2879 THEN
            sigmoid_f := 403;
        ELSIF x =- 2878 THEN
            sigmoid_f := 403;
        ELSIF x =- 2877 THEN
            sigmoid_f := 403;
        ELSIF x =- 2876 THEN
            sigmoid_f := 403;
        ELSIF x =- 2875 THEN
            sigmoid_f := 404;
        ELSIF x =- 2874 THEN
            sigmoid_f := 404;
        ELSIF x =- 2873 THEN
            sigmoid_f := 404;
        ELSIF x =- 2872 THEN
            sigmoid_f := 404;
        ELSIF x =- 2871 THEN
            sigmoid_f := 404;
        ELSIF x =- 2870 THEN
            sigmoid_f := 404;
        ELSIF x =- 2869 THEN
            sigmoid_f := 405;
        ELSIF x =- 2868 THEN
            sigmoid_f := 405;
        ELSIF x =- 2867 THEN
            sigmoid_f := 405;
        ELSIF x =- 2866 THEN
            sigmoid_f := 405;
        ELSIF x =- 2865 THEN
            sigmoid_f := 405;
        ELSIF x =- 2864 THEN
            sigmoid_f := 405;
        ELSIF x =- 2863 THEN
            sigmoid_f := 406;
        ELSIF x =- 2862 THEN
            sigmoid_f := 406;
        ELSIF x =- 2861 THEN
            sigmoid_f := 406;
        ELSIF x =- 2860 THEN
            sigmoid_f := 406;
        ELSIF x =- 2859 THEN
            sigmoid_f := 406;
        ELSIF x =- 2858 THEN
            sigmoid_f := 406;
        ELSIF x =- 2857 THEN
            sigmoid_f := 407;
        ELSIF x =- 2856 THEN
            sigmoid_f := 407;
        ELSIF x =- 2855 THEN
            sigmoid_f := 407;
        ELSIF x =- 2854 THEN
            sigmoid_f := 407;
        ELSIF x =- 2853 THEN
            sigmoid_f := 407;
        ELSIF x =- 2852 THEN
            sigmoid_f := 407;
        ELSIF x =- 2851 THEN
            sigmoid_f := 408;
        ELSIF x =- 2850 THEN
            sigmoid_f := 408;
        ELSIF x =- 2849 THEN
            sigmoid_f := 408;
        ELSIF x =- 2848 THEN
            sigmoid_f := 408;
        ELSIF x =- 2847 THEN
            sigmoid_f := 408;
        ELSIF x =- 2846 THEN
            sigmoid_f := 408;
        ELSIF x =- 2845 THEN
            sigmoid_f := 408;
        ELSIF x =- 2844 THEN
            sigmoid_f := 409;
        ELSIF x =- 2843 THEN
            sigmoid_f := 409;
        ELSIF x =- 2842 THEN
            sigmoid_f := 409;
        ELSIF x =- 2841 THEN
            sigmoid_f := 409;
        ELSIF x =- 2840 THEN
            sigmoid_f := 409;
        ELSIF x =- 2839 THEN
            sigmoid_f := 409;
        ELSIF x =- 2838 THEN
            sigmoid_f := 410;
        ELSIF x =- 2837 THEN
            sigmoid_f := 410;
        ELSIF x =- 2836 THEN
            sigmoid_f := 410;
        ELSIF x =- 2835 THEN
            sigmoid_f := 410;
        ELSIF x =- 2834 THEN
            sigmoid_f := 410;
        ELSIF x =- 2833 THEN
            sigmoid_f := 410;
        ELSIF x =- 2832 THEN
            sigmoid_f := 411;
        ELSIF x =- 2831 THEN
            sigmoid_f := 411;
        ELSIF x =- 2830 THEN
            sigmoid_f := 411;
        ELSIF x =- 2829 THEN
            sigmoid_f := 411;
        ELSIF x =- 2828 THEN
            sigmoid_f := 411;
        ELSIF x =- 2827 THEN
            sigmoid_f := 411;
        ELSIF x =- 2826 THEN
            sigmoid_f := 412;
        ELSIF x =- 2825 THEN
            sigmoid_f := 412;
        ELSIF x =- 2824 THEN
            sigmoid_f := 412;
        ELSIF x =- 2823 THEN
            sigmoid_f := 412;
        ELSIF x =- 2822 THEN
            sigmoid_f := 412;
        ELSIF x =- 2821 THEN
            sigmoid_f := 412;
        ELSIF x =- 2820 THEN
            sigmoid_f := 412;
        ELSIF x =- 2819 THEN
            sigmoid_f := 413;
        ELSIF x =- 2818 THEN
            sigmoid_f := 413;
        ELSIF x =- 2817 THEN
            sigmoid_f := 413;
        ELSIF x =- 2816 THEN
            sigmoid_f := 413;
        ELSIF x =- 2815 THEN
            sigmoid_f := 413;
        ELSIF x =- 2814 THEN
            sigmoid_f := 413;
        ELSIF x =- 2813 THEN
            sigmoid_f := 414;
        ELSIF x =- 2812 THEN
            sigmoid_f := 414;
        ELSIF x =- 2811 THEN
            sigmoid_f := 414;
        ELSIF x =- 2810 THEN
            sigmoid_f := 414;
        ELSIF x =- 2809 THEN
            sigmoid_f := 414;
        ELSIF x =- 2808 THEN
            sigmoid_f := 414;
        ELSIF x =- 2807 THEN
            sigmoid_f := 415;
        ELSIF x =- 2806 THEN
            sigmoid_f := 415;
        ELSIF x =- 2805 THEN
            sigmoid_f := 415;
        ELSIF x =- 2804 THEN
            sigmoid_f := 415;
        ELSIF x =- 2803 THEN
            sigmoid_f := 415;
        ELSIF x =- 2802 THEN
            sigmoid_f := 415;
        ELSIF x =- 2801 THEN
            sigmoid_f := 416;
        ELSIF x =- 2800 THEN
            sigmoid_f := 416;
        ELSIF x =- 2799 THEN
            sigmoid_f := 416;
        ELSIF x =- 2798 THEN
            sigmoid_f := 416;
        ELSIF x =- 2797 THEN
            sigmoid_f := 416;
        ELSIF x =- 2796 THEN
            sigmoid_f := 416;
        ELSIF x =- 2795 THEN
            sigmoid_f := 416;
        ELSIF x =- 2794 THEN
            sigmoid_f := 417;
        ELSIF x =- 2793 THEN
            sigmoid_f := 417;
        ELSIF x =- 2792 THEN
            sigmoid_f := 417;
        ELSIF x =- 2791 THEN
            sigmoid_f := 417;
        ELSIF x =- 2790 THEN
            sigmoid_f := 417;
        ELSIF x =- 2789 THEN
            sigmoid_f := 417;
        ELSIF x =- 2788 THEN
            sigmoid_f := 418;
        ELSIF x =- 2787 THEN
            sigmoid_f := 418;
        ELSIF x =- 2786 THEN
            sigmoid_f := 418;
        ELSIF x =- 2785 THEN
            sigmoid_f := 418;
        ELSIF x =- 2784 THEN
            sigmoid_f := 418;
        ELSIF x =- 2783 THEN
            sigmoid_f := 418;
        ELSIF x =- 2782 THEN
            sigmoid_f := 419;
        ELSIF x =- 2781 THEN
            sigmoid_f := 419;
        ELSIF x =- 2780 THEN
            sigmoid_f := 419;
        ELSIF x =- 2779 THEN
            sigmoid_f := 419;
        ELSIF x =- 2778 THEN
            sigmoid_f := 419;
        ELSIF x =- 2777 THEN
            sigmoid_f := 419;
        ELSIF x =- 2776 THEN
            sigmoid_f := 420;
        ELSIF x =- 2775 THEN
            sigmoid_f := 420;
        ELSIF x =- 2774 THEN
            sigmoid_f := 420;
        ELSIF x =- 2773 THEN
            sigmoid_f := 420;
        ELSIF x =- 2772 THEN
            sigmoid_f := 420;
        ELSIF x =- 2771 THEN
            sigmoid_f := 420;
        ELSIF x =- 2770 THEN
            sigmoid_f := 421;
        ELSIF x =- 2769 THEN
            sigmoid_f := 421;
        ELSIF x =- 2768 THEN
            sigmoid_f := 421;
        ELSIF x =- 2767 THEN
            sigmoid_f := 421;
        ELSIF x =- 2766 THEN
            sigmoid_f := 421;
        ELSIF x =- 2765 THEN
            sigmoid_f := 421;
        ELSIF x =- 2764 THEN
            sigmoid_f := 421;
        ELSIF x =- 2763 THEN
            sigmoid_f := 422;
        ELSIF x =- 2762 THEN
            sigmoid_f := 422;
        ELSIF x =- 2761 THEN
            sigmoid_f := 422;
        ELSIF x =- 2760 THEN
            sigmoid_f := 422;
        ELSIF x =- 2759 THEN
            sigmoid_f := 422;
        ELSIF x =- 2758 THEN
            sigmoid_f := 422;
        ELSIF x =- 2757 THEN
            sigmoid_f := 423;
        ELSIF x =- 2756 THEN
            sigmoid_f := 423;
        ELSIF x =- 2755 THEN
            sigmoid_f := 423;
        ELSIF x =- 2754 THEN
            sigmoid_f := 423;
        ELSIF x =- 2753 THEN
            sigmoid_f := 423;
        ELSIF x =- 2752 THEN
            sigmoid_f := 423;
        ELSIF x =- 2751 THEN
            sigmoid_f := 424;
        ELSIF x =- 2750 THEN
            sigmoid_f := 424;
        ELSIF x =- 2749 THEN
            sigmoid_f := 424;
        ELSIF x =- 2748 THEN
            sigmoid_f := 424;
        ELSIF x =- 2747 THEN
            sigmoid_f := 424;
        ELSIF x =- 2746 THEN
            sigmoid_f := 424;
        ELSIF x =- 2745 THEN
            sigmoid_f := 425;
        ELSIF x =- 2744 THEN
            sigmoid_f := 425;
        ELSIF x =- 2743 THEN
            sigmoid_f := 425;
        ELSIF x =- 2742 THEN
            sigmoid_f := 425;
        ELSIF x =- 2741 THEN
            sigmoid_f := 425;
        ELSIF x =- 2740 THEN
            sigmoid_f := 425;
        ELSIF x =- 2739 THEN
            sigmoid_f := 425;
        ELSIF x =- 2738 THEN
            sigmoid_f := 426;
        ELSIF x =- 2737 THEN
            sigmoid_f := 426;
        ELSIF x =- 2736 THEN
            sigmoid_f := 426;
        ELSIF x =- 2735 THEN
            sigmoid_f := 426;
        ELSIF x =- 2734 THEN
            sigmoid_f := 426;
        ELSIF x =- 2733 THEN
            sigmoid_f := 426;
        ELSIF x =- 2732 THEN
            sigmoid_f := 427;
        ELSIF x =- 2731 THEN
            sigmoid_f := 427;
        ELSIF x =- 2730 THEN
            sigmoid_f := 427;
        ELSIF x =- 2729 THEN
            sigmoid_f := 427;
        ELSIF x =- 2728 THEN
            sigmoid_f := 427;
        ELSIF x =- 2727 THEN
            sigmoid_f := 427;
        ELSIF x =- 2726 THEN
            sigmoid_f := 428;
        ELSIF x =- 2725 THEN
            sigmoid_f := 428;
        ELSIF x =- 2724 THEN
            sigmoid_f := 428;
        ELSIF x =- 2723 THEN
            sigmoid_f := 428;
        ELSIF x =- 2722 THEN
            sigmoid_f := 428;
        ELSIF x =- 2721 THEN
            sigmoid_f := 428;
        ELSIF x =- 2720 THEN
            sigmoid_f := 429;
        ELSIF x =- 2719 THEN
            sigmoid_f := 429;
        ELSIF x =- 2718 THEN
            sigmoid_f := 429;
        ELSIF x =- 2717 THEN
            sigmoid_f := 429;
        ELSIF x =- 2716 THEN
            sigmoid_f := 429;
        ELSIF x =- 2715 THEN
            sigmoid_f := 429;
        ELSIF x =- 2714 THEN
            sigmoid_f := 430;
        ELSIF x =- 2713 THEN
            sigmoid_f := 430;
        ELSIF x =- 2712 THEN
            sigmoid_f := 430;
        ELSIF x =- 2711 THEN
            sigmoid_f := 430;
        ELSIF x =- 2710 THEN
            sigmoid_f := 430;
        ELSIF x =- 2709 THEN
            sigmoid_f := 430;
        ELSIF x =- 2708 THEN
            sigmoid_f := 430;
        ELSIF x =- 2707 THEN
            sigmoid_f := 431;
        ELSIF x =- 2706 THEN
            sigmoid_f := 431;
        ELSIF x =- 2705 THEN
            sigmoid_f := 431;
        ELSIF x =- 2704 THEN
            sigmoid_f := 431;
        ELSIF x =- 2703 THEN
            sigmoid_f := 431;
        ELSIF x =- 2702 THEN
            sigmoid_f := 431;
        ELSIF x =- 2701 THEN
            sigmoid_f := 432;
        ELSIF x =- 2700 THEN
            sigmoid_f := 432;
        ELSIF x =- 2699 THEN
            sigmoid_f := 432;
        ELSIF x =- 2698 THEN
            sigmoid_f := 432;
        ELSIF x =- 2697 THEN
            sigmoid_f := 432;
        ELSIF x =- 2696 THEN
            sigmoid_f := 432;
        ELSIF x =- 2695 THEN
            sigmoid_f := 433;
        ELSIF x =- 2694 THEN
            sigmoid_f := 433;
        ELSIF x =- 2693 THEN
            sigmoid_f := 433;
        ELSIF x =- 2692 THEN
            sigmoid_f := 433;
        ELSIF x =- 2691 THEN
            sigmoid_f := 433;
        ELSIF x =- 2690 THEN
            sigmoid_f := 433;
        ELSIF x =- 2689 THEN
            sigmoid_f := 434;
        ELSIF x =- 2688 THEN
            sigmoid_f := 434;
        ELSIF x =- 2687 THEN
            sigmoid_f := 434;
        ELSIF x =- 2686 THEN
            sigmoid_f := 434;
        ELSIF x =- 2685 THEN
            sigmoid_f := 434;
        ELSIF x =- 2684 THEN
            sigmoid_f := 434;
        ELSIF x =- 2683 THEN
            sigmoid_f := 434;
        ELSIF x =- 2682 THEN
            sigmoid_f := 435;
        ELSIF x =- 2681 THEN
            sigmoid_f := 435;
        ELSIF x =- 2680 THEN
            sigmoid_f := 435;
        ELSIF x =- 2679 THEN
            sigmoid_f := 435;
        ELSIF x =- 2678 THEN
            sigmoid_f := 435;
        ELSIF x =- 2677 THEN
            sigmoid_f := 435;
        ELSIF x =- 2676 THEN
            sigmoid_f := 436;
        ELSIF x =- 2675 THEN
            sigmoid_f := 436;
        ELSIF x =- 2674 THEN
            sigmoid_f := 436;
        ELSIF x =- 2673 THEN
            sigmoid_f := 436;
        ELSIF x =- 2672 THEN
            sigmoid_f := 436;
        ELSIF x =- 2671 THEN
            sigmoid_f := 436;
        ELSIF x =- 2670 THEN
            sigmoid_f := 437;
        ELSIF x =- 2669 THEN
            sigmoid_f := 437;
        ELSIF x =- 2668 THEN
            sigmoid_f := 437;
        ELSIF x =- 2667 THEN
            sigmoid_f := 437;
        ELSIF x =- 2666 THEN
            sigmoid_f := 437;
        ELSIF x =- 2665 THEN
            sigmoid_f := 437;
        ELSIF x =- 2664 THEN
            sigmoid_f := 438;
        ELSIF x =- 2663 THEN
            sigmoid_f := 438;
        ELSIF x =- 2662 THEN
            sigmoid_f := 438;
        ELSIF x =- 2661 THEN
            sigmoid_f := 438;
        ELSIF x =- 2660 THEN
            sigmoid_f := 438;
        ELSIF x =- 2659 THEN
            sigmoid_f := 438;
        ELSIF x =- 2658 THEN
            sigmoid_f := 439;
        ELSIF x =- 2657 THEN
            sigmoid_f := 439;
        ELSIF x =- 2656 THEN
            sigmoid_f := 439;
        ELSIF x =- 2655 THEN
            sigmoid_f := 439;
        ELSIF x =- 2654 THEN
            sigmoid_f := 439;
        ELSIF x =- 2653 THEN
            sigmoid_f := 439;
        ELSIF x =- 2652 THEN
            sigmoid_f := 439;
        ELSIF x =- 2651 THEN
            sigmoid_f := 440;
        ELSIF x =- 2650 THEN
            sigmoid_f := 440;
        ELSIF x =- 2649 THEN
            sigmoid_f := 440;
        ELSIF x =- 2648 THEN
            sigmoid_f := 440;
        ELSIF x =- 2647 THEN
            sigmoid_f := 440;
        ELSIF x =- 2646 THEN
            sigmoid_f := 440;
        ELSIF x =- 2645 THEN
            sigmoid_f := 441;
        ELSIF x =- 2644 THEN
            sigmoid_f := 441;
        ELSIF x =- 2643 THEN
            sigmoid_f := 441;
        ELSIF x =- 2642 THEN
            sigmoid_f := 441;
        ELSIF x =- 2641 THEN
            sigmoid_f := 441;
        ELSIF x =- 2640 THEN
            sigmoid_f := 441;
        ELSIF x =- 2639 THEN
            sigmoid_f := 442;
        ELSIF x =- 2638 THEN
            sigmoid_f := 442;
        ELSIF x =- 2637 THEN
            sigmoid_f := 442;
        ELSIF x =- 2636 THEN
            sigmoid_f := 442;
        ELSIF x =- 2635 THEN
            sigmoid_f := 442;
        ELSIF x =- 2634 THEN
            sigmoid_f := 442;
        ELSIF x =- 2633 THEN
            sigmoid_f := 443;
        ELSIF x =- 2632 THEN
            sigmoid_f := 443;
        ELSIF x =- 2631 THEN
            sigmoid_f := 443;
        ELSIF x =- 2630 THEN
            sigmoid_f := 443;
        ELSIF x =- 2629 THEN
            sigmoid_f := 443;
        ELSIF x =- 2628 THEN
            sigmoid_f := 443;
        ELSIF x =- 2627 THEN
            sigmoid_f := 443;
        ELSIF x =- 2626 THEN
            sigmoid_f := 444;
        ELSIF x =- 2625 THEN
            sigmoid_f := 444;
        ELSIF x =- 2624 THEN
            sigmoid_f := 444;
        ELSIF x =- 2623 THEN
            sigmoid_f := 444;
        ELSIF x =- 2622 THEN
            sigmoid_f := 444;
        ELSIF x =- 2621 THEN
            sigmoid_f := 444;
        ELSIF x =- 2620 THEN
            sigmoid_f := 445;
        ELSIF x =- 2619 THEN
            sigmoid_f := 445;
        ELSIF x =- 2618 THEN
            sigmoid_f := 445;
        ELSIF x =- 2617 THEN
            sigmoid_f := 445;
        ELSIF x =- 2616 THEN
            sigmoid_f := 445;
        ELSIF x =- 2615 THEN
            sigmoid_f := 445;
        ELSIF x =- 2614 THEN
            sigmoid_f := 446;
        ELSIF x =- 2613 THEN
            sigmoid_f := 446;
        ELSIF x =- 2612 THEN
            sigmoid_f := 446;
        ELSIF x =- 2611 THEN
            sigmoid_f := 446;
        ELSIF x =- 2610 THEN
            sigmoid_f := 446;
        ELSIF x =- 2609 THEN
            sigmoid_f := 446;
        ELSIF x =- 2608 THEN
            sigmoid_f := 447;
        ELSIF x =- 2607 THEN
            sigmoid_f := 447;
        ELSIF x =- 2606 THEN
            sigmoid_f := 447;
        ELSIF x =- 2605 THEN
            sigmoid_f := 447;
        ELSIF x =- 2604 THEN
            sigmoid_f := 447;
        ELSIF x =- 2603 THEN
            sigmoid_f := 447;
        ELSIF x =- 2602 THEN
            sigmoid_f := 448;
        ELSIF x =- 2601 THEN
            sigmoid_f := 448;
        ELSIF x =- 2600 THEN
            sigmoid_f := 448;
        ELSIF x =- 2599 THEN
            sigmoid_f := 448;
        ELSIF x =- 2598 THEN
            sigmoid_f := 448;
        ELSIF x =- 2597 THEN
            sigmoid_f := 448;
        ELSIF x =- 2596 THEN
            sigmoid_f := 448;
        ELSIF x =- 2595 THEN
            sigmoid_f := 449;
        ELSIF x =- 2594 THEN
            sigmoid_f := 449;
        ELSIF x =- 2593 THEN
            sigmoid_f := 449;
        ELSIF x =- 2592 THEN
            sigmoid_f := 449;
        ELSIF x =- 2591 THEN
            sigmoid_f := 449;
        ELSIF x =- 2590 THEN
            sigmoid_f := 449;
        ELSIF x =- 2589 THEN
            sigmoid_f := 450;
        ELSIF x =- 2588 THEN
            sigmoid_f := 450;
        ELSIF x =- 2587 THEN
            sigmoid_f := 450;
        ELSIF x =- 2586 THEN
            sigmoid_f := 450;
        ELSIF x =- 2585 THEN
            sigmoid_f := 450;
        ELSIF x =- 2584 THEN
            sigmoid_f := 450;
        ELSIF x =- 2583 THEN
            sigmoid_f := 451;
        ELSIF x =- 2582 THEN
            sigmoid_f := 451;
        ELSIF x =- 2581 THEN
            sigmoid_f := 451;
        ELSIF x =- 2580 THEN
            sigmoid_f := 451;
        ELSIF x =- 2579 THEN
            sigmoid_f := 451;
        ELSIF x =- 2578 THEN
            sigmoid_f := 451;
        ELSIF x =- 2577 THEN
            sigmoid_f := 452;
        ELSIF x =- 2576 THEN
            sigmoid_f := 452;
        ELSIF x =- 2575 THEN
            sigmoid_f := 452;
        ELSIF x =- 2574 THEN
            sigmoid_f := 452;
        ELSIF x =- 2573 THEN
            sigmoid_f := 452;
        ELSIF x =- 2572 THEN
            sigmoid_f := 452;
        ELSIF x =- 2571 THEN
            sigmoid_f := 452;
        ELSIF x =- 2570 THEN
            sigmoid_f := 453;
        ELSIF x =- 2569 THEN
            sigmoid_f := 453;
        ELSIF x =- 2568 THEN
            sigmoid_f := 453;
        ELSIF x =- 2567 THEN
            sigmoid_f := 453;
        ELSIF x =- 2566 THEN
            sigmoid_f := 453;
        ELSIF x =- 2565 THEN
            sigmoid_f := 453;
        ELSIF x =- 2564 THEN
            sigmoid_f := 454;
        ELSIF x =- 2563 THEN
            sigmoid_f := 454;
        ELSIF x =- 2562 THEN
            sigmoid_f := 454;
        ELSIF x =- 2561 THEN
            sigmoid_f := 454;
        ELSIF x =- 2560 THEN
            sigmoid_f := 454;
        ELSIF x =- 2559 THEN
            sigmoid_f := 454;
        ELSIF x =- 2558 THEN
            sigmoid_f := 455;
        ELSIF x =- 2557 THEN
            sigmoid_f := 455;
        ELSIF x =- 2556 THEN
            sigmoid_f := 455;
        ELSIF x =- 2555 THEN
            sigmoid_f := 455;
        ELSIF x =- 2554 THEN
            sigmoid_f := 455;
        ELSIF x =- 2553 THEN
            sigmoid_f := 456;
        ELSIF x =- 2552 THEN
            sigmoid_f := 456;
        ELSIF x =- 2551 THEN
            sigmoid_f := 456;
        ELSIF x =- 2550 THEN
            sigmoid_f := 456;
        ELSIF x =- 2549 THEN
            sigmoid_f := 456;
        ELSIF x =- 2548 THEN
            sigmoid_f := 456;
        ELSIF x =- 2547 THEN
            sigmoid_f := 457;
        ELSIF x =- 2546 THEN
            sigmoid_f := 457;
        ELSIF x =- 2545 THEN
            sigmoid_f := 457;
        ELSIF x =- 2544 THEN
            sigmoid_f := 457;
        ELSIF x =- 2543 THEN
            sigmoid_f := 457;
        ELSIF x =- 2542 THEN
            sigmoid_f := 458;
        ELSIF x =- 2541 THEN
            sigmoid_f := 458;
        ELSIF x =- 2540 THEN
            sigmoid_f := 458;
        ELSIF x =- 2539 THEN
            sigmoid_f := 458;
        ELSIF x =- 2538 THEN
            sigmoid_f := 458;
        ELSIF x =- 2537 THEN
            sigmoid_f := 459;
        ELSIF x =- 2536 THEN
            sigmoid_f := 459;
        ELSIF x =- 2535 THEN
            sigmoid_f := 459;
        ELSIF x =- 2534 THEN
            sigmoid_f := 459;
        ELSIF x =- 2533 THEN
            sigmoid_f := 459;
        ELSIF x =- 2532 THEN
            sigmoid_f := 459;
        ELSIF x =- 2531 THEN
            sigmoid_f := 460;
        ELSIF x =- 2530 THEN
            sigmoid_f := 460;
        ELSIF x =- 2529 THEN
            sigmoid_f := 460;
        ELSIF x =- 2528 THEN
            sigmoid_f := 460;
        ELSIF x =- 2527 THEN
            sigmoid_f := 460;
        ELSIF x =- 2526 THEN
            sigmoid_f := 461;
        ELSIF x =- 2525 THEN
            sigmoid_f := 461;
        ELSIF x =- 2524 THEN
            sigmoid_f := 461;
        ELSIF x =- 2523 THEN
            sigmoid_f := 461;
        ELSIF x =- 2522 THEN
            sigmoid_f := 461;
        ELSIF x =- 2521 THEN
            sigmoid_f := 462;
        ELSIF x =- 2520 THEN
            sigmoid_f := 462;
        ELSIF x =- 2519 THEN
            sigmoid_f := 462;
        ELSIF x =- 2518 THEN
            sigmoid_f := 462;
        ELSIF x =- 2517 THEN
            sigmoid_f := 462;
        ELSIF x =- 2516 THEN
            sigmoid_f := 462;
        ELSIF x =- 2515 THEN
            sigmoid_f := 463;
        ELSIF x =- 2514 THEN
            sigmoid_f := 463;
        ELSIF x =- 2513 THEN
            sigmoid_f := 463;
        ELSIF x =- 2512 THEN
            sigmoid_f := 463;
        ELSIF x =- 2511 THEN
            sigmoid_f := 463;
        ELSIF x =- 2510 THEN
            sigmoid_f := 464;
        ELSIF x =- 2509 THEN
            sigmoid_f := 464;
        ELSIF x =- 2508 THEN
            sigmoid_f := 464;
        ELSIF x =- 2507 THEN
            sigmoid_f := 464;
        ELSIF x =- 2506 THEN
            sigmoid_f := 464;
        ELSIF x =- 2505 THEN
            sigmoid_f := 464;
        ELSIF x =- 2504 THEN
            sigmoid_f := 465;
        ELSIF x =- 2503 THEN
            sigmoid_f := 465;
        ELSIF x =- 2502 THEN
            sigmoid_f := 465;
        ELSIF x =- 2501 THEN
            sigmoid_f := 465;
        ELSIF x =- 2500 THEN
            sigmoid_f := 465;
        ELSIF x =- 2499 THEN
            sigmoid_f := 466;
        ELSIF x =- 2498 THEN
            sigmoid_f := 466;
        ELSIF x =- 2497 THEN
            sigmoid_f := 466;
        ELSIF x =- 2496 THEN
            sigmoid_f := 466;
        ELSIF x =- 2495 THEN
            sigmoid_f := 466;
        ELSIF x =- 2494 THEN
            sigmoid_f := 467;
        ELSIF x =- 2493 THEN
            sigmoid_f := 467;
        ELSIF x =- 2492 THEN
            sigmoid_f := 467;
        ELSIF x =- 2491 THEN
            sigmoid_f := 467;
        ELSIF x =- 2490 THEN
            sigmoid_f := 467;
        ELSIF x =- 2489 THEN
            sigmoid_f := 467;
        ELSIF x =- 2488 THEN
            sigmoid_f := 468;
        ELSIF x =- 2487 THEN
            sigmoid_f := 468;
        ELSIF x =- 2486 THEN
            sigmoid_f := 468;
        ELSIF x =- 2485 THEN
            sigmoid_f := 468;
        ELSIF x =- 2484 THEN
            sigmoid_f := 468;
        ELSIF x =- 2483 THEN
            sigmoid_f := 469;
        ELSIF x =- 2482 THEN
            sigmoid_f := 469;
        ELSIF x =- 2481 THEN
            sigmoid_f := 469;
        ELSIF x =- 2480 THEN
            sigmoid_f := 469;
        ELSIF x =- 2479 THEN
            sigmoid_f := 469;
        ELSIF x =- 2478 THEN
            sigmoid_f := 470;
        ELSIF x =- 2477 THEN
            sigmoid_f := 470;
        ELSIF x =- 2476 THEN
            sigmoid_f := 470;
        ELSIF x =- 2475 THEN
            sigmoid_f := 470;
        ELSIF x =- 2474 THEN
            sigmoid_f := 470;
        ELSIF x =- 2473 THEN
            sigmoid_f := 470;
        ELSIF x =- 2472 THEN
            sigmoid_f := 471;
        ELSIF x =- 2471 THEN
            sigmoid_f := 471;
        ELSIF x =- 2470 THEN
            sigmoid_f := 471;
        ELSIF x =- 2469 THEN
            sigmoid_f := 471;
        ELSIF x =- 2468 THEN
            sigmoid_f := 471;
        ELSIF x =- 2467 THEN
            sigmoid_f := 472;
        ELSIF x =- 2466 THEN
            sigmoid_f := 472;
        ELSIF x =- 2465 THEN
            sigmoid_f := 472;
        ELSIF x =- 2464 THEN
            sigmoid_f := 472;
        ELSIF x =- 2463 THEN
            sigmoid_f := 472;
        ELSIF x =- 2462 THEN
            sigmoid_f := 472;
        ELSIF x =- 2461 THEN
            sigmoid_f := 473;
        ELSIF x =- 2460 THEN
            sigmoid_f := 473;
        ELSIF x =- 2459 THEN
            sigmoid_f := 473;
        ELSIF x =- 2458 THEN
            sigmoid_f := 473;
        ELSIF x =- 2457 THEN
            sigmoid_f := 473;
        ELSIF x =- 2456 THEN
            sigmoid_f := 474;
        ELSIF x =- 2455 THEN
            sigmoid_f := 474;
        ELSIF x =- 2454 THEN
            sigmoid_f := 474;
        ELSIF x =- 2453 THEN
            sigmoid_f := 474;
        ELSIF x =- 2452 THEN
            sigmoid_f := 474;
        ELSIF x =- 2451 THEN
            sigmoid_f := 475;
        ELSIF x =- 2450 THEN
            sigmoid_f := 475;
        ELSIF x =- 2449 THEN
            sigmoid_f := 475;
        ELSIF x =- 2448 THEN
            sigmoid_f := 475;
        ELSIF x =- 2447 THEN
            sigmoid_f := 475;
        ELSIF x =- 2446 THEN
            sigmoid_f := 475;
        ELSIF x =- 2445 THEN
            sigmoid_f := 476;
        ELSIF x =- 2444 THEN
            sigmoid_f := 476;
        ELSIF x =- 2443 THEN
            sigmoid_f := 476;
        ELSIF x =- 2442 THEN
            sigmoid_f := 476;
        ELSIF x =- 2441 THEN
            sigmoid_f := 476;
        ELSIF x =- 2440 THEN
            sigmoid_f := 477;
        ELSIF x =- 2439 THEN
            sigmoid_f := 477;
        ELSIF x =- 2438 THEN
            sigmoid_f := 477;
        ELSIF x =- 2437 THEN
            sigmoid_f := 477;
        ELSIF x =- 2436 THEN
            sigmoid_f := 477;
        ELSIF x =- 2435 THEN
            sigmoid_f := 478;
        ELSIF x =- 2434 THEN
            sigmoid_f := 478;
        ELSIF x =- 2433 THEN
            sigmoid_f := 478;
        ELSIF x =- 2432 THEN
            sigmoid_f := 478;
        ELSIF x =- 2431 THEN
            sigmoid_f := 478;
        ELSIF x =- 2430 THEN
            sigmoid_f := 478;
        ELSIF x =- 2429 THEN
            sigmoid_f := 479;
        ELSIF x =- 2428 THEN
            sigmoid_f := 479;
        ELSIF x =- 2427 THEN
            sigmoid_f := 479;
        ELSIF x =- 2426 THEN
            sigmoid_f := 479;
        ELSIF x =- 2425 THEN
            sigmoid_f := 479;
        ELSIF x =- 2424 THEN
            sigmoid_f := 480;
        ELSIF x =- 2423 THEN
            sigmoid_f := 480;
        ELSIF x =- 2422 THEN
            sigmoid_f := 480;
        ELSIF x =- 2421 THEN
            sigmoid_f := 480;
        ELSIF x =- 2420 THEN
            sigmoid_f := 480;
        ELSIF x =- 2419 THEN
            sigmoid_f := 480;
        ELSIF x =- 2418 THEN
            sigmoid_f := 481;
        ELSIF x =- 2417 THEN
            sigmoid_f := 481;
        ELSIF x =- 2416 THEN
            sigmoid_f := 481;
        ELSIF x =- 2415 THEN
            sigmoid_f := 481;
        ELSIF x =- 2414 THEN
            sigmoid_f := 481;
        ELSIF x =- 2413 THEN
            sigmoid_f := 482;
        ELSIF x =- 2412 THEN
            sigmoid_f := 482;
        ELSIF x =- 2411 THEN
            sigmoid_f := 482;
        ELSIF x =- 2410 THEN
            sigmoid_f := 482;
        ELSIF x =- 2409 THEN
            sigmoid_f := 482;
        ELSIF x =- 2408 THEN
            sigmoid_f := 483;
        ELSIF x =- 2407 THEN
            sigmoid_f := 483;
        ELSIF x =- 2406 THEN
            sigmoid_f := 483;
        ELSIF x =- 2405 THEN
            sigmoid_f := 483;
        ELSIF x =- 2404 THEN
            sigmoid_f := 483;
        ELSIF x =- 2403 THEN
            sigmoid_f := 483;
        ELSIF x =- 2402 THEN
            sigmoid_f := 484;
        ELSIF x =- 2401 THEN
            sigmoid_f := 484;
        ELSIF x =- 2400 THEN
            sigmoid_f := 484;
        ELSIF x =- 2399 THEN
            sigmoid_f := 484;
        ELSIF x =- 2398 THEN
            sigmoid_f := 484;
        ELSIF x =- 2397 THEN
            sigmoid_f := 485;
        ELSIF x =- 2396 THEN
            sigmoid_f := 485;
        ELSIF x =- 2395 THEN
            sigmoid_f := 485;
        ELSIF x =- 2394 THEN
            sigmoid_f := 485;
        ELSIF x =- 2393 THEN
            sigmoid_f := 485;
        ELSIF x =- 2392 THEN
            sigmoid_f := 486;
        ELSIF x =- 2391 THEN
            sigmoid_f := 486;
        ELSIF x =- 2390 THEN
            sigmoid_f := 486;
        ELSIF x =- 2389 THEN
            sigmoid_f := 486;
        ELSIF x =- 2388 THEN
            sigmoid_f := 486;
        ELSIF x =- 2387 THEN
            sigmoid_f := 486;
        ELSIF x =- 2386 THEN
            sigmoid_f := 487;
        ELSIF x =- 2385 THEN
            sigmoid_f := 487;
        ELSIF x =- 2384 THEN
            sigmoid_f := 487;
        ELSIF x =- 2383 THEN
            sigmoid_f := 487;
        ELSIF x =- 2382 THEN
            sigmoid_f := 487;
        ELSIF x =- 2381 THEN
            sigmoid_f := 488;
        ELSIF x =- 2380 THEN
            sigmoid_f := 488;
        ELSIF x =- 2379 THEN
            sigmoid_f := 488;
        ELSIF x =- 2378 THEN
            sigmoid_f := 488;
        ELSIF x =- 2377 THEN
            sigmoid_f := 488;
        ELSIF x =- 2376 THEN
            sigmoid_f := 488;
        ELSIF x =- 2375 THEN
            sigmoid_f := 489;
        ELSIF x =- 2374 THEN
            sigmoid_f := 489;
        ELSIF x =- 2373 THEN
            sigmoid_f := 489;
        ELSIF x =- 2372 THEN
            sigmoid_f := 489;
        ELSIF x =- 2371 THEN
            sigmoid_f := 489;
        ELSIF x =- 2370 THEN
            sigmoid_f := 490;
        ELSIF x =- 2369 THEN
            sigmoid_f := 490;
        ELSIF x =- 2368 THEN
            sigmoid_f := 490;
        ELSIF x =- 2367 THEN
            sigmoid_f := 490;
        ELSIF x =- 2366 THEN
            sigmoid_f := 490;
        ELSIF x =- 2365 THEN
            sigmoid_f := 491;
        ELSIF x =- 2364 THEN
            sigmoid_f := 491;
        ELSIF x =- 2363 THEN
            sigmoid_f := 491;
        ELSIF x =- 2362 THEN
            sigmoid_f := 491;
        ELSIF x =- 2361 THEN
            sigmoid_f := 491;
        ELSIF x =- 2360 THEN
            sigmoid_f := 491;
        ELSIF x =- 2359 THEN
            sigmoid_f := 492;
        ELSIF x =- 2358 THEN
            sigmoid_f := 492;
        ELSIF x =- 2357 THEN
            sigmoid_f := 492;
        ELSIF x =- 2356 THEN
            sigmoid_f := 492;
        ELSIF x =- 2355 THEN
            sigmoid_f := 492;
        ELSIF x =- 2354 THEN
            sigmoid_f := 493;
        ELSIF x =- 2353 THEN
            sigmoid_f := 493;
        ELSIF x =- 2352 THEN
            sigmoid_f := 493;
        ELSIF x =- 2351 THEN
            sigmoid_f := 493;
        ELSIF x =- 2350 THEN
            sigmoid_f := 493;
        ELSIF x =- 2349 THEN
            sigmoid_f := 494;
        ELSIF x =- 2348 THEN
            sigmoid_f := 494;
        ELSIF x =- 2347 THEN
            sigmoid_f := 494;
        ELSIF x =- 2346 THEN
            sigmoid_f := 494;
        ELSIF x =- 2345 THEN
            sigmoid_f := 494;
        ELSIF x =- 2344 THEN
            sigmoid_f := 494;
        ELSIF x =- 2343 THEN
            sigmoid_f := 495;
        ELSIF x =- 2342 THEN
            sigmoid_f := 495;
        ELSIF x =- 2341 THEN
            sigmoid_f := 495;
        ELSIF x =- 2340 THEN
            sigmoid_f := 495;
        ELSIF x =- 2339 THEN
            sigmoid_f := 495;
        ELSIF x =- 2338 THEN
            sigmoid_f := 496;
        ELSIF x =- 2337 THEN
            sigmoid_f := 496;
        ELSIF x =- 2336 THEN
            sigmoid_f := 496;
        ELSIF x =- 2335 THEN
            sigmoid_f := 496;
        ELSIF x =- 2334 THEN
            sigmoid_f := 496;
        ELSIF x =- 2333 THEN
            sigmoid_f := 496;
        ELSIF x =- 2332 THEN
            sigmoid_f := 497;
        ELSIF x =- 2331 THEN
            sigmoid_f := 497;
        ELSIF x =- 2330 THEN
            sigmoid_f := 497;
        ELSIF x =- 2329 THEN
            sigmoid_f := 497;
        ELSIF x =- 2328 THEN
            sigmoid_f := 497;
        ELSIF x =- 2327 THEN
            sigmoid_f := 498;
        ELSIF x =- 2326 THEN
            sigmoid_f := 498;
        ELSIF x =- 2325 THEN
            sigmoid_f := 498;
        ELSIF x =- 2324 THEN
            sigmoid_f := 498;
        ELSIF x =- 2323 THEN
            sigmoid_f := 498;
        ELSIF x =- 2322 THEN
            sigmoid_f := 499;
        ELSIF x =- 2321 THEN
            sigmoid_f := 499;
        ELSIF x =- 2320 THEN
            sigmoid_f := 499;
        ELSIF x =- 2319 THEN
            sigmoid_f := 499;
        ELSIF x =- 2318 THEN
            sigmoid_f := 499;
        ELSIF x =- 2317 THEN
            sigmoid_f := 499;
        ELSIF x =- 2316 THEN
            sigmoid_f := 500;
        ELSIF x =- 2315 THEN
            sigmoid_f := 500;
        ELSIF x =- 2314 THEN
            sigmoid_f := 500;
        ELSIF x =- 2313 THEN
            sigmoid_f := 500;
        ELSIF x =- 2312 THEN
            sigmoid_f := 500;
        ELSIF x =- 2311 THEN
            sigmoid_f := 501;
        ELSIF x =- 2310 THEN
            sigmoid_f := 501;
        ELSIF x =- 2309 THEN
            sigmoid_f := 501;
        ELSIF x =- 2308 THEN
            sigmoid_f := 501;
        ELSIF x =- 2307 THEN
            sigmoid_f := 501;
        ELSIF x =- 2306 THEN
            sigmoid_f := 502;
        ELSIF x =- 2305 THEN
            sigmoid_f := 502;
        ELSIF x =- 2304 THEN
            sigmoid_f := 502;
        ELSIF x =- 2303 THEN
            sigmoid_f := 502;
        ELSIF x =- 2302 THEN
            sigmoid_f := 502;
        ELSIF x =- 2301 THEN
            sigmoid_f := 502;
        ELSIF x =- 2300 THEN
            sigmoid_f := 503;
        ELSIF x =- 2299 THEN
            sigmoid_f := 503;
        ELSIF x =- 2298 THEN
            sigmoid_f := 503;
        ELSIF x =- 2297 THEN
            sigmoid_f := 503;
        ELSIF x =- 2296 THEN
            sigmoid_f := 503;
        ELSIF x =- 2295 THEN
            sigmoid_f := 504;
        ELSIF x =- 2294 THEN
            sigmoid_f := 504;
        ELSIF x =- 2293 THEN
            sigmoid_f := 504;
        ELSIF x =- 2292 THEN
            sigmoid_f := 504;
        ELSIF x =- 2291 THEN
            sigmoid_f := 504;
        ELSIF x =- 2290 THEN
            sigmoid_f := 504;
        ELSIF x =- 2289 THEN
            sigmoid_f := 505;
        ELSIF x =- 2288 THEN
            sigmoid_f := 505;
        ELSIF x =- 2287 THEN
            sigmoid_f := 505;
        ELSIF x =- 2286 THEN
            sigmoid_f := 505;
        ELSIF x =- 2285 THEN
            sigmoid_f := 505;
        ELSIF x =- 2284 THEN
            sigmoid_f := 506;
        ELSIF x =- 2283 THEN
            sigmoid_f := 506;
        ELSIF x =- 2282 THEN
            sigmoid_f := 506;
        ELSIF x =- 2281 THEN
            sigmoid_f := 506;
        ELSIF x =- 2280 THEN
            sigmoid_f := 506;
        ELSIF x =- 2279 THEN
            sigmoid_f := 507;
        ELSIF x =- 2278 THEN
            sigmoid_f := 507;
        ELSIF x =- 2277 THEN
            sigmoid_f := 507;
        ELSIF x =- 2276 THEN
            sigmoid_f := 507;
        ELSIF x =- 2275 THEN
            sigmoid_f := 507;
        ELSIF x =- 2274 THEN
            sigmoid_f := 507;
        ELSIF x =- 2273 THEN
            sigmoid_f := 508;
        ELSIF x =- 2272 THEN
            sigmoid_f := 508;
        ELSIF x =- 2271 THEN
            sigmoid_f := 508;
        ELSIF x =- 2270 THEN
            sigmoid_f := 508;
        ELSIF x =- 2269 THEN
            sigmoid_f := 508;
        ELSIF x =- 2268 THEN
            sigmoid_f := 509;
        ELSIF x =- 2267 THEN
            sigmoid_f := 509;
        ELSIF x =- 2266 THEN
            sigmoid_f := 509;
        ELSIF x =- 2265 THEN
            sigmoid_f := 509;
        ELSIF x =- 2264 THEN
            sigmoid_f := 509;
        ELSIF x =- 2263 THEN
            sigmoid_f := 510;
        ELSIF x =- 2262 THEN
            sigmoid_f := 510;
        ELSIF x =- 2261 THEN
            sigmoid_f := 510;
        ELSIF x =- 2260 THEN
            sigmoid_f := 510;
        ELSIF x =- 2259 THEN
            sigmoid_f := 510;
        ELSIF x =- 2258 THEN
            sigmoid_f := 510;
        ELSIF x =- 2257 THEN
            sigmoid_f := 511;
        ELSIF x =- 2256 THEN
            sigmoid_f := 511;
        ELSIF x =- 2255 THEN
            sigmoid_f := 511;
        ELSIF x =- 2254 THEN
            sigmoid_f := 511;
        ELSIF x =- 2253 THEN
            sigmoid_f := 511;
        ELSIF x =- 2252 THEN
            sigmoid_f := 512;
        ELSIF x =- 2251 THEN
            sigmoid_f := 512;
        ELSIF x =- 2250 THEN
            sigmoid_f := 512;
        ELSIF x =- 2249 THEN
            sigmoid_f := 512;
        ELSIF x =- 2248 THEN
            sigmoid_f := 512;
        ELSIF x =- 2247 THEN
            sigmoid_f := 512;
        ELSIF x =- 2246 THEN
            sigmoid_f := 513;
        ELSIF x =- 2245 THEN
            sigmoid_f := 513;
        ELSIF x =- 2244 THEN
            sigmoid_f := 513;
        ELSIF x =- 2243 THEN
            sigmoid_f := 513;
        ELSIF x =- 2242 THEN
            sigmoid_f := 513;
        ELSIF x =- 2241 THEN
            sigmoid_f := 514;
        ELSIF x =- 2240 THEN
            sigmoid_f := 514;
        ELSIF x =- 2239 THEN
            sigmoid_f := 514;
        ELSIF x =- 2238 THEN
            sigmoid_f := 514;
        ELSIF x =- 2237 THEN
            sigmoid_f := 514;
        ELSIF x =- 2236 THEN
            sigmoid_f := 515;
        ELSIF x =- 2235 THEN
            sigmoid_f := 515;
        ELSIF x =- 2234 THEN
            sigmoid_f := 515;
        ELSIF x =- 2233 THEN
            sigmoid_f := 515;
        ELSIF x =- 2232 THEN
            sigmoid_f := 515;
        ELSIF x =- 2231 THEN
            sigmoid_f := 515;
        ELSIF x =- 2230 THEN
            sigmoid_f := 516;
        ELSIF x =- 2229 THEN
            sigmoid_f := 516;
        ELSIF x =- 2228 THEN
            sigmoid_f := 516;
        ELSIF x =- 2227 THEN
            sigmoid_f := 516;
        ELSIF x =- 2226 THEN
            sigmoid_f := 516;
        ELSIF x =- 2225 THEN
            sigmoid_f := 517;
        ELSIF x =- 2224 THEN
            sigmoid_f := 517;
        ELSIF x =- 2223 THEN
            sigmoid_f := 517;
        ELSIF x =- 2222 THEN
            sigmoid_f := 517;
        ELSIF x =- 2221 THEN
            sigmoid_f := 517;
        ELSIF x =- 2220 THEN
            sigmoid_f := 518;
        ELSIF x =- 2219 THEN
            sigmoid_f := 518;
        ELSIF x =- 2218 THEN
            sigmoid_f := 518;
        ELSIF x =- 2217 THEN
            sigmoid_f := 518;
        ELSIF x =- 2216 THEN
            sigmoid_f := 518;
        ELSIF x =- 2215 THEN
            sigmoid_f := 518;
        ELSIF x =- 2214 THEN
            sigmoid_f := 519;
        ELSIF x =- 2213 THEN
            sigmoid_f := 519;
        ELSIF x =- 2212 THEN
            sigmoid_f := 519;
        ELSIF x =- 2211 THEN
            sigmoid_f := 519;
        ELSIF x =- 2210 THEN
            sigmoid_f := 519;
        ELSIF x =- 2209 THEN
            sigmoid_f := 520;
        ELSIF x =- 2208 THEN
            sigmoid_f := 520;
        ELSIF x =- 2207 THEN
            sigmoid_f := 520;
        ELSIF x =- 2206 THEN
            sigmoid_f := 520;
        ELSIF x =- 2205 THEN
            sigmoid_f := 520;
        ELSIF x =- 2204 THEN
            sigmoid_f := 520;
        ELSIF x =- 2203 THEN
            sigmoid_f := 521;
        ELSIF x =- 2202 THEN
            sigmoid_f := 521;
        ELSIF x =- 2201 THEN
            sigmoid_f := 521;
        ELSIF x =- 2200 THEN
            sigmoid_f := 521;
        ELSIF x =- 2199 THEN
            sigmoid_f := 521;
        ELSIF x =- 2198 THEN
            sigmoid_f := 522;
        ELSIF x =- 2197 THEN
            sigmoid_f := 522;
        ELSIF x =- 2196 THEN
            sigmoid_f := 522;
        ELSIF x =- 2195 THEN
            sigmoid_f := 522;
        ELSIF x =- 2194 THEN
            sigmoid_f := 522;
        ELSIF x =- 2193 THEN
            sigmoid_f := 523;
        ELSIF x =- 2192 THEN
            sigmoid_f := 523;
        ELSIF x =- 2191 THEN
            sigmoid_f := 523;
        ELSIF x =- 2190 THEN
            sigmoid_f := 523;
        ELSIF x =- 2189 THEN
            sigmoid_f := 523;
        ELSIF x =- 2188 THEN
            sigmoid_f := 523;
        ELSIF x =- 2187 THEN
            sigmoid_f := 524;
        ELSIF x =- 2186 THEN
            sigmoid_f := 524;
        ELSIF x =- 2185 THEN
            sigmoid_f := 524;
        ELSIF x =- 2184 THEN
            sigmoid_f := 524;
        ELSIF x =- 2183 THEN
            sigmoid_f := 524;
        ELSIF x =- 2182 THEN
            sigmoid_f := 525;
        ELSIF x =- 2181 THEN
            sigmoid_f := 525;
        ELSIF x =- 2180 THEN
            sigmoid_f := 525;
        ELSIF x =- 2179 THEN
            sigmoid_f := 525;
        ELSIF x =- 2178 THEN
            sigmoid_f := 525;
        ELSIF x =- 2177 THEN
            sigmoid_f := 526;
        ELSIF x =- 2176 THEN
            sigmoid_f := 526;
        ELSIF x =- 2175 THEN
            sigmoid_f := 526;
        ELSIF x =- 2174 THEN
            sigmoid_f := 526;
        ELSIF x =- 2173 THEN
            sigmoid_f := 526;
        ELSIF x =- 2172 THEN
            sigmoid_f := 526;
        ELSIF x =- 2171 THEN
            sigmoid_f := 527;
        ELSIF x =- 2170 THEN
            sigmoid_f := 527;
        ELSIF x =- 2169 THEN
            sigmoid_f := 527;
        ELSIF x =- 2168 THEN
            sigmoid_f := 527;
        ELSIF x =- 2167 THEN
            sigmoid_f := 527;
        ELSIF x =- 2166 THEN
            sigmoid_f := 528;
        ELSIF x =- 2165 THEN
            sigmoid_f := 528;
        ELSIF x =- 2164 THEN
            sigmoid_f := 528;
        ELSIF x =- 2163 THEN
            sigmoid_f := 528;
        ELSIF x =- 2162 THEN
            sigmoid_f := 528;
        ELSIF x =- 2161 THEN
            sigmoid_f := 528;
        ELSIF x =- 2160 THEN
            sigmoid_f := 529;
        ELSIF x =- 2159 THEN
            sigmoid_f := 529;
        ELSIF x =- 2158 THEN
            sigmoid_f := 529;
        ELSIF x =- 2157 THEN
            sigmoid_f := 529;
        ELSIF x =- 2156 THEN
            sigmoid_f := 529;
        ELSIF x =- 2155 THEN
            sigmoid_f := 530;
        ELSIF x =- 2154 THEN
            sigmoid_f := 530;
        ELSIF x =- 2153 THEN
            sigmoid_f := 530;
        ELSIF x =- 2152 THEN
            sigmoid_f := 530;
        ELSIF x =- 2151 THEN
            sigmoid_f := 530;
        ELSIF x =- 2150 THEN
            sigmoid_f := 531;
        ELSIF x =- 2149 THEN
            sigmoid_f := 531;
        ELSIF x =- 2148 THEN
            sigmoid_f := 531;
        ELSIF x =- 2147 THEN
            sigmoid_f := 531;
        ELSIF x =- 2146 THEN
            sigmoid_f := 531;
        ELSIF x =- 2145 THEN
            sigmoid_f := 531;
        ELSIF x =- 2144 THEN
            sigmoid_f := 532;
        ELSIF x =- 2143 THEN
            sigmoid_f := 532;
        ELSIF x =- 2142 THEN
            sigmoid_f := 532;
        ELSIF x =- 2141 THEN
            sigmoid_f := 532;
        ELSIF x =- 2140 THEN
            sigmoid_f := 532;
        ELSIF x =- 2139 THEN
            sigmoid_f := 533;
        ELSIF x =- 2138 THEN
            sigmoid_f := 533;
        ELSIF x =- 2137 THEN
            sigmoid_f := 533;
        ELSIF x =- 2136 THEN
            sigmoid_f := 533;
        ELSIF x =- 2135 THEN
            sigmoid_f := 533;
        ELSIF x =- 2134 THEN
            sigmoid_f := 534;
        ELSIF x =- 2133 THEN
            sigmoid_f := 534;
        ELSIF x =- 2132 THEN
            sigmoid_f := 534;
        ELSIF x =- 2131 THEN
            sigmoid_f := 534;
        ELSIF x =- 2130 THEN
            sigmoid_f := 534;
        ELSIF x =- 2129 THEN
            sigmoid_f := 534;
        ELSIF x =- 2128 THEN
            sigmoid_f := 535;
        ELSIF x =- 2127 THEN
            sigmoid_f := 535;
        ELSIF x =- 2126 THEN
            sigmoid_f := 535;
        ELSIF x =- 2125 THEN
            sigmoid_f := 535;
        ELSIF x =- 2124 THEN
            sigmoid_f := 535;
        ELSIF x =- 2123 THEN
            sigmoid_f := 536;
        ELSIF x =- 2122 THEN
            sigmoid_f := 536;
        ELSIF x =- 2121 THEN
            sigmoid_f := 536;
        ELSIF x =- 2120 THEN
            sigmoid_f := 536;
        ELSIF x =- 2119 THEN
            sigmoid_f := 536;
        ELSIF x =- 2118 THEN
            sigmoid_f := 536;
        ELSIF x =- 2117 THEN
            sigmoid_f := 537;
        ELSIF x =- 2116 THEN
            sigmoid_f := 537;
        ELSIF x =- 2115 THEN
            sigmoid_f := 537;
        ELSIF x =- 2114 THEN
            sigmoid_f := 537;
        ELSIF x =- 2113 THEN
            sigmoid_f := 537;
        ELSIF x =- 2112 THEN
            sigmoid_f := 538;
        ELSIF x =- 2111 THEN
            sigmoid_f := 538;
        ELSIF x =- 2110 THEN
            sigmoid_f := 538;
        ELSIF x =- 2109 THEN
            sigmoid_f := 538;
        ELSIF x =- 2108 THEN
            sigmoid_f := 538;
        ELSIF x =- 2107 THEN
            sigmoid_f := 539;
        ELSIF x =- 2106 THEN
            sigmoid_f := 539;
        ELSIF x =- 2105 THEN
            sigmoid_f := 539;
        ELSIF x =- 2104 THEN
            sigmoid_f := 539;
        ELSIF x =- 2103 THEN
            sigmoid_f := 539;
        ELSIF x =- 2102 THEN
            sigmoid_f := 539;
        ELSIF x =- 2101 THEN
            sigmoid_f := 540;
        ELSIF x =- 2100 THEN
            sigmoid_f := 540;
        ELSIF x =- 2099 THEN
            sigmoid_f := 540;
        ELSIF x =- 2098 THEN
            sigmoid_f := 540;
        ELSIF x =- 2097 THEN
            sigmoid_f := 540;
        ELSIF x =- 2096 THEN
            sigmoid_f := 541;
        ELSIF x =- 2095 THEN
            sigmoid_f := 541;
        ELSIF x =- 2094 THEN
            sigmoid_f := 541;
        ELSIF x =- 2093 THEN
            sigmoid_f := 541;
        ELSIF x =- 2092 THEN
            sigmoid_f := 541;
        ELSIF x =- 2091 THEN
            sigmoid_f := 542;
        ELSIF x =- 2090 THEN
            sigmoid_f := 542;
        ELSIF x =- 2089 THEN
            sigmoid_f := 542;
        ELSIF x =- 2088 THEN
            sigmoid_f := 542;
        ELSIF x =- 2087 THEN
            sigmoid_f := 542;
        ELSIF x =- 2086 THEN
            sigmoid_f := 542;
        ELSIF x =- 2085 THEN
            sigmoid_f := 543;
        ELSIF x =- 2084 THEN
            sigmoid_f := 543;
        ELSIF x =- 2083 THEN
            sigmoid_f := 543;
        ELSIF x =- 2082 THEN
            sigmoid_f := 543;
        ELSIF x =- 2081 THEN
            sigmoid_f := 543;
        ELSIF x =- 2080 THEN
            sigmoid_f := 544;
        ELSIF x =- 2079 THEN
            sigmoid_f := 544;
        ELSIF x =- 2078 THEN
            sigmoid_f := 544;
        ELSIF x =- 2077 THEN
            sigmoid_f := 544;
        ELSIF x =- 2076 THEN
            sigmoid_f := 544;
        ELSIF x =- 2075 THEN
            sigmoid_f := 544;
        ELSIF x =- 2074 THEN
            sigmoid_f := 545;
        ELSIF x =- 2073 THEN
            sigmoid_f := 545;
        ELSIF x =- 2072 THEN
            sigmoid_f := 545;
        ELSIF x =- 2071 THEN
            sigmoid_f := 545;
        ELSIF x =- 2070 THEN
            sigmoid_f := 545;
        ELSIF x =- 2069 THEN
            sigmoid_f := 546;
        ELSIF x =- 2068 THEN
            sigmoid_f := 546;
        ELSIF x =- 2067 THEN
            sigmoid_f := 546;
        ELSIF x =- 2066 THEN
            sigmoid_f := 546;
        ELSIF x =- 2065 THEN
            sigmoid_f := 546;
        ELSIF x =- 2064 THEN
            sigmoid_f := 547;
        ELSIF x =- 2063 THEN
            sigmoid_f := 547;
        ELSIF x =- 2062 THEN
            sigmoid_f := 547;
        ELSIF x =- 2061 THEN
            sigmoid_f := 547;
        ELSIF x =- 2060 THEN
            sigmoid_f := 547;
        ELSIF x =- 2059 THEN
            sigmoid_f := 547;
        ELSIF x =- 2058 THEN
            sigmoid_f := 548;
        ELSIF x =- 2057 THEN
            sigmoid_f := 548;
        ELSIF x =- 2056 THEN
            sigmoid_f := 548;
        ELSIF x =- 2055 THEN
            sigmoid_f := 548;
        ELSIF x =- 2054 THEN
            sigmoid_f := 548;
        ELSIF x =- 2053 THEN
            sigmoid_f := 549;
        ELSIF x =- 2052 THEN
            sigmoid_f := 549;
        ELSIF x =- 2051 THEN
            sigmoid_f := 549;
        ELSIF x =- 2050 THEN
            sigmoid_f := 549;
        ELSIF x =- 2049 THEN
            sigmoid_f := 549;
        ELSIF x =- 2048 THEN
            sigmoid_f := 550;
        ELSIF x =- 2047 THEN
            sigmoid_f := 550;
        ELSIF x =- 2046 THEN
            sigmoid_f := 550;
        ELSIF x =- 2045 THEN
            sigmoid_f := 550;
        ELSIF x =- 2044 THEN
            sigmoid_f := 550;
        ELSIF x =- 2043 THEN
            sigmoid_f := 551;
        ELSIF x =- 2042 THEN
            sigmoid_f := 551;
        ELSIF x =- 2041 THEN
            sigmoid_f := 551;
        ELSIF x =- 2040 THEN
            sigmoid_f := 551;
        ELSIF x =- 2039 THEN
            sigmoid_f := 551;
        ELSIF x =- 2038 THEN
            sigmoid_f := 552;
        ELSIF x =- 2037 THEN
            sigmoid_f := 552;
        ELSIF x =- 2036 THEN
            sigmoid_f := 552;
        ELSIF x =- 2035 THEN
            sigmoid_f := 552;
        ELSIF x =- 2034 THEN
            sigmoid_f := 552;
        ELSIF x =- 2033 THEN
            sigmoid_f := 553;
        ELSIF x =- 2032 THEN
            sigmoid_f := 553;
        ELSIF x =- 2031 THEN
            sigmoid_f := 553;
        ELSIF x =- 2030 THEN
            sigmoid_f := 553;
        ELSIF x =- 2029 THEN
            sigmoid_f := 553;
        ELSIF x =- 2028 THEN
            sigmoid_f := 554;
        ELSIF x =- 2027 THEN
            sigmoid_f := 554;
        ELSIF x =- 2026 THEN
            sigmoid_f := 554;
        ELSIF x =- 2025 THEN
            sigmoid_f := 554;
        ELSIF x =- 2024 THEN
            sigmoid_f := 554;
        ELSIF x =- 2023 THEN
            sigmoid_f := 555;
        ELSIF x =- 2022 THEN
            sigmoid_f := 555;
        ELSIF x =- 2021 THEN
            sigmoid_f := 555;
        ELSIF x =- 2020 THEN
            sigmoid_f := 555;
        ELSIF x =- 2019 THEN
            sigmoid_f := 556;
        ELSIF x =- 2018 THEN
            sigmoid_f := 556;
        ELSIF x =- 2017 THEN
            sigmoid_f := 556;
        ELSIF x =- 2016 THEN
            sigmoid_f := 556;
        ELSIF x =- 2015 THEN
            sigmoid_f := 556;
        ELSIF x =- 2014 THEN
            sigmoid_f := 557;
        ELSIF x =- 2013 THEN
            sigmoid_f := 557;
        ELSIF x =- 2012 THEN
            sigmoid_f := 557;
        ELSIF x =- 2011 THEN
            sigmoid_f := 557;
        ELSIF x =- 2010 THEN
            sigmoid_f := 557;
        ELSIF x =- 2009 THEN
            sigmoid_f := 558;
        ELSIF x =- 2008 THEN
            sigmoid_f := 558;
        ELSIF x =- 2007 THEN
            sigmoid_f := 558;
        ELSIF x =- 2006 THEN
            sigmoid_f := 558;
        ELSIF x =- 2005 THEN
            sigmoid_f := 558;
        ELSIF x =- 2004 THEN
            sigmoid_f := 559;
        ELSIF x =- 2003 THEN
            sigmoid_f := 559;
        ELSIF x =- 2002 THEN
            sigmoid_f := 559;
        ELSIF x =- 2001 THEN
            sigmoid_f := 559;
        ELSIF x =- 2000 THEN
            sigmoid_f := 559;
        ELSIF x =- 1999 THEN
            sigmoid_f := 560;
        ELSIF x =- 1998 THEN
            sigmoid_f := 560;
        ELSIF x =- 1997 THEN
            sigmoid_f := 560;
        ELSIF x =- 1996 THEN
            sigmoid_f := 560;
        ELSIF x =- 1995 THEN
            sigmoid_f := 560;
        ELSIF x =- 1994 THEN
            sigmoid_f := 561;
        ELSIF x =- 1993 THEN
            sigmoid_f := 561;
        ELSIF x =- 1992 THEN
            sigmoid_f := 561;
        ELSIF x =- 1991 THEN
            sigmoid_f := 561;
        ELSIF x =- 1990 THEN
            sigmoid_f := 562;
        ELSIF x =- 1989 THEN
            sigmoid_f := 562;
        ELSIF x =- 1988 THEN
            sigmoid_f := 562;
        ELSIF x =- 1987 THEN
            sigmoid_f := 562;
        ELSIF x =- 1986 THEN
            sigmoid_f := 562;
        ELSIF x =- 1985 THEN
            sigmoid_f := 563;
        ELSIF x =- 1984 THEN
            sigmoid_f := 563;
        ELSIF x =- 1983 THEN
            sigmoid_f := 563;
        ELSIF x =- 1982 THEN
            sigmoid_f := 563;
        ELSIF x =- 1981 THEN
            sigmoid_f := 563;
        ELSIF x =- 1980 THEN
            sigmoid_f := 564;
        ELSIF x =- 1979 THEN
            sigmoid_f := 564;
        ELSIF x =- 1978 THEN
            sigmoid_f := 564;
        ELSIF x =- 1977 THEN
            sigmoid_f := 564;
        ELSIF x =- 1976 THEN
            sigmoid_f := 564;
        ELSIF x =- 1975 THEN
            sigmoid_f := 565;
        ELSIF x =- 1974 THEN
            sigmoid_f := 565;
        ELSIF x =- 1973 THEN
            sigmoid_f := 565;
        ELSIF x =- 1972 THEN
            sigmoid_f := 565;
        ELSIF x =- 1971 THEN
            sigmoid_f := 565;
        ELSIF x =- 1970 THEN
            sigmoid_f := 566;
        ELSIF x =- 1969 THEN
            sigmoid_f := 566;
        ELSIF x =- 1968 THEN
            sigmoid_f := 566;
        ELSIF x =- 1967 THEN
            sigmoid_f := 566;
        ELSIF x =- 1966 THEN
            sigmoid_f := 566;
        ELSIF x =- 1965 THEN
            sigmoid_f := 567;
        ELSIF x =- 1964 THEN
            sigmoid_f := 567;
        ELSIF x =- 1963 THEN
            sigmoid_f := 567;
        ELSIF x =- 1962 THEN
            sigmoid_f := 567;
        ELSIF x =- 1961 THEN
            sigmoid_f := 568;
        ELSIF x =- 1960 THEN
            sigmoid_f := 568;
        ELSIF x =- 1959 THEN
            sigmoid_f := 568;
        ELSIF x =- 1958 THEN
            sigmoid_f := 568;
        ELSIF x =- 1957 THEN
            sigmoid_f := 568;
        ELSIF x =- 1956 THEN
            sigmoid_f := 569;
        ELSIF x =- 1955 THEN
            sigmoid_f := 569;
        ELSIF x =- 1954 THEN
            sigmoid_f := 569;
        ELSIF x =- 1953 THEN
            sigmoid_f := 569;
        ELSIF x =- 1952 THEN
            sigmoid_f := 569;
        ELSIF x =- 1951 THEN
            sigmoid_f := 570;
        ELSIF x =- 1950 THEN
            sigmoid_f := 570;
        ELSIF x =- 1949 THEN
            sigmoid_f := 570;
        ELSIF x =- 1948 THEN
            sigmoid_f := 570;
        ELSIF x =- 1947 THEN
            sigmoid_f := 570;
        ELSIF x =- 1946 THEN
            sigmoid_f := 571;
        ELSIF x =- 1945 THEN
            sigmoid_f := 571;
        ELSIF x =- 1944 THEN
            sigmoid_f := 571;
        ELSIF x =- 1943 THEN
            sigmoid_f := 571;
        ELSIF x =- 1942 THEN
            sigmoid_f := 571;
        ELSIF x =- 1941 THEN
            sigmoid_f := 572;
        ELSIF x =- 1940 THEN
            sigmoid_f := 572;
        ELSIF x =- 1939 THEN
            sigmoid_f := 572;
        ELSIF x =- 1938 THEN
            sigmoid_f := 572;
        ELSIF x =- 1937 THEN
            sigmoid_f := 572;
        ELSIF x =- 1936 THEN
            sigmoid_f := 573;
        ELSIF x =- 1935 THEN
            sigmoid_f := 573;
        ELSIF x =- 1934 THEN
            sigmoid_f := 573;
        ELSIF x =- 1933 THEN
            sigmoid_f := 573;
        ELSIF x =- 1932 THEN
            sigmoid_f := 574;
        ELSIF x =- 1931 THEN
            sigmoid_f := 574;
        ELSIF x =- 1930 THEN
            sigmoid_f := 574;
        ELSIF x =- 1929 THEN
            sigmoid_f := 574;
        ELSIF x =- 1928 THEN
            sigmoid_f := 574;
        ELSIF x =- 1927 THEN
            sigmoid_f := 575;
        ELSIF x =- 1926 THEN
            sigmoid_f := 575;
        ELSIF x =- 1925 THEN
            sigmoid_f := 575;
        ELSIF x =- 1924 THEN
            sigmoid_f := 575;
        ELSIF x =- 1923 THEN
            sigmoid_f := 575;
        ELSIF x =- 1922 THEN
            sigmoid_f := 576;
        ELSIF x =- 1921 THEN
            sigmoid_f := 576;
        ELSIF x =- 1920 THEN
            sigmoid_f := 576;
        ELSIF x =- 1919 THEN
            sigmoid_f := 576;
        ELSIF x =- 1918 THEN
            sigmoid_f := 576;
        ELSIF x =- 1917 THEN
            sigmoid_f := 577;
        ELSIF x =- 1916 THEN
            sigmoid_f := 577;
        ELSIF x =- 1915 THEN
            sigmoid_f := 577;
        ELSIF x =- 1914 THEN
            sigmoid_f := 577;
        ELSIF x =- 1913 THEN
            sigmoid_f := 577;
        ELSIF x =- 1912 THEN
            sigmoid_f := 578;
        ELSIF x =- 1911 THEN
            sigmoid_f := 578;
        ELSIF x =- 1910 THEN
            sigmoid_f := 578;
        ELSIF x =- 1909 THEN
            sigmoid_f := 578;
        ELSIF x =- 1908 THEN
            sigmoid_f := 578;
        ELSIF x =- 1907 THEN
            sigmoid_f := 579;
        ELSIF x =- 1906 THEN
            sigmoid_f := 579;
        ELSIF x =- 1905 THEN
            sigmoid_f := 579;
        ELSIF x =- 1904 THEN
            sigmoid_f := 579;
        ELSIF x =- 1903 THEN
            sigmoid_f := 580;
        ELSIF x =- 1902 THEN
            sigmoid_f := 580;
        ELSIF x =- 1901 THEN
            sigmoid_f := 580;
        ELSIF x =- 1900 THEN
            sigmoid_f := 580;
        ELSIF x =- 1899 THEN
            sigmoid_f := 580;
        ELSIF x =- 1898 THEN
            sigmoid_f := 581;
        ELSIF x =- 1897 THEN
            sigmoid_f := 581;
        ELSIF x =- 1896 THEN
            sigmoid_f := 581;
        ELSIF x =- 1895 THEN
            sigmoid_f := 581;
        ELSIF x =- 1894 THEN
            sigmoid_f := 581;
        ELSIF x =- 1893 THEN
            sigmoid_f := 582;
        ELSIF x =- 1892 THEN
            sigmoid_f := 582;
        ELSIF x =- 1891 THEN
            sigmoid_f := 582;
        ELSIF x =- 1890 THEN
            sigmoid_f := 582;
        ELSIF x =- 1889 THEN
            sigmoid_f := 582;
        ELSIF x =- 1888 THEN
            sigmoid_f := 583;
        ELSIF x =- 1887 THEN
            sigmoid_f := 583;
        ELSIF x =- 1886 THEN
            sigmoid_f := 583;
        ELSIF x =- 1885 THEN
            sigmoid_f := 583;
        ELSIF x =- 1884 THEN
            sigmoid_f := 583;
        ELSIF x =- 1883 THEN
            sigmoid_f := 584;
        ELSIF x =- 1882 THEN
            sigmoid_f := 584;
        ELSIF x =- 1881 THEN
            sigmoid_f := 584;
        ELSIF x =- 1880 THEN
            sigmoid_f := 584;
        ELSIF x =- 1879 THEN
            sigmoid_f := 584;
        ELSIF x =- 1878 THEN
            sigmoid_f := 585;
        ELSIF x =- 1877 THEN
            sigmoid_f := 585;
        ELSIF x =- 1876 THEN
            sigmoid_f := 585;
        ELSIF x =- 1875 THEN
            sigmoid_f := 585;
        ELSIF x =- 1874 THEN
            sigmoid_f := 586;
        ELSIF x =- 1873 THEN
            sigmoid_f := 586;
        ELSIF x =- 1872 THEN
            sigmoid_f := 586;
        ELSIF x =- 1871 THEN
            sigmoid_f := 586;
        ELSIF x =- 1870 THEN
            sigmoid_f := 586;
        ELSIF x =- 1869 THEN
            sigmoid_f := 587;
        ELSIF x =- 1868 THEN
            sigmoid_f := 587;
        ELSIF x =- 1867 THEN
            sigmoid_f := 587;
        ELSIF x =- 1866 THEN
            sigmoid_f := 587;
        ELSIF x =- 1865 THEN
            sigmoid_f := 587;
        ELSIF x =- 1864 THEN
            sigmoid_f := 588;
        ELSIF x =- 1863 THEN
            sigmoid_f := 588;
        ELSIF x =- 1862 THEN
            sigmoid_f := 588;
        ELSIF x =- 1861 THEN
            sigmoid_f := 588;
        ELSIF x =- 1860 THEN
            sigmoid_f := 588;
        ELSIF x =- 1859 THEN
            sigmoid_f := 589;
        ELSIF x =- 1858 THEN
            sigmoid_f := 589;
        ELSIF x =- 1857 THEN
            sigmoid_f := 589;
        ELSIF x =- 1856 THEN
            sigmoid_f := 589;
        ELSIF x =- 1855 THEN
            sigmoid_f := 589;
        ELSIF x =- 1854 THEN
            sigmoid_f := 590;
        ELSIF x =- 1853 THEN
            sigmoid_f := 590;
        ELSIF x =- 1852 THEN
            sigmoid_f := 590;
        ELSIF x =- 1851 THEN
            sigmoid_f := 590;
        ELSIF x =- 1850 THEN
            sigmoid_f := 590;
        ELSIF x =- 1849 THEN
            sigmoid_f := 591;
        ELSIF x =- 1848 THEN
            sigmoid_f := 591;
        ELSIF x =- 1847 THEN
            sigmoid_f := 591;
        ELSIF x =- 1846 THEN
            sigmoid_f := 591;
        ELSIF x =- 1845 THEN
            sigmoid_f := 592;
        ELSIF x =- 1844 THEN
            sigmoid_f := 592;
        ELSIF x =- 1843 THEN
            sigmoid_f := 592;
        ELSIF x =- 1842 THEN
            sigmoid_f := 592;
        ELSIF x =- 1841 THEN
            sigmoid_f := 592;
        ELSIF x =- 1840 THEN
            sigmoid_f := 593;
        ELSIF x =- 1839 THEN
            sigmoid_f := 593;
        ELSIF x =- 1838 THEN
            sigmoid_f := 593;
        ELSIF x =- 1837 THEN
            sigmoid_f := 593;
        ELSIF x =- 1836 THEN
            sigmoid_f := 593;
        ELSIF x =- 1835 THEN
            sigmoid_f := 594;
        ELSIF x =- 1834 THEN
            sigmoid_f := 594;
        ELSIF x =- 1833 THEN
            sigmoid_f := 594;
        ELSIF x =- 1832 THEN
            sigmoid_f := 594;
        ELSIF x =- 1831 THEN
            sigmoid_f := 594;
        ELSIF x =- 1830 THEN
            sigmoid_f := 595;
        ELSIF x =- 1829 THEN
            sigmoid_f := 595;
        ELSIF x =- 1828 THEN
            sigmoid_f := 595;
        ELSIF x =- 1827 THEN
            sigmoid_f := 595;
        ELSIF x =- 1826 THEN
            sigmoid_f := 595;
        ELSIF x =- 1825 THEN
            sigmoid_f := 596;
        ELSIF x =- 1824 THEN
            sigmoid_f := 596;
        ELSIF x =- 1823 THEN
            sigmoid_f := 596;
        ELSIF x =- 1822 THEN
            sigmoid_f := 596;
        ELSIF x =- 1821 THEN
            sigmoid_f := 596;
        ELSIF x =- 1820 THEN
            sigmoid_f := 597;
        ELSIF x =- 1819 THEN
            sigmoid_f := 597;
        ELSIF x =- 1818 THEN
            sigmoid_f := 597;
        ELSIF x =- 1817 THEN
            sigmoid_f := 597;
        ELSIF x =- 1816 THEN
            sigmoid_f := 598;
        ELSIF x =- 1815 THEN
            sigmoid_f := 598;
        ELSIF x =- 1814 THEN
            sigmoid_f := 598;
        ELSIF x =- 1813 THEN
            sigmoid_f := 598;
        ELSIF x =- 1812 THEN
            sigmoid_f := 598;
        ELSIF x =- 1811 THEN
            sigmoid_f := 599;
        ELSIF x =- 1810 THEN
            sigmoid_f := 599;
        ELSIF x =- 1809 THEN
            sigmoid_f := 599;
        ELSIF x =- 1808 THEN
            sigmoid_f := 599;
        ELSIF x =- 1807 THEN
            sigmoid_f := 599;
        ELSIF x =- 1806 THEN
            sigmoid_f := 600;
        ELSIF x =- 1805 THEN
            sigmoid_f := 600;
        ELSIF x =- 1804 THEN
            sigmoid_f := 600;
        ELSIF x =- 1803 THEN
            sigmoid_f := 600;
        ELSIF x =- 1802 THEN
            sigmoid_f := 600;
        ELSIF x =- 1801 THEN
            sigmoid_f := 601;
        ELSIF x =- 1800 THEN
            sigmoid_f := 601;
        ELSIF x =- 1799 THEN
            sigmoid_f := 601;
        ELSIF x =- 1798 THEN
            sigmoid_f := 601;
        ELSIF x =- 1797 THEN
            sigmoid_f := 601;
        ELSIF x =- 1796 THEN
            sigmoid_f := 602;
        ELSIF x =- 1795 THEN
            sigmoid_f := 602;
        ELSIF x =- 1794 THEN
            sigmoid_f := 602;
        ELSIF x =- 1793 THEN
            sigmoid_f := 602;
        ELSIF x =- 1792 THEN
            sigmoid_f := 603;
        ELSIF x =- 1791 THEN
            sigmoid_f := 603;
        ELSIF x =- 1790 THEN
            sigmoid_f := 603;
        ELSIF x =- 1789 THEN
            sigmoid_f := 603;
        ELSIF x =- 1788 THEN
            sigmoid_f := 603;
        ELSIF x =- 1787 THEN
            sigmoid_f := 604;
        ELSIF x =- 1786 THEN
            sigmoid_f := 604;
        ELSIF x =- 1785 THEN
            sigmoid_f := 604;
        ELSIF x =- 1784 THEN
            sigmoid_f := 604;
        ELSIF x =- 1783 THEN
            sigmoid_f := 604;
        ELSIF x =- 1782 THEN
            sigmoid_f := 605;
        ELSIF x =- 1781 THEN
            sigmoid_f := 605;
        ELSIF x =- 1780 THEN
            sigmoid_f := 605;
        ELSIF x =- 1779 THEN
            sigmoid_f := 605;
        ELSIF x =- 1778 THEN
            sigmoid_f := 605;
        ELSIF x =- 1777 THEN
            sigmoid_f := 606;
        ELSIF x =- 1776 THEN
            sigmoid_f := 606;
        ELSIF x =- 1775 THEN
            sigmoid_f := 606;
        ELSIF x =- 1774 THEN
            sigmoid_f := 606;
        ELSIF x =- 1773 THEN
            sigmoid_f := 606;
        ELSIF x =- 1772 THEN
            sigmoid_f := 607;
        ELSIF x =- 1771 THEN
            sigmoid_f := 607;
        ELSIF x =- 1770 THEN
            sigmoid_f := 607;
        ELSIF x =- 1769 THEN
            sigmoid_f := 607;
        ELSIF x =- 1768 THEN
            sigmoid_f := 607;
        ELSIF x =- 1767 THEN
            sigmoid_f := 608;
        ELSIF x =- 1766 THEN
            sigmoid_f := 608;
        ELSIF x =- 1765 THEN
            sigmoid_f := 608;
        ELSIF x =- 1764 THEN
            sigmoid_f := 608;
        ELSIF x =- 1763 THEN
            sigmoid_f := 609;
        ELSIF x =- 1762 THEN
            sigmoid_f := 609;
        ELSIF x =- 1761 THEN
            sigmoid_f := 609;
        ELSIF x =- 1760 THEN
            sigmoid_f := 609;
        ELSIF x =- 1759 THEN
            sigmoid_f := 609;
        ELSIF x =- 1758 THEN
            sigmoid_f := 610;
        ELSIF x =- 1757 THEN
            sigmoid_f := 610;
        ELSIF x =- 1756 THEN
            sigmoid_f := 610;
        ELSIF x =- 1755 THEN
            sigmoid_f := 610;
        ELSIF x =- 1754 THEN
            sigmoid_f := 610;
        ELSIF x =- 1753 THEN
            sigmoid_f := 611;
        ELSIF x =- 1752 THEN
            sigmoid_f := 611;
        ELSIF x =- 1751 THEN
            sigmoid_f := 611;
        ELSIF x =- 1750 THEN
            sigmoid_f := 611;
        ELSIF x =- 1749 THEN
            sigmoid_f := 611;
        ELSIF x =- 1748 THEN
            sigmoid_f := 612;
        ELSIF x =- 1747 THEN
            sigmoid_f := 612;
        ELSIF x =- 1746 THEN
            sigmoid_f := 612;
        ELSIF x =- 1745 THEN
            sigmoid_f := 612;
        ELSIF x =- 1744 THEN
            sigmoid_f := 612;
        ELSIF x =- 1743 THEN
            sigmoid_f := 613;
        ELSIF x =- 1742 THEN
            sigmoid_f := 613;
        ELSIF x =- 1741 THEN
            sigmoid_f := 613;
        ELSIF x =- 1740 THEN
            sigmoid_f := 613;
        ELSIF x =- 1739 THEN
            sigmoid_f := 613;
        ELSIF x =- 1738 THEN
            sigmoid_f := 614;
        ELSIF x =- 1737 THEN
            sigmoid_f := 614;
        ELSIF x =- 1736 THEN
            sigmoid_f := 614;
        ELSIF x =- 1735 THEN
            sigmoid_f := 614;
        ELSIF x =- 1734 THEN
            sigmoid_f := 615;
        ELSIF x =- 1733 THEN
            sigmoid_f := 615;
        ELSIF x =- 1732 THEN
            sigmoid_f := 615;
        ELSIF x =- 1731 THEN
            sigmoid_f := 615;
        ELSIF x =- 1730 THEN
            sigmoid_f := 615;
        ELSIF x =- 1729 THEN
            sigmoid_f := 616;
        ELSIF x =- 1728 THEN
            sigmoid_f := 616;
        ELSIF x =- 1727 THEN
            sigmoid_f := 616;
        ELSIF x =- 1726 THEN
            sigmoid_f := 616;
        ELSIF x =- 1725 THEN
            sigmoid_f := 616;
        ELSIF x =- 1724 THEN
            sigmoid_f := 617;
        ELSIF x =- 1723 THEN
            sigmoid_f := 617;
        ELSIF x =- 1722 THEN
            sigmoid_f := 617;
        ELSIF x =- 1721 THEN
            sigmoid_f := 617;
        ELSIF x =- 1720 THEN
            sigmoid_f := 617;
        ELSIF x =- 1719 THEN
            sigmoid_f := 618;
        ELSIF x =- 1718 THEN
            sigmoid_f := 618;
        ELSIF x =- 1717 THEN
            sigmoid_f := 618;
        ELSIF x =- 1716 THEN
            sigmoid_f := 618;
        ELSIF x =- 1715 THEN
            sigmoid_f := 618;
        ELSIF x =- 1714 THEN
            sigmoid_f := 619;
        ELSIF x =- 1713 THEN
            sigmoid_f := 619;
        ELSIF x =- 1712 THEN
            sigmoid_f := 619;
        ELSIF x =- 1711 THEN
            sigmoid_f := 619;
        ELSIF x =- 1710 THEN
            sigmoid_f := 619;
        ELSIF x =- 1709 THEN
            sigmoid_f := 620;
        ELSIF x =- 1708 THEN
            sigmoid_f := 620;
        ELSIF x =- 1707 THEN
            sigmoid_f := 620;
        ELSIF x =- 1706 THEN
            sigmoid_f := 620;
        ELSIF x =- 1705 THEN
            sigmoid_f := 621;
        ELSIF x =- 1704 THEN
            sigmoid_f := 621;
        ELSIF x =- 1703 THEN
            sigmoid_f := 621;
        ELSIF x =- 1702 THEN
            sigmoid_f := 621;
        ELSIF x =- 1701 THEN
            sigmoid_f := 621;
        ELSIF x =- 1700 THEN
            sigmoid_f := 622;
        ELSIF x =- 1699 THEN
            sigmoid_f := 622;
        ELSIF x =- 1698 THEN
            sigmoid_f := 622;
        ELSIF x =- 1697 THEN
            sigmoid_f := 622;
        ELSIF x =- 1696 THEN
            sigmoid_f := 622;
        ELSIF x =- 1695 THEN
            sigmoid_f := 623;
        ELSIF x =- 1694 THEN
            sigmoid_f := 623;
        ELSIF x =- 1693 THEN
            sigmoid_f := 623;
        ELSIF x =- 1692 THEN
            sigmoid_f := 623;
        ELSIF x =- 1691 THEN
            sigmoid_f := 623;
        ELSIF x =- 1690 THEN
            sigmoid_f := 624;
        ELSIF x =- 1689 THEN
            sigmoid_f := 624;
        ELSIF x =- 1688 THEN
            sigmoid_f := 624;
        ELSIF x =- 1687 THEN
            sigmoid_f := 624;
        ELSIF x =- 1686 THEN
            sigmoid_f := 624;
        ELSIF x =- 1685 THEN
            sigmoid_f := 625;
        ELSIF x =- 1684 THEN
            sigmoid_f := 625;
        ELSIF x =- 1683 THEN
            sigmoid_f := 625;
        ELSIF x =- 1682 THEN
            sigmoid_f := 625;
        ELSIF x =- 1681 THEN
            sigmoid_f := 625;
        ELSIF x =- 1680 THEN
            sigmoid_f := 626;
        ELSIF x =- 1679 THEN
            sigmoid_f := 626;
        ELSIF x =- 1678 THEN
            sigmoid_f := 626;
        ELSIF x =- 1677 THEN
            sigmoid_f := 626;
        ELSIF x =- 1676 THEN
            sigmoid_f := 627;
        ELSIF x =- 1675 THEN
            sigmoid_f := 627;
        ELSIF x =- 1674 THEN
            sigmoid_f := 627;
        ELSIF x =- 1673 THEN
            sigmoid_f := 627;
        ELSIF x =- 1672 THEN
            sigmoid_f := 627;
        ELSIF x =- 1671 THEN
            sigmoid_f := 628;
        ELSIF x =- 1670 THEN
            sigmoid_f := 628;
        ELSIF x =- 1669 THEN
            sigmoid_f := 628;
        ELSIF x =- 1668 THEN
            sigmoid_f := 628;
        ELSIF x =- 1667 THEN
            sigmoid_f := 628;
        ELSIF x =- 1666 THEN
            sigmoid_f := 629;
        ELSIF x =- 1665 THEN
            sigmoid_f := 629;
        ELSIF x =- 1664 THEN
            sigmoid_f := 629;
        ELSIF x =- 1663 THEN
            sigmoid_f := 629;
        ELSIF x =- 1662 THEN
            sigmoid_f := 629;
        ELSIF x =- 1661 THEN
            sigmoid_f := 630;
        ELSIF x =- 1660 THEN
            sigmoid_f := 630;
        ELSIF x =- 1659 THEN
            sigmoid_f := 630;
        ELSIF x =- 1658 THEN
            sigmoid_f := 630;
        ELSIF x =- 1657 THEN
            sigmoid_f := 630;
        ELSIF x =- 1656 THEN
            sigmoid_f := 631;
        ELSIF x =- 1655 THEN
            sigmoid_f := 631;
        ELSIF x =- 1654 THEN
            sigmoid_f := 631;
        ELSIF x =- 1653 THEN
            sigmoid_f := 631;
        ELSIF x =- 1652 THEN
            sigmoid_f := 631;
        ELSIF x =- 1651 THEN
            sigmoid_f := 632;
        ELSIF x =- 1650 THEN
            sigmoid_f := 632;
        ELSIF x =- 1649 THEN
            sigmoid_f := 632;
        ELSIF x =- 1648 THEN
            sigmoid_f := 632;
        ELSIF x =- 1647 THEN
            sigmoid_f := 633;
        ELSIF x =- 1646 THEN
            sigmoid_f := 633;
        ELSIF x =- 1645 THEN
            sigmoid_f := 633;
        ELSIF x =- 1644 THEN
            sigmoid_f := 633;
        ELSIF x =- 1643 THEN
            sigmoid_f := 633;
        ELSIF x =- 1642 THEN
            sigmoid_f := 634;
        ELSIF x =- 1641 THEN
            sigmoid_f := 634;
        ELSIF x =- 1640 THEN
            sigmoid_f := 634;
        ELSIF x =- 1639 THEN
            sigmoid_f := 634;
        ELSIF x =- 1638 THEN
            sigmoid_f := 634;
        ELSIF x =- 1637 THEN
            sigmoid_f := 635;
        ELSIF x =- 1636 THEN
            sigmoid_f := 635;
        ELSIF x =- 1635 THEN
            sigmoid_f := 635;
        ELSIF x =- 1634 THEN
            sigmoid_f := 635;
        ELSIF x =- 1633 THEN
            sigmoid_f := 635;
        ELSIF x =- 1632 THEN
            sigmoid_f := 636;
        ELSIF x =- 1631 THEN
            sigmoid_f := 636;
        ELSIF x =- 1630 THEN
            sigmoid_f := 636;
        ELSIF x =- 1629 THEN
            sigmoid_f := 636;
        ELSIF x =- 1628 THEN
            sigmoid_f := 636;
        ELSIF x =- 1627 THEN
            sigmoid_f := 637;
        ELSIF x =- 1626 THEN
            sigmoid_f := 637;
        ELSIF x =- 1625 THEN
            sigmoid_f := 637;
        ELSIF x =- 1624 THEN
            sigmoid_f := 637;
        ELSIF x =- 1623 THEN
            sigmoid_f := 637;
        ELSIF x =- 1622 THEN
            sigmoid_f := 638;
        ELSIF x =- 1621 THEN
            sigmoid_f := 638;
        ELSIF x =- 1620 THEN
            sigmoid_f := 638;
        ELSIF x =- 1619 THEN
            sigmoid_f := 638;
        ELSIF x =- 1618 THEN
            sigmoid_f := 639;
        ELSIF x =- 1617 THEN
            sigmoid_f := 639;
        ELSIF x =- 1616 THEN
            sigmoid_f := 639;
        ELSIF x =- 1615 THEN
            sigmoid_f := 639;
        ELSIF x =- 1614 THEN
            sigmoid_f := 639;
        ELSIF x =- 1613 THEN
            sigmoid_f := 640;
        ELSIF x =- 1612 THEN
            sigmoid_f := 640;
        ELSIF x =- 1611 THEN
            sigmoid_f := 640;
        ELSIF x =- 1610 THEN
            sigmoid_f := 640;
        ELSIF x =- 1609 THEN
            sigmoid_f := 640;
        ELSIF x =- 1608 THEN
            sigmoid_f := 641;
        ELSIF x =- 1607 THEN
            sigmoid_f := 641;
        ELSIF x =- 1606 THEN
            sigmoid_f := 641;
        ELSIF x =- 1605 THEN
            sigmoid_f := 641;
        ELSIF x =- 1604 THEN
            sigmoid_f := 641;
        ELSIF x =- 1603 THEN
            sigmoid_f := 642;
        ELSIF x =- 1602 THEN
            sigmoid_f := 642;
        ELSIF x =- 1601 THEN
            sigmoid_f := 642;
        ELSIF x =- 1600 THEN
            sigmoid_f := 642;
        ELSIF x =- 1599 THEN
            sigmoid_f := 642;
        ELSIF x =- 1598 THEN
            sigmoid_f := 643;
        ELSIF x =- 1597 THEN
            sigmoid_f := 643;
        ELSIF x =- 1596 THEN
            sigmoid_f := 643;
        ELSIF x =- 1595 THEN
            sigmoid_f := 643;
        ELSIF x =- 1594 THEN
            sigmoid_f := 643;
        ELSIF x =- 1593 THEN
            sigmoid_f := 644;
        ELSIF x =- 1592 THEN
            sigmoid_f := 644;
        ELSIF x =- 1591 THEN
            sigmoid_f := 644;
        ELSIF x =- 1590 THEN
            sigmoid_f := 644;
        ELSIF x =- 1589 THEN
            sigmoid_f := 645;
        ELSIF x =- 1588 THEN
            sigmoid_f := 645;
        ELSIF x =- 1587 THEN
            sigmoid_f := 645;
        ELSIF x =- 1586 THEN
            sigmoid_f := 645;
        ELSIF x =- 1585 THEN
            sigmoid_f := 645;
        ELSIF x =- 1584 THEN
            sigmoid_f := 646;
        ELSIF x =- 1583 THEN
            sigmoid_f := 646;
        ELSIF x =- 1582 THEN
            sigmoid_f := 646;
        ELSIF x =- 1581 THEN
            sigmoid_f := 646;
        ELSIF x =- 1580 THEN
            sigmoid_f := 646;
        ELSIF x =- 1579 THEN
            sigmoid_f := 647;
        ELSIF x =- 1578 THEN
            sigmoid_f := 647;
        ELSIF x =- 1577 THEN
            sigmoid_f := 647;
        ELSIF x =- 1576 THEN
            sigmoid_f := 647;
        ELSIF x =- 1575 THEN
            sigmoid_f := 647;
        ELSIF x =- 1574 THEN
            sigmoid_f := 648;
        ELSIF x =- 1573 THEN
            sigmoid_f := 648;
        ELSIF x =- 1572 THEN
            sigmoid_f := 648;
        ELSIF x =- 1571 THEN
            sigmoid_f := 648;
        ELSIF x =- 1570 THEN
            sigmoid_f := 648;
        ELSIF x =- 1569 THEN
            sigmoid_f := 649;
        ELSIF x =- 1568 THEN
            sigmoid_f := 649;
        ELSIF x =- 1567 THEN
            sigmoid_f := 649;
        ELSIF x =- 1566 THEN
            sigmoid_f := 649;
        ELSIF x =- 1565 THEN
            sigmoid_f := 649;
        ELSIF x =- 1564 THEN
            sigmoid_f := 650;
        ELSIF x =- 1563 THEN
            sigmoid_f := 650;
        ELSIF x =- 1562 THEN
            sigmoid_f := 650;
        ELSIF x =- 1561 THEN
            sigmoid_f := 650;
        ELSIF x =- 1560 THEN
            sigmoid_f := 651;
        ELSIF x =- 1559 THEN
            sigmoid_f := 651;
        ELSIF x =- 1558 THEN
            sigmoid_f := 651;
        ELSIF x =- 1557 THEN
            sigmoid_f := 651;
        ELSIF x =- 1556 THEN
            sigmoid_f := 651;
        ELSIF x =- 1555 THEN
            sigmoid_f := 652;
        ELSIF x =- 1554 THEN
            sigmoid_f := 652;
        ELSIF x =- 1553 THEN
            sigmoid_f := 652;
        ELSIF x =- 1552 THEN
            sigmoid_f := 652;
        ELSIF x =- 1551 THEN
            sigmoid_f := 652;
        ELSIF x =- 1550 THEN
            sigmoid_f := 653;
        ELSIF x =- 1549 THEN
            sigmoid_f := 653;
        ELSIF x =- 1548 THEN
            sigmoid_f := 653;
        ELSIF x =- 1547 THEN
            sigmoid_f := 653;
        ELSIF x =- 1546 THEN
            sigmoid_f := 653;
        ELSIF x =- 1545 THEN
            sigmoid_f := 654;
        ELSIF x =- 1544 THEN
            sigmoid_f := 654;
        ELSIF x =- 1543 THEN
            sigmoid_f := 654;
        ELSIF x =- 1542 THEN
            sigmoid_f := 654;
        ELSIF x =- 1541 THEN
            sigmoid_f := 654;
        ELSIF x =- 1540 THEN
            sigmoid_f := 655;
        ELSIF x =- 1539 THEN
            sigmoid_f := 655;
        ELSIF x =- 1538 THEN
            sigmoid_f := 655;
        ELSIF x =- 1537 THEN
            sigmoid_f := 655;
        ELSIF x =- 1536 THEN
            sigmoid_f := 656;
        ELSIF x =- 1535 THEN
            sigmoid_f := 656;
        ELSIF x =- 1534 THEN
            sigmoid_f := 656;
        ELSIF x =- 1533 THEN
            sigmoid_f := 656;
        ELSIF x =- 1532 THEN
            sigmoid_f := 657;
        ELSIF x =- 1531 THEN
            sigmoid_f := 657;
        ELSIF x =- 1530 THEN
            sigmoid_f := 657;
        ELSIF x =- 1529 THEN
            sigmoid_f := 657;
        ELSIF x =- 1528 THEN
            sigmoid_f := 658;
        ELSIF x =- 1527 THEN
            sigmoid_f := 658;
        ELSIF x =- 1526 THEN
            sigmoid_f := 658;
        ELSIF x =- 1525 THEN
            sigmoid_f := 658;
        ELSIF x =- 1524 THEN
            sigmoid_f := 658;
        ELSIF x =- 1523 THEN
            sigmoid_f := 659;
        ELSIF x =- 1522 THEN
            sigmoid_f := 659;
        ELSIF x =- 1521 THEN
            sigmoid_f := 659;
        ELSIF x =- 1520 THEN
            sigmoid_f := 659;
        ELSIF x =- 1519 THEN
            sigmoid_f := 660;
        ELSIF x =- 1518 THEN
            sigmoid_f := 660;
        ELSIF x =- 1517 THEN
            sigmoid_f := 660;
        ELSIF x =- 1516 THEN
            sigmoid_f := 660;
        ELSIF x =- 1515 THEN
            sigmoid_f := 661;
        ELSIF x =- 1514 THEN
            sigmoid_f := 661;
        ELSIF x =- 1513 THEN
            sigmoid_f := 661;
        ELSIF x =- 1512 THEN
            sigmoid_f := 661;
        ELSIF x =- 1511 THEN
            sigmoid_f := 661;
        ELSIF x =- 1510 THEN
            sigmoid_f := 662;
        ELSIF x =- 1509 THEN
            sigmoid_f := 662;
        ELSIF x =- 1508 THEN
            sigmoid_f := 662;
        ELSIF x =- 1507 THEN
            sigmoid_f := 662;
        ELSIF x =- 1506 THEN
            sigmoid_f := 663;
        ELSIF x =- 1505 THEN
            sigmoid_f := 663;
        ELSIF x =- 1504 THEN
            sigmoid_f := 663;
        ELSIF x =- 1503 THEN
            sigmoid_f := 663;
        ELSIF x =- 1502 THEN
            sigmoid_f := 663;
        ELSIF x =- 1501 THEN
            sigmoid_f := 664;
        ELSIF x =- 1500 THEN
            sigmoid_f := 664;
        ELSIF x =- 1499 THEN
            sigmoid_f := 664;
        ELSIF x =- 1498 THEN
            sigmoid_f := 664;
        ELSIF x =- 1497 THEN
            sigmoid_f := 665;
        ELSIF x =- 1496 THEN
            sigmoid_f := 665;
        ELSIF x =- 1495 THEN
            sigmoid_f := 665;
        ELSIF x =- 1494 THEN
            sigmoid_f := 665;
        ELSIF x =- 1493 THEN
            sigmoid_f := 666;
        ELSIF x =- 1492 THEN
            sigmoid_f := 666;
        ELSIF x =- 1491 THEN
            sigmoid_f := 666;
        ELSIF x =- 1490 THEN
            sigmoid_f := 666;
        ELSIF x =- 1489 THEN
            sigmoid_f := 666;
        ELSIF x =- 1488 THEN
            sigmoid_f := 667;
        ELSIF x =- 1487 THEN
            sigmoid_f := 667;
        ELSIF x =- 1486 THEN
            sigmoid_f := 667;
        ELSIF x =- 1485 THEN
            sigmoid_f := 667;
        ELSIF x =- 1484 THEN
            sigmoid_f := 668;
        ELSIF x =- 1483 THEN
            sigmoid_f := 668;
        ELSIF x =- 1482 THEN
            sigmoid_f := 668;
        ELSIF x =- 1481 THEN
            sigmoid_f := 668;
        ELSIF x =- 1480 THEN
            sigmoid_f := 668;
        ELSIF x =- 1479 THEN
            sigmoid_f := 669;
        ELSIF x =- 1478 THEN
            sigmoid_f := 669;
        ELSIF x =- 1477 THEN
            sigmoid_f := 669;
        ELSIF x =- 1476 THEN
            sigmoid_f := 669;
        ELSIF x =- 1475 THEN
            sigmoid_f := 670;
        ELSIF x =- 1474 THEN
            sigmoid_f := 670;
        ELSIF x =- 1473 THEN
            sigmoid_f := 670;
        ELSIF x =- 1472 THEN
            sigmoid_f := 670;
        ELSIF x =- 1471 THEN
            sigmoid_f := 671;
        ELSIF x =- 1470 THEN
            sigmoid_f := 671;
        ELSIF x =- 1469 THEN
            sigmoid_f := 671;
        ELSIF x =- 1468 THEN
            sigmoid_f := 671;
        ELSIF x =- 1467 THEN
            sigmoid_f := 671;
        ELSIF x =- 1466 THEN
            sigmoid_f := 672;
        ELSIF x =- 1465 THEN
            sigmoid_f := 672;
        ELSIF x =- 1464 THEN
            sigmoid_f := 672;
        ELSIF x =- 1463 THEN
            sigmoid_f := 672;
        ELSIF x =- 1462 THEN
            sigmoid_f := 673;
        ELSIF x =- 1461 THEN
            sigmoid_f := 673;
        ELSIF x =- 1460 THEN
            sigmoid_f := 673;
        ELSIF x =- 1459 THEN
            sigmoid_f := 673;
        ELSIF x =- 1458 THEN
            sigmoid_f := 673;
        ELSIF x =- 1457 THEN
            sigmoid_f := 674;
        ELSIF x =- 1456 THEN
            sigmoid_f := 674;
        ELSIF x =- 1455 THEN
            sigmoid_f := 674;
        ELSIF x =- 1454 THEN
            sigmoid_f := 674;
        ELSIF x =- 1453 THEN
            sigmoid_f := 675;
        ELSIF x =- 1452 THEN
            sigmoid_f := 675;
        ELSIF x =- 1451 THEN
            sigmoid_f := 675;
        ELSIF x =- 1450 THEN
            sigmoid_f := 675;
        ELSIF x =- 1449 THEN
            sigmoid_f := 676;
        ELSIF x =- 1448 THEN
            sigmoid_f := 676;
        ELSIF x =- 1447 THEN
            sigmoid_f := 676;
        ELSIF x =- 1446 THEN
            sigmoid_f := 676;
        ELSIF x =- 1445 THEN
            sigmoid_f := 676;
        ELSIF x =- 1444 THEN
            sigmoid_f := 677;
        ELSIF x =- 1443 THEN
            sigmoid_f := 677;
        ELSIF x =- 1442 THEN
            sigmoid_f := 677;
        ELSIF x =- 1441 THEN
            sigmoid_f := 677;
        ELSIF x =- 1440 THEN
            sigmoid_f := 678;
        ELSIF x =- 1439 THEN
            sigmoid_f := 678;
        ELSIF x =- 1438 THEN
            sigmoid_f := 678;
        ELSIF x =- 1437 THEN
            sigmoid_f := 678;
        ELSIF x =- 1436 THEN
            sigmoid_f := 678;
        ELSIF x =- 1435 THEN
            sigmoid_f := 679;
        ELSIF x =- 1434 THEN
            sigmoid_f := 679;
        ELSIF x =- 1433 THEN
            sigmoid_f := 679;
        ELSIF x =- 1432 THEN
            sigmoid_f := 679;
        ELSIF x =- 1431 THEN
            sigmoid_f := 680;
        ELSIF x =- 1430 THEN
            sigmoid_f := 680;
        ELSIF x =- 1429 THEN
            sigmoid_f := 680;
        ELSIF x =- 1428 THEN
            sigmoid_f := 680;
        ELSIF x =- 1427 THEN
            sigmoid_f := 680;
        ELSIF x =- 1426 THEN
            sigmoid_f := 681;
        ELSIF x =- 1425 THEN
            sigmoid_f := 681;
        ELSIF x =- 1424 THEN
            sigmoid_f := 681;
        ELSIF x =- 1423 THEN
            sigmoid_f := 681;
        ELSIF x =- 1422 THEN
            sigmoid_f := 682;
        ELSIF x =- 1421 THEN
            sigmoid_f := 682;
        ELSIF x =- 1420 THEN
            sigmoid_f := 682;
        ELSIF x =- 1419 THEN
            sigmoid_f := 682;
        ELSIF x =- 1418 THEN
            sigmoid_f := 683;
        ELSIF x =- 1417 THEN
            sigmoid_f := 683;
        ELSIF x =- 1416 THEN
            sigmoid_f := 683;
        ELSIF x =- 1415 THEN
            sigmoid_f := 683;
        ELSIF x =- 1414 THEN
            sigmoid_f := 683;
        ELSIF x =- 1413 THEN
            sigmoid_f := 684;
        ELSIF x =- 1412 THEN
            sigmoid_f := 684;
        ELSIF x =- 1411 THEN
            sigmoid_f := 684;
        ELSIF x =- 1410 THEN
            sigmoid_f := 684;
        ELSIF x =- 1409 THEN
            sigmoid_f := 685;
        ELSIF x =- 1408 THEN
            sigmoid_f := 685;
        ELSIF x =- 1407 THEN
            sigmoid_f := 685;
        ELSIF x =- 1406 THEN
            sigmoid_f := 685;
        ELSIF x =- 1405 THEN
            sigmoid_f := 685;
        ELSIF x =- 1404 THEN
            sigmoid_f := 686;
        ELSIF x =- 1403 THEN
            sigmoid_f := 686;
        ELSIF x =- 1402 THEN
            sigmoid_f := 686;
        ELSIF x =- 1401 THEN
            sigmoid_f := 686;
        ELSIF x =- 1400 THEN
            sigmoid_f := 687;
        ELSIF x =- 1399 THEN
            sigmoid_f := 687;
        ELSIF x =- 1398 THEN
            sigmoid_f := 687;
        ELSIF x =- 1397 THEN
            sigmoid_f := 687;
        ELSIF x =- 1396 THEN
            sigmoid_f := 688;
        ELSIF x =- 1395 THEN
            sigmoid_f := 688;
        ELSIF x =- 1394 THEN
            sigmoid_f := 688;
        ELSIF x =- 1393 THEN
            sigmoid_f := 688;
        ELSIF x =- 1392 THEN
            sigmoid_f := 688;
        ELSIF x =- 1391 THEN
            sigmoid_f := 689;
        ELSIF x =- 1390 THEN
            sigmoid_f := 689;
        ELSIF x =- 1389 THEN
            sigmoid_f := 689;
        ELSIF x =- 1388 THEN
            sigmoid_f := 689;
        ELSIF x =- 1387 THEN
            sigmoid_f := 690;
        ELSIF x =- 1386 THEN
            sigmoid_f := 690;
        ELSIF x =- 1385 THEN
            sigmoid_f := 690;
        ELSIF x =- 1384 THEN
            sigmoid_f := 690;
        ELSIF x =- 1383 THEN
            sigmoid_f := 690;
        ELSIF x =- 1382 THEN
            sigmoid_f := 691;
        ELSIF x =- 1381 THEN
            sigmoid_f := 691;
        ELSIF x =- 1380 THEN
            sigmoid_f := 691;
        ELSIF x =- 1379 THEN
            sigmoid_f := 691;
        ELSIF x =- 1378 THEN
            sigmoid_f := 692;
        ELSIF x =- 1377 THEN
            sigmoid_f := 692;
        ELSIF x =- 1376 THEN
            sigmoid_f := 692;
        ELSIF x =- 1375 THEN
            sigmoid_f := 692;
        ELSIF x =- 1374 THEN
            sigmoid_f := 693;
        ELSIF x =- 1373 THEN
            sigmoid_f := 693;
        ELSIF x =- 1372 THEN
            sigmoid_f := 693;
        ELSIF x =- 1371 THEN
            sigmoid_f := 693;
        ELSIF x =- 1370 THEN
            sigmoid_f := 693;
        ELSIF x =- 1369 THEN
            sigmoid_f := 694;
        ELSIF x =- 1368 THEN
            sigmoid_f := 694;
        ELSIF x =- 1367 THEN
            sigmoid_f := 694;
        ELSIF x =- 1366 THEN
            sigmoid_f := 694;
        ELSIF x =- 1365 THEN
            sigmoid_f := 695;
        ELSIF x =- 1364 THEN
            sigmoid_f := 695;
        ELSIF x =- 1363 THEN
            sigmoid_f := 695;
        ELSIF x =- 1362 THEN
            sigmoid_f := 695;
        ELSIF x =- 1361 THEN
            sigmoid_f := 695;
        ELSIF x =- 1360 THEN
            sigmoid_f := 696;
        ELSIF x =- 1359 THEN
            sigmoid_f := 696;
        ELSIF x =- 1358 THEN
            sigmoid_f := 696;
        ELSIF x =- 1357 THEN
            sigmoid_f := 696;
        ELSIF x =- 1356 THEN
            sigmoid_f := 697;
        ELSIF x =- 1355 THEN
            sigmoid_f := 697;
        ELSIF x =- 1354 THEN
            sigmoid_f := 697;
        ELSIF x =- 1353 THEN
            sigmoid_f := 697;
        ELSIF x =- 1352 THEN
            sigmoid_f := 698;
        ELSIF x =- 1351 THEN
            sigmoid_f := 698;
        ELSIF x =- 1350 THEN
            sigmoid_f := 698;
        ELSIF x =- 1349 THEN
            sigmoid_f := 698;
        ELSIF x =- 1348 THEN
            sigmoid_f := 698;
        ELSIF x =- 1347 THEN
            sigmoid_f := 699;
        ELSIF x =- 1346 THEN
            sigmoid_f := 699;
        ELSIF x =- 1345 THEN
            sigmoid_f := 699;
        ELSIF x =- 1344 THEN
            sigmoid_f := 699;
        ELSIF x =- 1343 THEN
            sigmoid_f := 700;
        ELSIF x =- 1342 THEN
            sigmoid_f := 700;
        ELSIF x =- 1341 THEN
            sigmoid_f := 700;
        ELSIF x =- 1340 THEN
            sigmoid_f := 700;
        ELSIF x =- 1339 THEN
            sigmoid_f := 700;
        ELSIF x =- 1338 THEN
            sigmoid_f := 701;
        ELSIF x =- 1337 THEN
            sigmoid_f := 701;
        ELSIF x =- 1336 THEN
            sigmoid_f := 701;
        ELSIF x =- 1335 THEN
            sigmoid_f := 701;
        ELSIF x =- 1334 THEN
            sigmoid_f := 702;
        ELSIF x =- 1333 THEN
            sigmoid_f := 702;
        ELSIF x =- 1332 THEN
            sigmoid_f := 702;
        ELSIF x =- 1331 THEN
            sigmoid_f := 702;
        ELSIF x =- 1330 THEN
            sigmoid_f := 703;
        ELSIF x =- 1329 THEN
            sigmoid_f := 703;
        ELSIF x =- 1328 THEN
            sigmoid_f := 703;
        ELSIF x =- 1327 THEN
            sigmoid_f := 703;
        ELSIF x =- 1326 THEN
            sigmoid_f := 703;
        ELSIF x =- 1325 THEN
            sigmoid_f := 704;
        ELSIF x =- 1324 THEN
            sigmoid_f := 704;
        ELSIF x =- 1323 THEN
            sigmoid_f := 704;
        ELSIF x =- 1322 THEN
            sigmoid_f := 704;
        ELSIF x =- 1321 THEN
            sigmoid_f := 705;
        ELSIF x =- 1320 THEN
            sigmoid_f := 705;
        ELSIF x =- 1319 THEN
            sigmoid_f := 705;
        ELSIF x =- 1318 THEN
            sigmoid_f := 705;
        ELSIF x =- 1317 THEN
            sigmoid_f := 705;
        ELSIF x =- 1316 THEN
            sigmoid_f := 706;
        ELSIF x =- 1315 THEN
            sigmoid_f := 706;
        ELSIF x =- 1314 THEN
            sigmoid_f := 706;
        ELSIF x =- 1313 THEN
            sigmoid_f := 706;
        ELSIF x =- 1312 THEN
            sigmoid_f := 707;
        ELSIF x =- 1311 THEN
            sigmoid_f := 707;
        ELSIF x =- 1310 THEN
            sigmoid_f := 707;
        ELSIF x =- 1309 THEN
            sigmoid_f := 707;
        ELSIF x =- 1308 THEN
            sigmoid_f := 708;
        ELSIF x =- 1307 THEN
            sigmoid_f := 708;
        ELSIF x =- 1306 THEN
            sigmoid_f := 708;
        ELSIF x =- 1305 THEN
            sigmoid_f := 708;
        ELSIF x =- 1304 THEN
            sigmoid_f := 708;
        ELSIF x =- 1303 THEN
            sigmoid_f := 709;
        ELSIF x =- 1302 THEN
            sigmoid_f := 709;
        ELSIF x =- 1301 THEN
            sigmoid_f := 709;
        ELSIF x =- 1300 THEN
            sigmoid_f := 709;
        ELSIF x =- 1299 THEN
            sigmoid_f := 710;
        ELSIF x =- 1298 THEN
            sigmoid_f := 710;
        ELSIF x =- 1297 THEN
            sigmoid_f := 710;
        ELSIF x =- 1296 THEN
            sigmoid_f := 710;
        ELSIF x =- 1295 THEN
            sigmoid_f := 710;
        ELSIF x =- 1294 THEN
            sigmoid_f := 711;
        ELSIF x =- 1293 THEN
            sigmoid_f := 711;
        ELSIF x =- 1292 THEN
            sigmoid_f := 711;
        ELSIF x =- 1291 THEN
            sigmoid_f := 711;
        ELSIF x =- 1290 THEN
            sigmoid_f := 712;
        ELSIF x =- 1289 THEN
            sigmoid_f := 712;
        ELSIF x =- 1288 THEN
            sigmoid_f := 712;
        ELSIF x =- 1287 THEN
            sigmoid_f := 712;
        ELSIF x =- 1286 THEN
            sigmoid_f := 713;
        ELSIF x =- 1285 THEN
            sigmoid_f := 713;
        ELSIF x =- 1284 THEN
            sigmoid_f := 713;
        ELSIF x =- 1283 THEN
            sigmoid_f := 713;
        ELSIF x =- 1282 THEN
            sigmoid_f := 713;
        ELSIF x =- 1281 THEN
            sigmoid_f := 714;
        ELSIF x =- 1280 THEN
            sigmoid_f := 714;
        ELSIF x =- 1279 THEN
            sigmoid_f := 714;
        ELSIF x =- 1278 THEN
            sigmoid_f := 714;
        ELSIF x =- 1277 THEN
            sigmoid_f := 715;
        ELSIF x =- 1276 THEN
            sigmoid_f := 715;
        ELSIF x =- 1275 THEN
            sigmoid_f := 715;
        ELSIF x =- 1274 THEN
            sigmoid_f := 715;
        ELSIF x =- 1273 THEN
            sigmoid_f := 715;
        ELSIF x =- 1272 THEN
            sigmoid_f := 716;
        ELSIF x =- 1271 THEN
            sigmoid_f := 716;
        ELSIF x =- 1270 THEN
            sigmoid_f := 716;
        ELSIF x =- 1269 THEN
            sigmoid_f := 716;
        ELSIF x =- 1268 THEN
            sigmoid_f := 717;
        ELSIF x =- 1267 THEN
            sigmoid_f := 717;
        ELSIF x =- 1266 THEN
            sigmoid_f := 717;
        ELSIF x =- 1265 THEN
            sigmoid_f := 717;
        ELSIF x =- 1264 THEN
            sigmoid_f := 718;
        ELSIF x =- 1263 THEN
            sigmoid_f := 718;
        ELSIF x =- 1262 THEN
            sigmoid_f := 718;
        ELSIF x =- 1261 THEN
            sigmoid_f := 718;
        ELSIF x =- 1260 THEN
            sigmoid_f := 718;
        ELSIF x =- 1259 THEN
            sigmoid_f := 719;
        ELSIF x =- 1258 THEN
            sigmoid_f := 719;
        ELSIF x =- 1257 THEN
            sigmoid_f := 719;
        ELSIF x =- 1256 THEN
            sigmoid_f := 719;
        ELSIF x =- 1255 THEN
            sigmoid_f := 720;
        ELSIF x =- 1254 THEN
            sigmoid_f := 720;
        ELSIF x =- 1253 THEN
            sigmoid_f := 720;
        ELSIF x =- 1252 THEN
            sigmoid_f := 720;
        ELSIF x =- 1251 THEN
            sigmoid_f := 720;
        ELSIF x =- 1250 THEN
            sigmoid_f := 721;
        ELSIF x =- 1249 THEN
            sigmoid_f := 721;
        ELSIF x =- 1248 THEN
            sigmoid_f := 721;
        ELSIF x =- 1247 THEN
            sigmoid_f := 721;
        ELSIF x =- 1246 THEN
            sigmoid_f := 722;
        ELSIF x =- 1245 THEN
            sigmoid_f := 722;
        ELSIF x =- 1244 THEN
            sigmoid_f := 722;
        ELSIF x =- 1243 THEN
            sigmoid_f := 722;
        ELSIF x =- 1242 THEN
            sigmoid_f := 723;
        ELSIF x =- 1241 THEN
            sigmoid_f := 723;
        ELSIF x =- 1240 THEN
            sigmoid_f := 723;
        ELSIF x =- 1239 THEN
            sigmoid_f := 723;
        ELSIF x =- 1238 THEN
            sigmoid_f := 723;
        ELSIF x =- 1237 THEN
            sigmoid_f := 724;
        ELSIF x =- 1236 THEN
            sigmoid_f := 724;
        ELSIF x =- 1235 THEN
            sigmoid_f := 724;
        ELSIF x =- 1234 THEN
            sigmoid_f := 724;
        ELSIF x =- 1233 THEN
            sigmoid_f := 725;
        ELSIF x =- 1232 THEN
            sigmoid_f := 725;
        ELSIF x =- 1231 THEN
            sigmoid_f := 725;
        ELSIF x =- 1230 THEN
            sigmoid_f := 725;
        ELSIF x =- 1229 THEN
            sigmoid_f := 725;
        ELSIF x =- 1228 THEN
            sigmoid_f := 726;
        ELSIF x =- 1227 THEN
            sigmoid_f := 726;
        ELSIF x =- 1226 THEN
            sigmoid_f := 726;
        ELSIF x =- 1225 THEN
            sigmoid_f := 726;
        ELSIF x =- 1224 THEN
            sigmoid_f := 727;
        ELSIF x =- 1223 THEN
            sigmoid_f := 727;
        ELSIF x =- 1222 THEN
            sigmoid_f := 727;
        ELSIF x =- 1221 THEN
            sigmoid_f := 727;
        ELSIF x =- 1220 THEN
            sigmoid_f := 727;
        ELSIF x =- 1219 THEN
            sigmoid_f := 728;
        ELSIF x =- 1218 THEN
            sigmoid_f := 728;
        ELSIF x =- 1217 THEN
            sigmoid_f := 728;
        ELSIF x =- 1216 THEN
            sigmoid_f := 728;
        ELSIF x =- 1215 THEN
            sigmoid_f := 729;
        ELSIF x =- 1214 THEN
            sigmoid_f := 729;
        ELSIF x =- 1213 THEN
            sigmoid_f := 729;
        ELSIF x =- 1212 THEN
            sigmoid_f := 729;
        ELSIF x =- 1211 THEN
            sigmoid_f := 730;
        ELSIF x =- 1210 THEN
            sigmoid_f := 730;
        ELSIF x =- 1209 THEN
            sigmoid_f := 730;
        ELSIF x =- 1208 THEN
            sigmoid_f := 730;
        ELSIF x =- 1207 THEN
            sigmoid_f := 730;
        ELSIF x =- 1206 THEN
            sigmoid_f := 731;
        ELSIF x =- 1205 THEN
            sigmoid_f := 731;
        ELSIF x =- 1204 THEN
            sigmoid_f := 731;
        ELSIF x =- 1203 THEN
            sigmoid_f := 731;
        ELSIF x =- 1202 THEN
            sigmoid_f := 732;
        ELSIF x =- 1201 THEN
            sigmoid_f := 732;
        ELSIF x =- 1200 THEN
            sigmoid_f := 732;
        ELSIF x =- 1199 THEN
            sigmoid_f := 732;
        ELSIF x =- 1198 THEN
            sigmoid_f := 732;
        ELSIF x =- 1197 THEN
            sigmoid_f := 733;
        ELSIF x =- 1196 THEN
            sigmoid_f := 733;
        ELSIF x =- 1195 THEN
            sigmoid_f := 733;
        ELSIF x =- 1194 THEN
            sigmoid_f := 733;
        ELSIF x =- 1193 THEN
            sigmoid_f := 734;
        ELSIF x =- 1192 THEN
            sigmoid_f := 734;
        ELSIF x =- 1191 THEN
            sigmoid_f := 734;
        ELSIF x =- 1190 THEN
            sigmoid_f := 734;
        ELSIF x =- 1189 THEN
            sigmoid_f := 735;
        ELSIF x =- 1188 THEN
            sigmoid_f := 735;
        ELSIF x =- 1187 THEN
            sigmoid_f := 735;
        ELSIF x =- 1186 THEN
            sigmoid_f := 735;
        ELSIF x =- 1185 THEN
            sigmoid_f := 735;
        ELSIF x =- 1184 THEN
            sigmoid_f := 736;
        ELSIF x =- 1183 THEN
            sigmoid_f := 736;
        ELSIF x =- 1182 THEN
            sigmoid_f := 736;
        ELSIF x =- 1181 THEN
            sigmoid_f := 736;
        ELSIF x =- 1180 THEN
            sigmoid_f := 737;
        ELSIF x =- 1179 THEN
            sigmoid_f := 737;
        ELSIF x =- 1178 THEN
            sigmoid_f := 737;
        ELSIF x =- 1177 THEN
            sigmoid_f := 737;
        ELSIF x =- 1176 THEN
            sigmoid_f := 737;
        ELSIF x =- 1175 THEN
            sigmoid_f := 738;
        ELSIF x =- 1174 THEN
            sigmoid_f := 738;
        ELSIF x =- 1173 THEN
            sigmoid_f := 738;
        ELSIF x =- 1172 THEN
            sigmoid_f := 738;
        ELSIF x =- 1171 THEN
            sigmoid_f := 739;
        ELSIF x =- 1170 THEN
            sigmoid_f := 739;
        ELSIF x =- 1169 THEN
            sigmoid_f := 739;
        ELSIF x =- 1168 THEN
            sigmoid_f := 739;
        ELSIF x =- 1167 THEN
            sigmoid_f := 740;
        ELSIF x =- 1166 THEN
            sigmoid_f := 740;
        ELSIF x =- 1165 THEN
            sigmoid_f := 740;
        ELSIF x =- 1164 THEN
            sigmoid_f := 740;
        ELSIF x =- 1163 THEN
            sigmoid_f := 740;
        ELSIF x =- 1162 THEN
            sigmoid_f := 741;
        ELSIF x =- 1161 THEN
            sigmoid_f := 741;
        ELSIF x =- 1160 THEN
            sigmoid_f := 741;
        ELSIF x =- 1159 THEN
            sigmoid_f := 741;
        ELSIF x =- 1158 THEN
            sigmoid_f := 742;
        ELSIF x =- 1157 THEN
            sigmoid_f := 742;
        ELSIF x =- 1156 THEN
            sigmoid_f := 742;
        ELSIF x =- 1155 THEN
            sigmoid_f := 742;
        ELSIF x =- 1154 THEN
            sigmoid_f := 742;
        ELSIF x =- 1153 THEN
            sigmoid_f := 743;
        ELSIF x =- 1152 THEN
            sigmoid_f := 743;
        ELSIF x =- 1151 THEN
            sigmoid_f := 743;
        ELSIF x =- 1150 THEN
            sigmoid_f := 743;
        ELSIF x =- 1149 THEN
            sigmoid_f := 744;
        ELSIF x =- 1148 THEN
            sigmoid_f := 744;
        ELSIF x =- 1147 THEN
            sigmoid_f := 744;
        ELSIF x =- 1146 THEN
            sigmoid_f := 744;
        ELSIF x =- 1145 THEN
            sigmoid_f := 745;
        ELSIF x =- 1144 THEN
            sigmoid_f := 745;
        ELSIF x =- 1143 THEN
            sigmoid_f := 745;
        ELSIF x =- 1142 THEN
            sigmoid_f := 745;
        ELSIF x =- 1141 THEN
            sigmoid_f := 745;
        ELSIF x =- 1140 THEN
            sigmoid_f := 746;
        ELSIF x =- 1139 THEN
            sigmoid_f := 746;
        ELSIF x =- 1138 THEN
            sigmoid_f := 746;
        ELSIF x =- 1137 THEN
            sigmoid_f := 746;
        ELSIF x =- 1136 THEN
            sigmoid_f := 747;
        ELSIF x =- 1135 THEN
            sigmoid_f := 747;
        ELSIF x =- 1134 THEN
            sigmoid_f := 747;
        ELSIF x =- 1133 THEN
            sigmoid_f := 747;
        ELSIF x =- 1132 THEN
            sigmoid_f := 747;
        ELSIF x =- 1131 THEN
            sigmoid_f := 748;
        ELSIF x =- 1130 THEN
            sigmoid_f := 748;
        ELSIF x =- 1129 THEN
            sigmoid_f := 748;
        ELSIF x =- 1128 THEN
            sigmoid_f := 748;
        ELSIF x =- 1127 THEN
            sigmoid_f := 749;
        ELSIF x =- 1126 THEN
            sigmoid_f := 749;
        ELSIF x =- 1125 THEN
            sigmoid_f := 749;
        ELSIF x =- 1124 THEN
            sigmoid_f := 749;
        ELSIF x =- 1123 THEN
            sigmoid_f := 750;
        ELSIF x =- 1122 THEN
            sigmoid_f := 750;
        ELSIF x =- 1121 THEN
            sigmoid_f := 750;
        ELSIF x =- 1120 THEN
            sigmoid_f := 750;
        ELSIF x =- 1119 THEN
            sigmoid_f := 750;
        ELSIF x =- 1118 THEN
            sigmoid_f := 751;
        ELSIF x =- 1117 THEN
            sigmoid_f := 751;
        ELSIF x =- 1116 THEN
            sigmoid_f := 751;
        ELSIF x =- 1115 THEN
            sigmoid_f := 751;
        ELSIF x =- 1114 THEN
            sigmoid_f := 752;
        ELSIF x =- 1113 THEN
            sigmoid_f := 752;
        ELSIF x =- 1112 THEN
            sigmoid_f := 752;
        ELSIF x =- 1111 THEN
            sigmoid_f := 752;
        ELSIF x =- 1110 THEN
            sigmoid_f := 752;
        ELSIF x =- 1109 THEN
            sigmoid_f := 753;
        ELSIF x =- 1108 THEN
            sigmoid_f := 753;
        ELSIF x =- 1107 THEN
            sigmoid_f := 753;
        ELSIF x =- 1106 THEN
            sigmoid_f := 753;
        ELSIF x =- 1105 THEN
            sigmoid_f := 754;
        ELSIF x =- 1104 THEN
            sigmoid_f := 754;
        ELSIF x =- 1103 THEN
            sigmoid_f := 754;
        ELSIF x =- 1102 THEN
            sigmoid_f := 754;
        ELSIF x =- 1101 THEN
            sigmoid_f := 755;
        ELSIF x =- 1100 THEN
            sigmoid_f := 755;
        ELSIF x =- 1099 THEN
            sigmoid_f := 755;
        ELSIF x =- 1098 THEN
            sigmoid_f := 755;
        ELSIF x =- 1097 THEN
            sigmoid_f := 755;
        ELSIF x =- 1096 THEN
            sigmoid_f := 756;
        ELSIF x =- 1095 THEN
            sigmoid_f := 756;
        ELSIF x =- 1094 THEN
            sigmoid_f := 756;
        ELSIF x =- 1093 THEN
            sigmoid_f := 756;
        ELSIF x =- 1092 THEN
            sigmoid_f := 757;
        ELSIF x =- 1091 THEN
            sigmoid_f := 757;
        ELSIF x =- 1090 THEN
            sigmoid_f := 757;
        ELSIF x =- 1089 THEN
            sigmoid_f := 757;
        ELSIF x =- 1088 THEN
            sigmoid_f := 757;
        ELSIF x =- 1087 THEN
            sigmoid_f := 758;
        ELSIF x =- 1086 THEN
            sigmoid_f := 758;
        ELSIF x =- 1085 THEN
            sigmoid_f := 758;
        ELSIF x =- 1084 THEN
            sigmoid_f := 758;
        ELSIF x =- 1083 THEN
            sigmoid_f := 759;
        ELSIF x =- 1082 THEN
            sigmoid_f := 759;
        ELSIF x =- 1081 THEN
            sigmoid_f := 759;
        ELSIF x =- 1080 THEN
            sigmoid_f := 759;
        ELSIF x =- 1079 THEN
            sigmoid_f := 760;
        ELSIF x =- 1078 THEN
            sigmoid_f := 760;
        ELSIF x =- 1077 THEN
            sigmoid_f := 760;
        ELSIF x =- 1076 THEN
            sigmoid_f := 760;
        ELSIF x =- 1075 THEN
            sigmoid_f := 760;
        ELSIF x =- 1074 THEN
            sigmoid_f := 761;
        ELSIF x =- 1073 THEN
            sigmoid_f := 761;
        ELSIF x =- 1072 THEN
            sigmoid_f := 761;
        ELSIF x =- 1071 THEN
            sigmoid_f := 761;
        ELSIF x =- 1070 THEN
            sigmoid_f := 762;
        ELSIF x =- 1069 THEN
            sigmoid_f := 762;
        ELSIF x =- 1068 THEN
            sigmoid_f := 762;
        ELSIF x =- 1067 THEN
            sigmoid_f := 762;
        ELSIF x =- 1066 THEN
            sigmoid_f := 762;
        ELSIF x =- 1065 THEN
            sigmoid_f := 763;
        ELSIF x =- 1064 THEN
            sigmoid_f := 763;
        ELSIF x =- 1063 THEN
            sigmoid_f := 763;
        ELSIF x =- 1062 THEN
            sigmoid_f := 763;
        ELSIF x =- 1061 THEN
            sigmoid_f := 764;
        ELSIF x =- 1060 THEN
            sigmoid_f := 764;
        ELSIF x =- 1059 THEN
            sigmoid_f := 764;
        ELSIF x =- 1058 THEN
            sigmoid_f := 764;
        ELSIF x =- 1057 THEN
            sigmoid_f := 765;
        ELSIF x =- 1056 THEN
            sigmoid_f := 765;
        ELSIF x =- 1055 THEN
            sigmoid_f := 765;
        ELSIF x =- 1054 THEN
            sigmoid_f := 765;
        ELSIF x =- 1053 THEN
            sigmoid_f := 765;
        ELSIF x =- 1052 THEN
            sigmoid_f := 766;
        ELSIF x =- 1051 THEN
            sigmoid_f := 766;
        ELSIF x =- 1050 THEN
            sigmoid_f := 766;
        ELSIF x =- 1049 THEN
            sigmoid_f := 766;
        ELSIF x =- 1048 THEN
            sigmoid_f := 767;
        ELSIF x =- 1047 THEN
            sigmoid_f := 767;
        ELSIF x =- 1046 THEN
            sigmoid_f := 767;
        ELSIF x =- 1045 THEN
            sigmoid_f := 767;
        ELSIF x =- 1044 THEN
            sigmoid_f := 767;
        ELSIF x =- 1043 THEN
            sigmoid_f := 768;
        ELSIF x =- 1042 THEN
            sigmoid_f := 768;
        ELSIF x =- 1041 THEN
            sigmoid_f := 768;
        ELSIF x =- 1040 THEN
            sigmoid_f := 768;
        ELSIF x =- 1039 THEN
            sigmoid_f := 769;
        ELSIF x =- 1038 THEN
            sigmoid_f := 769;
        ELSIF x =- 1037 THEN
            sigmoid_f := 769;
        ELSIF x =- 1036 THEN
            sigmoid_f := 769;
        ELSIF x =- 1035 THEN
            sigmoid_f := 770;
        ELSIF x =- 1034 THEN
            sigmoid_f := 770;
        ELSIF x =- 1033 THEN
            sigmoid_f := 770;
        ELSIF x =- 1032 THEN
            sigmoid_f := 770;
        ELSIF x =- 1031 THEN
            sigmoid_f := 770;
        ELSIF x =- 1030 THEN
            sigmoid_f := 771;
        ELSIF x =- 1029 THEN
            sigmoid_f := 771;
        ELSIF x =- 1028 THEN
            sigmoid_f := 771;
        ELSIF x =- 1027 THEN
            sigmoid_f := 771;
        ELSIF x =- 1026 THEN
            sigmoid_f := 772;
        ELSIF x =- 1025 THEN
            sigmoid_f := 772;
        ELSIF x =- 1024 THEN
            sigmoid_f := 772;
        ELSIF x =- 1023 THEN
            sigmoid_f := 772;
        ELSIF x =- 1022 THEN
            sigmoid_f := 772;
        ELSIF x =- 1021 THEN
            sigmoid_f := 773;
        ELSIF x =- 1020 THEN
            sigmoid_f := 773;
        ELSIF x =- 1019 THEN
            sigmoid_f := 773;
        ELSIF x =- 1018 THEN
            sigmoid_f := 773;
        ELSIF x =- 1017 THEN
            sigmoid_f := 774;
        ELSIF x =- 1016 THEN
            sigmoid_f := 774;
        ELSIF x =- 1015 THEN
            sigmoid_f := 774;
        ELSIF x =- 1014 THEN
            sigmoid_f := 774;
        ELSIF x =- 1013 THEN
            sigmoid_f := 775;
        ELSIF x =- 1012 THEN
            sigmoid_f := 775;
        ELSIF x =- 1011 THEN
            sigmoid_f := 775;
        ELSIF x =- 1010 THEN
            sigmoid_f := 775;
        ELSIF x =- 1009 THEN
            sigmoid_f := 776;
        ELSIF x =- 1008 THEN
            sigmoid_f := 776;
        ELSIF x =- 1007 THEN
            sigmoid_f := 776;
        ELSIF x =- 1006 THEN
            sigmoid_f := 776;
        ELSIF x =- 1005 THEN
            sigmoid_f := 777;
        ELSIF x =- 1004 THEN
            sigmoid_f := 777;
        ELSIF x =- 1003 THEN
            sigmoid_f := 777;
        ELSIF x =- 1002 THEN
            sigmoid_f := 777;
        ELSIF x =- 1001 THEN
            sigmoid_f := 778;
        ELSIF x =- 1000 THEN
            sigmoid_f := 778;
        ELSIF x =- 999 THEN
            sigmoid_f := 778;
        ELSIF x =- 998 THEN
            sigmoid_f := 778;
        ELSIF x =- 997 THEN
            sigmoid_f := 779;
        ELSIF x =- 996 THEN
            sigmoid_f := 779;
        ELSIF x =- 995 THEN
            sigmoid_f := 779;
        ELSIF x =- 994 THEN
            sigmoid_f := 779;
        ELSIF x =- 993 THEN
            sigmoid_f := 779;
        ELSIF x =- 992 THEN
            sigmoid_f := 780;
        ELSIF x =- 991 THEN
            sigmoid_f := 780;
        ELSIF x =- 990 THEN
            sigmoid_f := 780;
        ELSIF x =- 989 THEN
            sigmoid_f := 780;
        ELSIF x =- 988 THEN
            sigmoid_f := 781;
        ELSIF x =- 987 THEN
            sigmoid_f := 781;
        ELSIF x =- 986 THEN
            sigmoid_f := 781;
        ELSIF x =- 985 THEN
            sigmoid_f := 781;
        ELSIF x =- 984 THEN
            sigmoid_f := 782;
        ELSIF x =- 983 THEN
            sigmoid_f := 782;
        ELSIF x =- 982 THEN
            sigmoid_f := 782;
        ELSIF x =- 981 THEN
            sigmoid_f := 782;
        ELSIF x =- 980 THEN
            sigmoid_f := 783;
        ELSIF x =- 979 THEN
            sigmoid_f := 783;
        ELSIF x =- 978 THEN
            sigmoid_f := 783;
        ELSIF x =- 977 THEN
            sigmoid_f := 783;
        ELSIF x =- 976 THEN
            sigmoid_f := 784;
        ELSIF x =- 975 THEN
            sigmoid_f := 784;
        ELSIF x =- 974 THEN
            sigmoid_f := 784;
        ELSIF x =- 973 THEN
            sigmoid_f := 784;
        ELSIF x =- 972 THEN
            sigmoid_f := 785;
        ELSIF x =- 971 THEN
            sigmoid_f := 785;
        ELSIF x =- 970 THEN
            sigmoid_f := 785;
        ELSIF x =- 969 THEN
            sigmoid_f := 785;
        ELSIF x =- 968 THEN
            sigmoid_f := 786;
        ELSIF x =- 967 THEN
            sigmoid_f := 786;
        ELSIF x =- 966 THEN
            sigmoid_f := 786;
        ELSIF x =- 965 THEN
            sigmoid_f := 786;
        ELSIF x =- 964 THEN
            sigmoid_f := 787;
        ELSIF x =- 963 THEN
            sigmoid_f := 787;
        ELSIF x =- 962 THEN
            sigmoid_f := 787;
        ELSIF x =- 961 THEN
            sigmoid_f := 787;
        ELSIF x =- 960 THEN
            sigmoid_f := 787;
        ELSIF x =- 959 THEN
            sigmoid_f := 788;
        ELSIF x =- 958 THEN
            sigmoid_f := 788;
        ELSIF x =- 957 THEN
            sigmoid_f := 788;
        ELSIF x =- 956 THEN
            sigmoid_f := 788;
        ELSIF x =- 955 THEN
            sigmoid_f := 789;
        ELSIF x =- 954 THEN
            sigmoid_f := 789;
        ELSIF x =- 953 THEN
            sigmoid_f := 789;
        ELSIF x =- 952 THEN
            sigmoid_f := 789;
        ELSIF x =- 951 THEN
            sigmoid_f := 790;
        ELSIF x =- 950 THEN
            sigmoid_f := 790;
        ELSIF x =- 949 THEN
            sigmoid_f := 790;
        ELSIF x =- 948 THEN
            sigmoid_f := 790;
        ELSIF x =- 947 THEN
            sigmoid_f := 791;
        ELSIF x =- 946 THEN
            sigmoid_f := 791;
        ELSIF x =- 945 THEN
            sigmoid_f := 791;
        ELSIF x =- 944 THEN
            sigmoid_f := 791;
        ELSIF x =- 943 THEN
            sigmoid_f := 792;
        ELSIF x =- 942 THEN
            sigmoid_f := 792;
        ELSIF x =- 941 THEN
            sigmoid_f := 792;
        ELSIF x =- 940 THEN
            sigmoid_f := 792;
        ELSIF x =- 939 THEN
            sigmoid_f := 793;
        ELSIF x =- 938 THEN
            sigmoid_f := 793;
        ELSIF x =- 937 THEN
            sigmoid_f := 793;
        ELSIF x =- 936 THEN
            sigmoid_f := 793;
        ELSIF x =- 935 THEN
            sigmoid_f := 794;
        ELSIF x =- 934 THEN
            sigmoid_f := 794;
        ELSIF x =- 933 THEN
            sigmoid_f := 794;
        ELSIF x =- 932 THEN
            sigmoid_f := 794;
        ELSIF x =- 931 THEN
            sigmoid_f := 794;
        ELSIF x =- 930 THEN
            sigmoid_f := 795;
        ELSIF x =- 929 THEN
            sigmoid_f := 795;
        ELSIF x =- 928 THEN
            sigmoid_f := 795;
        ELSIF x =- 927 THEN
            sigmoid_f := 795;
        ELSIF x =- 926 THEN
            sigmoid_f := 796;
        ELSIF x =- 925 THEN
            sigmoid_f := 796;
        ELSIF x =- 924 THEN
            sigmoid_f := 796;
        ELSIF x =- 923 THEN
            sigmoid_f := 796;
        ELSIF x =- 922 THEN
            sigmoid_f := 797;
        ELSIF x =- 921 THEN
            sigmoid_f := 797;
        ELSIF x =- 920 THEN
            sigmoid_f := 797;
        ELSIF x =- 919 THEN
            sigmoid_f := 797;
        ELSIF x =- 918 THEN
            sigmoid_f := 798;
        ELSIF x =- 917 THEN
            sigmoid_f := 798;
        ELSIF x =- 916 THEN
            sigmoid_f := 798;
        ELSIF x =- 915 THEN
            sigmoid_f := 798;
        ELSIF x =- 914 THEN
            sigmoid_f := 799;
        ELSIF x =- 913 THEN
            sigmoid_f := 799;
        ELSIF x =- 912 THEN
            sigmoid_f := 799;
        ELSIF x =- 911 THEN
            sigmoid_f := 799;
        ELSIF x =- 910 THEN
            sigmoid_f := 800;
        ELSIF x =- 909 THEN
            sigmoid_f := 800;
        ELSIF x =- 908 THEN
            sigmoid_f := 800;
        ELSIF x =- 907 THEN
            sigmoid_f := 800;
        ELSIF x =- 906 THEN
            sigmoid_f := 801;
        ELSIF x =- 905 THEN
            sigmoid_f := 801;
        ELSIF x =- 904 THEN
            sigmoid_f := 801;
        ELSIF x =- 903 THEN
            sigmoid_f := 801;
        ELSIF x =- 902 THEN
            sigmoid_f := 801;
        ELSIF x =- 901 THEN
            sigmoid_f := 802;
        ELSIF x =- 900 THEN
            sigmoid_f := 802;
        ELSIF x =- 899 THEN
            sigmoid_f := 802;
        ELSIF x =- 898 THEN
            sigmoid_f := 802;
        ELSIF x =- 897 THEN
            sigmoid_f := 803;
        ELSIF x =- 896 THEN
            sigmoid_f := 803;
        ELSIF x =- 895 THEN
            sigmoid_f := 803;
        ELSIF x =- 894 THEN
            sigmoid_f := 803;
        ELSIF x =- 893 THEN
            sigmoid_f := 804;
        ELSIF x =- 892 THEN
            sigmoid_f := 804;
        ELSIF x =- 891 THEN
            sigmoid_f := 804;
        ELSIF x =- 890 THEN
            sigmoid_f := 804;
        ELSIF x =- 889 THEN
            sigmoid_f := 805;
        ELSIF x =- 888 THEN
            sigmoid_f := 805;
        ELSIF x =- 887 THEN
            sigmoid_f := 805;
        ELSIF x =- 886 THEN
            sigmoid_f := 805;
        ELSIF x =- 885 THEN
            sigmoid_f := 806;
        ELSIF x =- 884 THEN
            sigmoid_f := 806;
        ELSIF x =- 883 THEN
            sigmoid_f := 806;
        ELSIF x =- 882 THEN
            sigmoid_f := 806;
        ELSIF x =- 881 THEN
            sigmoid_f := 807;
        ELSIF x =- 880 THEN
            sigmoid_f := 807;
        ELSIF x =- 879 THEN
            sigmoid_f := 807;
        ELSIF x =- 878 THEN
            sigmoid_f := 807;
        ELSIF x =- 877 THEN
            sigmoid_f := 808;
        ELSIF x =- 876 THEN
            sigmoid_f := 808;
        ELSIF x =- 875 THEN
            sigmoid_f := 808;
        ELSIF x =- 874 THEN
            sigmoid_f := 808;
        ELSIF x =- 873 THEN
            sigmoid_f := 808;
        ELSIF x =- 872 THEN
            sigmoid_f := 809;
        ELSIF x =- 871 THEN
            sigmoid_f := 809;
        ELSIF x =- 870 THEN
            sigmoid_f := 809;
        ELSIF x =- 869 THEN
            sigmoid_f := 809;
        ELSIF x =- 868 THEN
            sigmoid_f := 810;
        ELSIF x =- 867 THEN
            sigmoid_f := 810;
        ELSIF x =- 866 THEN
            sigmoid_f := 810;
        ELSIF x =- 865 THEN
            sigmoid_f := 810;
        ELSIF x =- 864 THEN
            sigmoid_f := 811;
        ELSIF x =- 863 THEN
            sigmoid_f := 811;
        ELSIF x =- 862 THEN
            sigmoid_f := 811;
        ELSIF x =- 861 THEN
            sigmoid_f := 811;
        ELSIF x =- 860 THEN
            sigmoid_f := 812;
        ELSIF x =- 859 THEN
            sigmoid_f := 812;
        ELSIF x =- 858 THEN
            sigmoid_f := 812;
        ELSIF x =- 857 THEN
            sigmoid_f := 812;
        ELSIF x =- 856 THEN
            sigmoid_f := 813;
        ELSIF x =- 855 THEN
            sigmoid_f := 813;
        ELSIF x =- 854 THEN
            sigmoid_f := 813;
        ELSIF x =- 853 THEN
            sigmoid_f := 813;
        ELSIF x =- 852 THEN
            sigmoid_f := 814;
        ELSIF x =- 851 THEN
            sigmoid_f := 814;
        ELSIF x =- 850 THEN
            sigmoid_f := 814;
        ELSIF x =- 849 THEN
            sigmoid_f := 814;
        ELSIF x =- 848 THEN
            sigmoid_f := 815;
        ELSIF x =- 847 THEN
            sigmoid_f := 815;
        ELSIF x =- 846 THEN
            sigmoid_f := 815;
        ELSIF x =- 845 THEN
            sigmoid_f := 815;
        ELSIF x =- 844 THEN
            sigmoid_f := 816;
        ELSIF x =- 843 THEN
            sigmoid_f := 816;
        ELSIF x =- 842 THEN
            sigmoid_f := 816;
        ELSIF x =- 841 THEN
            sigmoid_f := 816;
        ELSIF x =- 840 THEN
            sigmoid_f := 816;
        ELSIF x =- 839 THEN
            sigmoid_f := 817;
        ELSIF x =- 838 THEN
            sigmoid_f := 817;
        ELSIF x =- 837 THEN
            sigmoid_f := 817;
        ELSIF x =- 836 THEN
            sigmoid_f := 817;
        ELSIF x =- 835 THEN
            sigmoid_f := 818;
        ELSIF x =- 834 THEN
            sigmoid_f := 818;
        ELSIF x =- 833 THEN
            sigmoid_f := 818;
        ELSIF x =- 832 THEN
            sigmoid_f := 818;
        ELSIF x =- 831 THEN
            sigmoid_f := 819;
        ELSIF x =- 830 THEN
            sigmoid_f := 819;
        ELSIF x =- 829 THEN
            sigmoid_f := 819;
        ELSIF x =- 828 THEN
            sigmoid_f := 819;
        ELSIF x =- 827 THEN
            sigmoid_f := 820;
        ELSIF x =- 826 THEN
            sigmoid_f := 820;
        ELSIF x =- 825 THEN
            sigmoid_f := 820;
        ELSIF x =- 824 THEN
            sigmoid_f := 820;
        ELSIF x =- 823 THEN
            sigmoid_f := 821;
        ELSIF x =- 822 THEN
            sigmoid_f := 821;
        ELSIF x =- 821 THEN
            sigmoid_f := 821;
        ELSIF x =- 820 THEN
            sigmoid_f := 821;
        ELSIF x =- 819 THEN
            sigmoid_f := 822;
        ELSIF x =- 818 THEN
            sigmoid_f := 822;
        ELSIF x =- 817 THEN
            sigmoid_f := 822;
        ELSIF x =- 816 THEN
            sigmoid_f := 822;
        ELSIF x =- 815 THEN
            sigmoid_f := 823;
        ELSIF x =- 814 THEN
            sigmoid_f := 823;
        ELSIF x =- 813 THEN
            sigmoid_f := 823;
        ELSIF x =- 812 THEN
            sigmoid_f := 823;
        ELSIF x =- 811 THEN
            sigmoid_f := 823;
        ELSIF x =- 810 THEN
            sigmoid_f := 824;
        ELSIF x =- 809 THEN
            sigmoid_f := 824;
        ELSIF x =- 808 THEN
            sigmoid_f := 824;
        ELSIF x =- 807 THEN
            sigmoid_f := 824;
        ELSIF x =- 806 THEN
            sigmoid_f := 825;
        ELSIF x =- 805 THEN
            sigmoid_f := 825;
        ELSIF x =- 804 THEN
            sigmoid_f := 825;
        ELSIF x =- 803 THEN
            sigmoid_f := 825;
        ELSIF x =- 802 THEN
            sigmoid_f := 826;
        ELSIF x =- 801 THEN
            sigmoid_f := 826;
        ELSIF x =- 800 THEN
            sigmoid_f := 826;
        ELSIF x =- 799 THEN
            sigmoid_f := 826;
        ELSIF x =- 798 THEN
            sigmoid_f := 827;
        ELSIF x =- 797 THEN
            sigmoid_f := 827;
        ELSIF x =- 796 THEN
            sigmoid_f := 827;
        ELSIF x =- 795 THEN
            sigmoid_f := 827;
        ELSIF x =- 794 THEN
            sigmoid_f := 828;
        ELSIF x =- 793 THEN
            sigmoid_f := 828;
        ELSIF x =- 792 THEN
            sigmoid_f := 828;
        ELSIF x =- 791 THEN
            sigmoid_f := 828;
        ELSIF x =- 790 THEN
            sigmoid_f := 829;
        ELSIF x =- 789 THEN
            sigmoid_f := 829;
        ELSIF x =- 788 THEN
            sigmoid_f := 829;
        ELSIF x =- 787 THEN
            sigmoid_f := 829;
        ELSIF x =- 786 THEN
            sigmoid_f := 830;
        ELSIF x =- 785 THEN
            sigmoid_f := 830;
        ELSIF x =- 784 THEN
            sigmoid_f := 830;
        ELSIF x =- 783 THEN
            sigmoid_f := 830;
        ELSIF x =- 782 THEN
            sigmoid_f := 830;
        ELSIF x =- 781 THEN
            sigmoid_f := 831;
        ELSIF x =- 780 THEN
            sigmoid_f := 831;
        ELSIF x =- 779 THEN
            sigmoid_f := 831;
        ELSIF x =- 778 THEN
            sigmoid_f := 831;
        ELSIF x =- 777 THEN
            sigmoid_f := 832;
        ELSIF x =- 776 THEN
            sigmoid_f := 832;
        ELSIF x =- 775 THEN
            sigmoid_f := 832;
        ELSIF x =- 774 THEN
            sigmoid_f := 832;
        ELSIF x =- 773 THEN
            sigmoid_f := 833;
        ELSIF x =- 772 THEN
            sigmoid_f := 833;
        ELSIF x =- 771 THEN
            sigmoid_f := 833;
        ELSIF x =- 770 THEN
            sigmoid_f := 833;
        ELSIF x =- 769 THEN
            sigmoid_f := 834;
        ELSIF x =- 768 THEN
            sigmoid_f := 834;
        ELSIF x =- 767 THEN
            sigmoid_f := 834;
        ELSIF x =- 766 THEN
            sigmoid_f := 834;
        ELSIF x =- 765 THEN
            sigmoid_f := 835;
        ELSIF x =- 764 THEN
            sigmoid_f := 835;
        ELSIF x =- 763 THEN
            sigmoid_f := 835;
        ELSIF x =- 762 THEN
            sigmoid_f := 835;
        ELSIF x =- 761 THEN
            sigmoid_f := 836;
        ELSIF x =- 760 THEN
            sigmoid_f := 836;
        ELSIF x =- 759 THEN
            sigmoid_f := 836;
        ELSIF x =- 758 THEN
            sigmoid_f := 836;
        ELSIF x =- 757 THEN
            sigmoid_f := 837;
        ELSIF x =- 756 THEN
            sigmoid_f := 837;
        ELSIF x =- 755 THEN
            sigmoid_f := 837;
        ELSIF x =- 754 THEN
            sigmoid_f := 837;
        ELSIF x =- 753 THEN
            sigmoid_f := 838;
        ELSIF x =- 752 THEN
            sigmoid_f := 838;
        ELSIF x =- 751 THEN
            sigmoid_f := 838;
        ELSIF x =- 750 THEN
            sigmoid_f := 838;
        ELSIF x =- 749 THEN
            sigmoid_f := 838;
        ELSIF x =- 748 THEN
            sigmoid_f := 839;
        ELSIF x =- 747 THEN
            sigmoid_f := 839;
        ELSIF x =- 746 THEN
            sigmoid_f := 839;
        ELSIF x =- 745 THEN
            sigmoid_f := 839;
        ELSIF x =- 744 THEN
            sigmoid_f := 840;
        ELSIF x =- 743 THEN
            sigmoid_f := 840;
        ELSIF x =- 742 THEN
            sigmoid_f := 840;
        ELSIF x =- 741 THEN
            sigmoid_f := 840;
        ELSIF x =- 740 THEN
            sigmoid_f := 841;
        ELSIF x =- 739 THEN
            sigmoid_f := 841;
        ELSIF x =- 738 THEN
            sigmoid_f := 841;
        ELSIF x =- 737 THEN
            sigmoid_f := 841;
        ELSIF x =- 736 THEN
            sigmoid_f := 842;
        ELSIF x =- 735 THEN
            sigmoid_f := 842;
        ELSIF x =- 734 THEN
            sigmoid_f := 842;
        ELSIF x =- 733 THEN
            sigmoid_f := 842;
        ELSIF x =- 732 THEN
            sigmoid_f := 843;
        ELSIF x =- 731 THEN
            sigmoid_f := 843;
        ELSIF x =- 730 THEN
            sigmoid_f := 843;
        ELSIF x =- 729 THEN
            sigmoid_f := 843;
        ELSIF x =- 728 THEN
            sigmoid_f := 844;
        ELSIF x =- 727 THEN
            sigmoid_f := 844;
        ELSIF x =- 726 THEN
            sigmoid_f := 844;
        ELSIF x =- 725 THEN
            sigmoid_f := 844;
        ELSIF x =- 724 THEN
            sigmoid_f := 845;
        ELSIF x =- 723 THEN
            sigmoid_f := 845;
        ELSIF x =- 722 THEN
            sigmoid_f := 845;
        ELSIF x =- 721 THEN
            sigmoid_f := 845;
        ELSIF x =- 720 THEN
            sigmoid_f := 845;
        ELSIF x =- 719 THEN
            sigmoid_f := 846;
        ELSIF x =- 718 THEN
            sigmoid_f := 846;
        ELSIF x =- 717 THEN
            sigmoid_f := 846;
        ELSIF x =- 716 THEN
            sigmoid_f := 846;
        ELSIF x =- 715 THEN
            sigmoid_f := 847;
        ELSIF x =- 714 THEN
            sigmoid_f := 847;
        ELSIF x =- 713 THEN
            sigmoid_f := 847;
        ELSIF x =- 712 THEN
            sigmoid_f := 847;
        ELSIF x =- 711 THEN
            sigmoid_f := 848;
        ELSIF x =- 710 THEN
            sigmoid_f := 848;
        ELSIF x =- 709 THEN
            sigmoid_f := 848;
        ELSIF x =- 708 THEN
            sigmoid_f := 848;
        ELSIF x =- 707 THEN
            sigmoid_f := 849;
        ELSIF x =- 706 THEN
            sigmoid_f := 849;
        ELSIF x =- 705 THEN
            sigmoid_f := 849;
        ELSIF x =- 704 THEN
            sigmoid_f := 849;
        ELSIF x =- 703 THEN
            sigmoid_f := 850;
        ELSIF x =- 702 THEN
            sigmoid_f := 850;
        ELSIF x =- 701 THEN
            sigmoid_f := 850;
        ELSIF x =- 700 THEN
            sigmoid_f := 850;
        ELSIF x =- 699 THEN
            sigmoid_f := 851;
        ELSIF x =- 698 THEN
            sigmoid_f := 851;
        ELSIF x =- 697 THEN
            sigmoid_f := 851;
        ELSIF x =- 696 THEN
            sigmoid_f := 851;
        ELSIF x =- 695 THEN
            sigmoid_f := 852;
        ELSIF x =- 694 THEN
            sigmoid_f := 852;
        ELSIF x =- 693 THEN
            sigmoid_f := 852;
        ELSIF x =- 692 THEN
            sigmoid_f := 852;
        ELSIF x =- 691 THEN
            sigmoid_f := 852;
        ELSIF x =- 690 THEN
            sigmoid_f := 853;
        ELSIF x =- 689 THEN
            sigmoid_f := 853;
        ELSIF x =- 688 THEN
            sigmoid_f := 853;
        ELSIF x =- 687 THEN
            sigmoid_f := 853;
        ELSIF x =- 686 THEN
            sigmoid_f := 854;
        ELSIF x =- 685 THEN
            sigmoid_f := 854;
        ELSIF x =- 684 THEN
            sigmoid_f := 854;
        ELSIF x =- 683 THEN
            sigmoid_f := 854;
        ELSIF x =- 682 THEN
            sigmoid_f := 855;
        ELSIF x =- 681 THEN
            sigmoid_f := 855;
        ELSIF x =- 680 THEN
            sigmoid_f := 855;
        ELSIF x =- 679 THEN
            sigmoid_f := 855;
        ELSIF x =- 678 THEN
            sigmoid_f := 856;
        ELSIF x =- 677 THEN
            sigmoid_f := 856;
        ELSIF x =- 676 THEN
            sigmoid_f := 856;
        ELSIF x =- 675 THEN
            sigmoid_f := 856;
        ELSIF x =- 674 THEN
            sigmoid_f := 857;
        ELSIF x =- 673 THEN
            sigmoid_f := 857;
        ELSIF x =- 672 THEN
            sigmoid_f := 857;
        ELSIF x =- 671 THEN
            sigmoid_f := 857;
        ELSIF x =- 670 THEN
            sigmoid_f := 858;
        ELSIF x =- 669 THEN
            sigmoid_f := 858;
        ELSIF x =- 668 THEN
            sigmoid_f := 858;
        ELSIF x =- 667 THEN
            sigmoid_f := 858;
        ELSIF x =- 666 THEN
            sigmoid_f := 859;
        ELSIF x =- 665 THEN
            sigmoid_f := 859;
        ELSIF x =- 664 THEN
            sigmoid_f := 859;
        ELSIF x =- 663 THEN
            sigmoid_f := 859;
        ELSIF x =- 662 THEN
            sigmoid_f := 859;
        ELSIF x =- 661 THEN
            sigmoid_f := 860;
        ELSIF x =- 660 THEN
            sigmoid_f := 860;
        ELSIF x =- 659 THEN
            sigmoid_f := 860;
        ELSIF x =- 658 THEN
            sigmoid_f := 860;
        ELSIF x =- 657 THEN
            sigmoid_f := 861;
        ELSIF x =- 656 THEN
            sigmoid_f := 861;
        ELSIF x =- 655 THEN
            sigmoid_f := 861;
        ELSIF x =- 654 THEN
            sigmoid_f := 861;
        ELSIF x =- 653 THEN
            sigmoid_f := 862;
        ELSIF x =- 652 THEN
            sigmoid_f := 862;
        ELSIF x =- 651 THEN
            sigmoid_f := 862;
        ELSIF x =- 650 THEN
            sigmoid_f := 862;
        ELSIF x =- 649 THEN
            sigmoid_f := 863;
        ELSIF x =- 648 THEN
            sigmoid_f := 863;
        ELSIF x =- 647 THEN
            sigmoid_f := 863;
        ELSIF x =- 646 THEN
            sigmoid_f := 863;
        ELSIF x =- 645 THEN
            sigmoid_f := 864;
        ELSIF x =- 644 THEN
            sigmoid_f := 864;
        ELSIF x =- 643 THEN
            sigmoid_f := 864;
        ELSIF x =- 642 THEN
            sigmoid_f := 864;
        ELSIF x =- 641 THEN
            sigmoid_f := 865;
        ELSIF x =- 640 THEN
            sigmoid_f := 865;
        ELSIF x =- 639 THEN
            sigmoid_f := 865;
        ELSIF x =- 638 THEN
            sigmoid_f := 865;
        ELSIF x =- 637 THEN
            sigmoid_f := 866;
        ELSIF x =- 636 THEN
            sigmoid_f := 866;
        ELSIF x =- 635 THEN
            sigmoid_f := 866;
        ELSIF x =- 634 THEN
            sigmoid_f := 866;
        ELSIF x =- 633 THEN
            sigmoid_f := 867;
        ELSIF x =- 632 THEN
            sigmoid_f := 867;
        ELSIF x =- 631 THEN
            sigmoid_f := 867;
        ELSIF x =- 630 THEN
            sigmoid_f := 867;
        ELSIF x =- 629 THEN
            sigmoid_f := 867;
        ELSIF x =- 628 THEN
            sigmoid_f := 868;
        ELSIF x =- 627 THEN
            sigmoid_f := 868;
        ELSIF x =- 626 THEN
            sigmoid_f := 868;
        ELSIF x =- 625 THEN
            sigmoid_f := 868;
        ELSIF x =- 624 THEN
            sigmoid_f := 869;
        ELSIF x =- 623 THEN
            sigmoid_f := 869;
        ELSIF x =- 622 THEN
            sigmoid_f := 869;
        ELSIF x =- 621 THEN
            sigmoid_f := 869;
        ELSIF x =- 620 THEN
            sigmoid_f := 870;
        ELSIF x =- 619 THEN
            sigmoid_f := 870;
        ELSIF x =- 618 THEN
            sigmoid_f := 870;
        ELSIF x =- 617 THEN
            sigmoid_f := 870;
        ELSIF x =- 616 THEN
            sigmoid_f := 871;
        ELSIF x =- 615 THEN
            sigmoid_f := 871;
        ELSIF x =- 614 THEN
            sigmoid_f := 871;
        ELSIF x =- 613 THEN
            sigmoid_f := 871;
        ELSIF x =- 612 THEN
            sigmoid_f := 872;
        ELSIF x =- 611 THEN
            sigmoid_f := 872;
        ELSIF x =- 610 THEN
            sigmoid_f := 872;
        ELSIF x =- 609 THEN
            sigmoid_f := 872;
        ELSIF x =- 608 THEN
            sigmoid_f := 873;
        ELSIF x =- 607 THEN
            sigmoid_f := 873;
        ELSIF x =- 606 THEN
            sigmoid_f := 873;
        ELSIF x =- 605 THEN
            sigmoid_f := 873;
        ELSIF x =- 604 THEN
            sigmoid_f := 874;
        ELSIF x =- 603 THEN
            sigmoid_f := 874;
        ELSIF x =- 602 THEN
            sigmoid_f := 874;
        ELSIF x =- 601 THEN
            sigmoid_f := 874;
        ELSIF x =- 600 THEN
            sigmoid_f := 874;
        ELSIF x =- 599 THEN
            sigmoid_f := 875;
        ELSIF x =- 598 THEN
            sigmoid_f := 875;
        ELSIF x =- 597 THEN
            sigmoid_f := 875;
        ELSIF x =- 596 THEN
            sigmoid_f := 875;
        ELSIF x =- 595 THEN
            sigmoid_f := 876;
        ELSIF x =- 594 THEN
            sigmoid_f := 876;
        ELSIF x =- 593 THEN
            sigmoid_f := 876;
        ELSIF x =- 592 THEN
            sigmoid_f := 876;
        ELSIF x =- 591 THEN
            sigmoid_f := 877;
        ELSIF x =- 590 THEN
            sigmoid_f := 877;
        ELSIF x =- 589 THEN
            sigmoid_f := 877;
        ELSIF x =- 588 THEN
            sigmoid_f := 877;
        ELSIF x =- 587 THEN
            sigmoid_f := 878;
        ELSIF x =- 586 THEN
            sigmoid_f := 878;
        ELSIF x =- 585 THEN
            sigmoid_f := 878;
        ELSIF x =- 584 THEN
            sigmoid_f := 878;
        ELSIF x =- 583 THEN
            sigmoid_f := 879;
        ELSIF x =- 582 THEN
            sigmoid_f := 879;
        ELSIF x =- 581 THEN
            sigmoid_f := 879;
        ELSIF x =- 580 THEN
            sigmoid_f := 879;
        ELSIF x =- 579 THEN
            sigmoid_f := 880;
        ELSIF x =- 578 THEN
            sigmoid_f := 880;
        ELSIF x =- 577 THEN
            sigmoid_f := 880;
        ELSIF x =- 576 THEN
            sigmoid_f := 880;
        ELSIF x =- 575 THEN
            sigmoid_f := 881;
        ELSIF x =- 574 THEN
            sigmoid_f := 881;
        ELSIF x =- 573 THEN
            sigmoid_f := 881;
        ELSIF x =- 572 THEN
            sigmoid_f := 881;
        ELSIF x =- 571 THEN
            sigmoid_f := 881;
        ELSIF x =- 570 THEN
            sigmoid_f := 882;
        ELSIF x =- 569 THEN
            sigmoid_f := 882;
        ELSIF x =- 568 THEN
            sigmoid_f := 882;
        ELSIF x =- 567 THEN
            sigmoid_f := 882;
        ELSIF x =- 566 THEN
            sigmoid_f := 883;
        ELSIF x =- 565 THEN
            sigmoid_f := 883;
        ELSIF x =- 564 THEN
            sigmoid_f := 883;
        ELSIF x =- 563 THEN
            sigmoid_f := 883;
        ELSIF x =- 562 THEN
            sigmoid_f := 884;
        ELSIF x =- 561 THEN
            sigmoid_f := 884;
        ELSIF x =- 560 THEN
            sigmoid_f := 884;
        ELSIF x =- 559 THEN
            sigmoid_f := 884;
        ELSIF x =- 558 THEN
            sigmoid_f := 885;
        ELSIF x =- 557 THEN
            sigmoid_f := 885;
        ELSIF x =- 556 THEN
            sigmoid_f := 885;
        ELSIF x =- 555 THEN
            sigmoid_f := 885;
        ELSIF x =- 554 THEN
            sigmoid_f := 886;
        ELSIF x =- 553 THEN
            sigmoid_f := 886;
        ELSIF x =- 552 THEN
            sigmoid_f := 886;
        ELSIF x =- 551 THEN
            sigmoid_f := 886;
        ELSIF x =- 550 THEN
            sigmoid_f := 887;
        ELSIF x =- 549 THEN
            sigmoid_f := 887;
        ELSIF x =- 548 THEN
            sigmoid_f := 887;
        ELSIF x =- 547 THEN
            sigmoid_f := 887;
        ELSIF x =- 546 THEN
            sigmoid_f := 888;
        ELSIF x =- 545 THEN
            sigmoid_f := 888;
        ELSIF x =- 544 THEN
            sigmoid_f := 888;
        ELSIF x =- 543 THEN
            sigmoid_f := 888;
        ELSIF x =- 542 THEN
            sigmoid_f := 888;
        ELSIF x =- 541 THEN
            sigmoid_f := 889;
        ELSIF x =- 540 THEN
            sigmoid_f := 889;
        ELSIF x =- 539 THEN
            sigmoid_f := 889;
        ELSIF x =- 538 THEN
            sigmoid_f := 889;
        ELSIF x =- 537 THEN
            sigmoid_f := 890;
        ELSIF x =- 536 THEN
            sigmoid_f := 890;
        ELSIF x =- 535 THEN
            sigmoid_f := 890;
        ELSIF x =- 534 THEN
            sigmoid_f := 890;
        ELSIF x =- 533 THEN
            sigmoid_f := 891;
        ELSIF x =- 532 THEN
            sigmoid_f := 891;
        ELSIF x =- 531 THEN
            sigmoid_f := 891;
        ELSIF x =- 530 THEN
            sigmoid_f := 891;
        ELSIF x =- 529 THEN
            sigmoid_f := 892;
        ELSIF x =- 528 THEN
            sigmoid_f := 892;
        ELSIF x =- 527 THEN
            sigmoid_f := 892;
        ELSIF x =- 526 THEN
            sigmoid_f := 892;
        ELSIF x =- 525 THEN
            sigmoid_f := 893;
        ELSIF x =- 524 THEN
            sigmoid_f := 893;
        ELSIF x =- 523 THEN
            sigmoid_f := 893;
        ELSIF x =- 522 THEN
            sigmoid_f := 893;
        ELSIF x =- 521 THEN
            sigmoid_f := 894;
        ELSIF x =- 520 THEN
            sigmoid_f := 894;
        ELSIF x =- 519 THEN
            sigmoid_f := 894;
        ELSIF x =- 518 THEN
            sigmoid_f := 894;
        ELSIF x =- 517 THEN
            sigmoid_f := 895;
        ELSIF x =- 516 THEN
            sigmoid_f := 895;
        ELSIF x =- 515 THEN
            sigmoid_f := 895;
        ELSIF x =- 514 THEN
            sigmoid_f := 895;
        ELSIF x =- 513 THEN
            sigmoid_f := 896;
        ELSIF x =- 512 THEN
            sigmoid_f := 896;
        ELSIF x =- 511 THEN
            sigmoid_f := 896;
        ELSIF x =- 510 THEN
            sigmoid_f := 896;
        ELSIF x =- 509 THEN
            sigmoid_f := 896;
        ELSIF x =- 508 THEN
            sigmoid_f := 897;
        ELSIF x =- 507 THEN
            sigmoid_f := 897;
        ELSIF x =- 506 THEN
            sigmoid_f := 897;
        ELSIF x =- 505 THEN
            sigmoid_f := 897;
        ELSIF x =- 504 THEN
            sigmoid_f := 898;
        ELSIF x =- 503 THEN
            sigmoid_f := 898;
        ELSIF x =- 502 THEN
            sigmoid_f := 898;
        ELSIF x =- 501 THEN
            sigmoid_f := 898;
        ELSIF x =- 500 THEN
            sigmoid_f := 899;
        ELSIF x =- 499 THEN
            sigmoid_f := 899;
        ELSIF x =- 498 THEN
            sigmoid_f := 899;
        ELSIF x =- 497 THEN
            sigmoid_f := 899;
        ELSIF x =- 496 THEN
            sigmoid_f := 900;
        ELSIF x =- 495 THEN
            sigmoid_f := 900;
        ELSIF x =- 494 THEN
            sigmoid_f := 900;
        ELSIF x =- 493 THEN
            sigmoid_f := 900;
        ELSIF x =- 492 THEN
            sigmoid_f := 901;
        ELSIF x =- 491 THEN
            sigmoid_f := 901;
        ELSIF x =- 490 THEN
            sigmoid_f := 901;
        ELSIF x =- 489 THEN
            sigmoid_f := 901;
        ELSIF x =- 488 THEN
            sigmoid_f := 902;
        ELSIF x =- 487 THEN
            sigmoid_f := 902;
        ELSIF x =- 486 THEN
            sigmoid_f := 902;
        ELSIF x =- 485 THEN
            sigmoid_f := 902;
        ELSIF x =- 484 THEN
            sigmoid_f := 903;
        ELSIF x =- 483 THEN
            sigmoid_f := 903;
        ELSIF x =- 482 THEN
            sigmoid_f := 903;
        ELSIF x =- 481 THEN
            sigmoid_f := 903;
        ELSIF x =- 480 THEN
            sigmoid_f := 904;
        ELSIF x =- 479 THEN
            sigmoid_f := 904;
        ELSIF x =- 478 THEN
            sigmoid_f := 904;
        ELSIF x =- 477 THEN
            sigmoid_f := 904;
        ELSIF x =- 476 THEN
            sigmoid_f := 905;
        ELSIF x =- 475 THEN
            sigmoid_f := 905;
        ELSIF x =- 474 THEN
            sigmoid_f := 905;
        ELSIF x =- 473 THEN
            sigmoid_f := 905;
        ELSIF x =- 472 THEN
            sigmoid_f := 906;
        ELSIF x =- 471 THEN
            sigmoid_f := 906;
        ELSIF x =- 470 THEN
            sigmoid_f := 906;
        ELSIF x =- 469 THEN
            sigmoid_f := 906;
        ELSIF x =- 468 THEN
            sigmoid_f := 907;
        ELSIF x =- 467 THEN
            sigmoid_f := 907;
        ELSIF x =- 466 THEN
            sigmoid_f := 907;
        ELSIF x =- 465 THEN
            sigmoid_f := 907;
        ELSIF x =- 464 THEN
            sigmoid_f := 908;
        ELSIF x =- 463 THEN
            sigmoid_f := 908;
        ELSIF x =- 462 THEN
            sigmoid_f := 908;
        ELSIF x =- 461 THEN
            sigmoid_f := 908;
        ELSIF x =- 460 THEN
            sigmoid_f := 909;
        ELSIF x =- 459 THEN
            sigmoid_f := 909;
        ELSIF x =- 458 THEN
            sigmoid_f := 909;
        ELSIF x =- 457 THEN
            sigmoid_f := 909;
        ELSIF x =- 456 THEN
            sigmoid_f := 910;
        ELSIF x =- 455 THEN
            sigmoid_f := 910;
        ELSIF x =- 454 THEN
            sigmoid_f := 910;
        ELSIF x =- 453 THEN
            sigmoid_f := 910;
        ELSIF x =- 452 THEN
            sigmoid_f := 911;
        ELSIF x =- 451 THEN
            sigmoid_f := 911;
        ELSIF x =- 450 THEN
            sigmoid_f := 911;
        ELSIF x =- 449 THEN
            sigmoid_f := 911;
        ELSIF x =- 448 THEN
            sigmoid_f := 912;
        ELSIF x =- 447 THEN
            sigmoid_f := 912;
        ELSIF x =- 446 THEN
            sigmoid_f := 912;
        ELSIF x =- 445 THEN
            sigmoid_f := 912;
        ELSIF x =- 444 THEN
            sigmoid_f := 913;
        ELSIF x =- 443 THEN
            sigmoid_f := 913;
        ELSIF x =- 442 THEN
            sigmoid_f := 913;
        ELSIF x =- 441 THEN
            sigmoid_f := 913;
        ELSIF x =- 440 THEN
            sigmoid_f := 914;
        ELSIF x =- 439 THEN
            sigmoid_f := 914;
        ELSIF x =- 438 THEN
            sigmoid_f := 914;
        ELSIF x =- 437 THEN
            sigmoid_f := 914;
        ELSIF x =- 436 THEN
            sigmoid_f := 915;
        ELSIF x =- 435 THEN
            sigmoid_f := 915;
        ELSIF x =- 434 THEN
            sigmoid_f := 915;
        ELSIF x =- 433 THEN
            sigmoid_f := 915;
        ELSIF x =- 432 THEN
            sigmoid_f := 916;
        ELSIF x =- 431 THEN
            sigmoid_f := 916;
        ELSIF x =- 430 THEN
            sigmoid_f := 916;
        ELSIF x =- 429 THEN
            sigmoid_f := 916;
        ELSIF x =- 428 THEN
            sigmoid_f := 917;
        ELSIF x =- 427 THEN
            sigmoid_f := 917;
        ELSIF x =- 426 THEN
            sigmoid_f := 917;
        ELSIF x =- 425 THEN
            sigmoid_f := 917;
        ELSIF x =- 424 THEN
            sigmoid_f := 918;
        ELSIF x =- 423 THEN
            sigmoid_f := 918;
        ELSIF x =- 422 THEN
            sigmoid_f := 918;
        ELSIF x =- 421 THEN
            sigmoid_f := 918;
        ELSIF x =- 420 THEN
            sigmoid_f := 919;
        ELSIF x =- 419 THEN
            sigmoid_f := 919;
        ELSIF x =- 418 THEN
            sigmoid_f := 919;
        ELSIF x =- 417 THEN
            sigmoid_f := 919;
        ELSIF x =- 416 THEN
            sigmoid_f := 920;
        ELSIF x =- 415 THEN
            sigmoid_f := 920;
        ELSIF x =- 414 THEN
            sigmoid_f := 920;
        ELSIF x =- 413 THEN
            sigmoid_f := 920;
        ELSIF x =- 412 THEN
            sigmoid_f := 921;
        ELSIF x =- 411 THEN
            sigmoid_f := 921;
        ELSIF x =- 410 THEN
            sigmoid_f := 921;
        ELSIF x =- 409 THEN
            sigmoid_f := 921;
        ELSIF x =- 408 THEN
            sigmoid_f := 922;
        ELSIF x =- 407 THEN
            sigmoid_f := 922;
        ELSIF x =- 406 THEN
            sigmoid_f := 922;
        ELSIF x =- 405 THEN
            sigmoid_f := 922;
        ELSIF x =- 404 THEN
            sigmoid_f := 923;
        ELSIF x =- 403 THEN
            sigmoid_f := 923;
        ELSIF x =- 402 THEN
            sigmoid_f := 923;
        ELSIF x =- 401 THEN
            sigmoid_f := 923;
        ELSIF x =- 400 THEN
            sigmoid_f := 924;
        ELSIF x =- 399 THEN
            sigmoid_f := 924;
        ELSIF x =- 398 THEN
            sigmoid_f := 924;
        ELSIF x =- 397 THEN
            sigmoid_f := 924;
        ELSIF x =- 396 THEN
            sigmoid_f := 925;
        ELSIF x =- 395 THEN
            sigmoid_f := 925;
        ELSIF x =- 394 THEN
            sigmoid_f := 925;
        ELSIF x =- 393 THEN
            sigmoid_f := 925;
        ELSIF x =- 392 THEN
            sigmoid_f := 926;
        ELSIF x =- 391 THEN
            sigmoid_f := 926;
        ELSIF x =- 390 THEN
            sigmoid_f := 926;
        ELSIF x =- 389 THEN
            sigmoid_f := 926;
        ELSIF x =- 388 THEN
            sigmoid_f := 927;
        ELSIF x =- 387 THEN
            sigmoid_f := 927;
        ELSIF x =- 386 THEN
            sigmoid_f := 927;
        ELSIF x =- 385 THEN
            sigmoid_f := 927;
        ELSIF x =- 384 THEN
            sigmoid_f := 928;
        ELSIF x =- 383 THEN
            sigmoid_f := 928;
        ELSIF x =- 382 THEN
            sigmoid_f := 928;
        ELSIF x =- 381 THEN
            sigmoid_f := 928;
        ELSIF x =- 380 THEN
            sigmoid_f := 929;
        ELSIF x =- 379 THEN
            sigmoid_f := 929;
        ELSIF x =- 378 THEN
            sigmoid_f := 929;
        ELSIF x =- 377 THEN
            sigmoid_f := 929;
        ELSIF x =- 376 THEN
            sigmoid_f := 930;
        ELSIF x =- 375 THEN
            sigmoid_f := 930;
        ELSIF x =- 374 THEN
            sigmoid_f := 930;
        ELSIF x =- 373 THEN
            sigmoid_f := 930;
        ELSIF x =- 372 THEN
            sigmoid_f := 931;
        ELSIF x =- 371 THEN
            sigmoid_f := 931;
        ELSIF x =- 370 THEN
            sigmoid_f := 931;
        ELSIF x =- 369 THEN
            sigmoid_f := 931;
        ELSIF x =- 368 THEN
            sigmoid_f := 932;
        ELSIF x =- 367 THEN
            sigmoid_f := 932;
        ELSIF x =- 366 THEN
            sigmoid_f := 932;
        ELSIF x =- 365 THEN
            sigmoid_f := 932;
        ELSIF x =- 364 THEN
            sigmoid_f := 933;
        ELSIF x =- 363 THEN
            sigmoid_f := 933;
        ELSIF x =- 362 THEN
            sigmoid_f := 933;
        ELSIF x =- 361 THEN
            sigmoid_f := 933;
        ELSIF x =- 360 THEN
            sigmoid_f := 934;
        ELSIF x =- 359 THEN
            sigmoid_f := 934;
        ELSIF x =- 358 THEN
            sigmoid_f := 934;
        ELSIF x =- 357 THEN
            sigmoid_f := 934;
        ELSIF x =- 356 THEN
            sigmoid_f := 935;
        ELSIF x =- 355 THEN
            sigmoid_f := 935;
        ELSIF x =- 354 THEN
            sigmoid_f := 935;
        ELSIF x =- 353 THEN
            sigmoid_f := 935;
        ELSIF x =- 352 THEN
            sigmoid_f := 936;
        ELSIF x =- 351 THEN
            sigmoid_f := 936;
        ELSIF x =- 350 THEN
            sigmoid_f := 936;
        ELSIF x =- 349 THEN
            sigmoid_f := 936;
        ELSIF x =- 348 THEN
            sigmoid_f := 937;
        ELSIF x =- 347 THEN
            sigmoid_f := 937;
        ELSIF x =- 346 THEN
            sigmoid_f := 937;
        ELSIF x =- 345 THEN
            sigmoid_f := 937;
        ELSIF x =- 344 THEN
            sigmoid_f := 938;
        ELSIF x =- 343 THEN
            sigmoid_f := 938;
        ELSIF x =- 342 THEN
            sigmoid_f := 938;
        ELSIF x =- 341 THEN
            sigmoid_f := 938;
        ELSIF x =- 340 THEN
            sigmoid_f := 939;
        ELSIF x =- 339 THEN
            sigmoid_f := 939;
        ELSIF x =- 338 THEN
            sigmoid_f := 939;
        ELSIF x =- 337 THEN
            sigmoid_f := 939;
        ELSIF x =- 336 THEN
            sigmoid_f := 940;
        ELSIF x =- 335 THEN
            sigmoid_f := 940;
        ELSIF x =- 334 THEN
            sigmoid_f := 940;
        ELSIF x =- 333 THEN
            sigmoid_f := 940;
        ELSIF x =- 332 THEN
            sigmoid_f := 941;
        ELSIF x =- 331 THEN
            sigmoid_f := 941;
        ELSIF x =- 330 THEN
            sigmoid_f := 941;
        ELSIF x =- 329 THEN
            sigmoid_f := 941;
        ELSIF x =- 328 THEN
            sigmoid_f := 942;
        ELSIF x =- 327 THEN
            sigmoid_f := 942;
        ELSIF x =- 326 THEN
            sigmoid_f := 942;
        ELSIF x =- 325 THEN
            sigmoid_f := 942;
        ELSIF x =- 324 THEN
            sigmoid_f := 943;
        ELSIF x =- 323 THEN
            sigmoid_f := 943;
        ELSIF x =- 322 THEN
            sigmoid_f := 943;
        ELSIF x =- 321 THEN
            sigmoid_f := 943;
        ELSIF x =- 320 THEN
            sigmoid_f := 944;
        ELSIF x =- 319 THEN
            sigmoid_f := 944;
        ELSIF x =- 318 THEN
            sigmoid_f := 944;
        ELSIF x =- 317 THEN
            sigmoid_f := 944;
        ELSIF x =- 316 THEN
            sigmoid_f := 945;
        ELSIF x =- 315 THEN
            sigmoid_f := 945;
        ELSIF x =- 314 THEN
            sigmoid_f := 945;
        ELSIF x =- 313 THEN
            sigmoid_f := 945;
        ELSIF x =- 312 THEN
            sigmoid_f := 946;
        ELSIF x =- 311 THEN
            sigmoid_f := 946;
        ELSIF x =- 310 THEN
            sigmoid_f := 946;
        ELSIF x =- 309 THEN
            sigmoid_f := 946;
        ELSIF x =- 308 THEN
            sigmoid_f := 947;
        ELSIF x =- 307 THEN
            sigmoid_f := 947;
        ELSIF x =- 306 THEN
            sigmoid_f := 947;
        ELSIF x =- 305 THEN
            sigmoid_f := 947;
        ELSIF x =- 304 THEN
            sigmoid_f := 948;
        ELSIF x =- 303 THEN
            sigmoid_f := 948;
        ELSIF x =- 302 THEN
            sigmoid_f := 948;
        ELSIF x =- 301 THEN
            sigmoid_f := 948;
        ELSIF x =- 300 THEN
            sigmoid_f := 949;
        ELSIF x =- 299 THEN
            sigmoid_f := 949;
        ELSIF x =- 298 THEN
            sigmoid_f := 949;
        ELSIF x =- 297 THEN
            sigmoid_f := 949;
        ELSIF x =- 296 THEN
            sigmoid_f := 950;
        ELSIF x =- 295 THEN
            sigmoid_f := 950;
        ELSIF x =- 294 THEN
            sigmoid_f := 950;
        ELSIF x =- 293 THEN
            sigmoid_f := 950;
        ELSIF x =- 292 THEN
            sigmoid_f := 951;
        ELSIF x =- 291 THEN
            sigmoid_f := 951;
        ELSIF x =- 290 THEN
            sigmoid_f := 951;
        ELSIF x =- 289 THEN
            sigmoid_f := 951;
        ELSIF x =- 288 THEN
            sigmoid_f := 952;
        ELSIF x =- 287 THEN
            sigmoid_f := 952;
        ELSIF x =- 286 THEN
            sigmoid_f := 952;
        ELSIF x =- 285 THEN
            sigmoid_f := 952;
        ELSIF x =- 284 THEN
            sigmoid_f := 953;
        ELSIF x =- 283 THEN
            sigmoid_f := 953;
        ELSIF x =- 282 THEN
            sigmoid_f := 953;
        ELSIF x =- 281 THEN
            sigmoid_f := 953;
        ELSIF x =- 280 THEN
            sigmoid_f := 954;
        ELSIF x =- 279 THEN
            sigmoid_f := 954;
        ELSIF x =- 278 THEN
            sigmoid_f := 954;
        ELSIF x =- 277 THEN
            sigmoid_f := 954;
        ELSIF x =- 276 THEN
            sigmoid_f := 955;
        ELSIF x =- 275 THEN
            sigmoid_f := 955;
        ELSIF x =- 274 THEN
            sigmoid_f := 955;
        ELSIF x =- 273 THEN
            sigmoid_f := 955;
        ELSIF x =- 272 THEN
            sigmoid_f := 956;
        ELSIF x =- 271 THEN
            sigmoid_f := 956;
        ELSIF x =- 270 THEN
            sigmoid_f := 956;
        ELSIF x =- 269 THEN
            sigmoid_f := 956;
        ELSIF x =- 268 THEN
            sigmoid_f := 957;
        ELSIF x =- 267 THEN
            sigmoid_f := 957;
        ELSIF x =- 266 THEN
            sigmoid_f := 957;
        ELSIF x =- 265 THEN
            sigmoid_f := 957;
        ELSIF x =- 264 THEN
            sigmoid_f := 958;
        ELSIF x =- 263 THEN
            sigmoid_f := 958;
        ELSIF x =- 262 THEN
            sigmoid_f := 958;
        ELSIF x =- 261 THEN
            sigmoid_f := 958;
        ELSIF x =- 260 THEN
            sigmoid_f := 959;
        ELSIF x =- 259 THEN
            sigmoid_f := 959;
        ELSIF x =- 258 THEN
            sigmoid_f := 959;
        ELSIF x =- 257 THEN
            sigmoid_f := 959;
        ELSIF x =- 256 THEN
            sigmoid_f := 960;
        ELSIF x =- 255 THEN
            sigmoid_f := 960;
        ELSIF x =- 254 THEN
            sigmoid_f := 960;
        ELSIF x =- 253 THEN
            sigmoid_f := 960;
        ELSIF x =- 252 THEN
            sigmoid_f := 961;
        ELSIF x =- 251 THEN
            sigmoid_f := 961;
        ELSIF x =- 250 THEN
            sigmoid_f := 961;
        ELSIF x =- 249 THEN
            sigmoid_f := 961;
        ELSIF x =- 248 THEN
            sigmoid_f := 962;
        ELSIF x =- 247 THEN
            sigmoid_f := 962;
        ELSIF x =- 246 THEN
            sigmoid_f := 962;
        ELSIF x =- 245 THEN
            sigmoid_f := 962;
        ELSIF x =- 244 THEN
            sigmoid_f := 963;
        ELSIF x =- 243 THEN
            sigmoid_f := 963;
        ELSIF x =- 242 THEN
            sigmoid_f := 963;
        ELSIF x =- 241 THEN
            sigmoid_f := 963;
        ELSIF x =- 240 THEN
            sigmoid_f := 964;
        ELSIF x =- 239 THEN
            sigmoid_f := 964;
        ELSIF x =- 238 THEN
            sigmoid_f := 964;
        ELSIF x =- 237 THEN
            sigmoid_f := 964;
        ELSIF x =- 236 THEN
            sigmoid_f := 965;
        ELSIF x =- 235 THEN
            sigmoid_f := 965;
        ELSIF x =- 234 THEN
            sigmoid_f := 965;
        ELSIF x =- 233 THEN
            sigmoid_f := 965;
        ELSIF x =- 232 THEN
            sigmoid_f := 966;
        ELSIF x =- 231 THEN
            sigmoid_f := 966;
        ELSIF x =- 230 THEN
            sigmoid_f := 966;
        ELSIF x =- 229 THEN
            sigmoid_f := 966;
        ELSIF x =- 228 THEN
            sigmoid_f := 967;
        ELSIF x =- 227 THEN
            sigmoid_f := 967;
        ELSIF x =- 226 THEN
            sigmoid_f := 967;
        ELSIF x =- 225 THEN
            sigmoid_f := 967;
        ELSIF x =- 224 THEN
            sigmoid_f := 968;
        ELSIF x =- 223 THEN
            sigmoid_f := 968;
        ELSIF x =- 222 THEN
            sigmoid_f := 968;
        ELSIF x =- 221 THEN
            sigmoid_f := 968;
        ELSIF x =- 220 THEN
            sigmoid_f := 969;
        ELSIF x =- 219 THEN
            sigmoid_f := 969;
        ELSIF x =- 218 THEN
            sigmoid_f := 969;
        ELSIF x =- 217 THEN
            sigmoid_f := 969;
        ELSIF x =- 216 THEN
            sigmoid_f := 970;
        ELSIF x =- 215 THEN
            sigmoid_f := 970;
        ELSIF x =- 214 THEN
            sigmoid_f := 970;
        ELSIF x =- 213 THEN
            sigmoid_f := 970;
        ELSIF x =- 212 THEN
            sigmoid_f := 971;
        ELSIF x =- 211 THEN
            sigmoid_f := 971;
        ELSIF x =- 210 THEN
            sigmoid_f := 971;
        ELSIF x =- 209 THEN
            sigmoid_f := 971;
        ELSIF x =- 208 THEN
            sigmoid_f := 972;
        ELSIF x =- 207 THEN
            sigmoid_f := 972;
        ELSIF x =- 206 THEN
            sigmoid_f := 972;
        ELSIF x =- 205 THEN
            sigmoid_f := 972;
        ELSIF x =- 204 THEN
            sigmoid_f := 973;
        ELSIF x =- 203 THEN
            sigmoid_f := 973;
        ELSIF x =- 202 THEN
            sigmoid_f := 973;
        ELSIF x =- 201 THEN
            sigmoid_f := 973;
        ELSIF x =- 200 THEN
            sigmoid_f := 974;
        ELSIF x =- 199 THEN
            sigmoid_f := 974;
        ELSIF x =- 198 THEN
            sigmoid_f := 974;
        ELSIF x =- 197 THEN
            sigmoid_f := 974;
        ELSIF x =- 196 THEN
            sigmoid_f := 975;
        ELSIF x =- 195 THEN
            sigmoid_f := 975;
        ELSIF x =- 194 THEN
            sigmoid_f := 975;
        ELSIF x =- 193 THEN
            sigmoid_f := 975;
        ELSIF x =- 192 THEN
            sigmoid_f := 976;
        ELSIF x =- 191 THEN
            sigmoid_f := 976;
        ELSIF x =- 190 THEN
            sigmoid_f := 976;
        ELSIF x =- 189 THEN
            sigmoid_f := 976;
        ELSIF x =- 188 THEN
            sigmoid_f := 977;
        ELSIF x =- 187 THEN
            sigmoid_f := 977;
        ELSIF x =- 186 THEN
            sigmoid_f := 977;
        ELSIF x =- 185 THEN
            sigmoid_f := 977;
        ELSIF x =- 184 THEN
            sigmoid_f := 978;
        ELSIF x =- 183 THEN
            sigmoid_f := 978;
        ELSIF x =- 182 THEN
            sigmoid_f := 978;
        ELSIF x =- 181 THEN
            sigmoid_f := 978;
        ELSIF x =- 180 THEN
            sigmoid_f := 979;
        ELSIF x =- 179 THEN
            sigmoid_f := 979;
        ELSIF x =- 178 THEN
            sigmoid_f := 979;
        ELSIF x =- 177 THEN
            sigmoid_f := 979;
        ELSIF x =- 176 THEN
            sigmoid_f := 980;
        ELSIF x =- 175 THEN
            sigmoid_f := 980;
        ELSIF x =- 174 THEN
            sigmoid_f := 980;
        ELSIF x =- 173 THEN
            sigmoid_f := 980;
        ELSIF x =- 172 THEN
            sigmoid_f := 981;
        ELSIF x =- 171 THEN
            sigmoid_f := 981;
        ELSIF x =- 170 THEN
            sigmoid_f := 981;
        ELSIF x =- 169 THEN
            sigmoid_f := 981;
        ELSIF x =- 168 THEN
            sigmoid_f := 982;
        ELSIF x =- 167 THEN
            sigmoid_f := 982;
        ELSIF x =- 166 THEN
            sigmoid_f := 982;
        ELSIF x =- 165 THEN
            sigmoid_f := 982;
        ELSIF x =- 164 THEN
            sigmoid_f := 983;
        ELSIF x =- 163 THEN
            sigmoid_f := 983;
        ELSIF x =- 162 THEN
            sigmoid_f := 983;
        ELSIF x =- 161 THEN
            sigmoid_f := 983;
        ELSIF x =- 160 THEN
            sigmoid_f := 984;
        ELSIF x =- 159 THEN
            sigmoid_f := 984;
        ELSIF x =- 158 THEN
            sigmoid_f := 984;
        ELSIF x =- 157 THEN
            sigmoid_f := 984;
        ELSIF x =- 156 THEN
            sigmoid_f := 985;
        ELSIF x =- 155 THEN
            sigmoid_f := 985;
        ELSIF x =- 154 THEN
            sigmoid_f := 985;
        ELSIF x =- 153 THEN
            sigmoid_f := 985;
        ELSIF x =- 152 THEN
            sigmoid_f := 986;
        ELSIF x =- 151 THEN
            sigmoid_f := 986;
        ELSIF x =- 150 THEN
            sigmoid_f := 986;
        ELSIF x =- 149 THEN
            sigmoid_f := 986;
        ELSIF x =- 148 THEN
            sigmoid_f := 987;
        ELSIF x =- 147 THEN
            sigmoid_f := 987;
        ELSIF x =- 146 THEN
            sigmoid_f := 987;
        ELSIF x =- 145 THEN
            sigmoid_f := 987;
        ELSIF x =- 144 THEN
            sigmoid_f := 988;
        ELSIF x =- 143 THEN
            sigmoid_f := 988;
        ELSIF x =- 142 THEN
            sigmoid_f := 988;
        ELSIF x =- 141 THEN
            sigmoid_f := 988;
        ELSIF x =- 140 THEN
            sigmoid_f := 989;
        ELSIF x =- 139 THEN
            sigmoid_f := 989;
        ELSIF x =- 138 THEN
            sigmoid_f := 989;
        ELSIF x =- 137 THEN
            sigmoid_f := 989;
        ELSIF x =- 136 THEN
            sigmoid_f := 990;
        ELSIF x =- 135 THEN
            sigmoid_f := 990;
        ELSIF x =- 134 THEN
            sigmoid_f := 990;
        ELSIF x =- 133 THEN
            sigmoid_f := 990;
        ELSIF x =- 132 THEN
            sigmoid_f := 991;
        ELSIF x =- 131 THEN
            sigmoid_f := 991;
        ELSIF x =- 130 THEN
            sigmoid_f := 991;
        ELSIF x =- 129 THEN
            sigmoid_f := 991;
        ELSIF x =- 128 THEN
            sigmoid_f := 992;
        ELSIF x =- 127 THEN
            sigmoid_f := 992;
        ELSIF x =- 126 THEN
            sigmoid_f := 992;
        ELSIF x =- 125 THEN
            sigmoid_f := 992;
        ELSIF x =- 124 THEN
            sigmoid_f := 993;
        ELSIF x =- 123 THEN
            sigmoid_f := 993;
        ELSIF x =- 122 THEN
            sigmoid_f := 993;
        ELSIF x =- 121 THEN
            sigmoid_f := 993;
        ELSIF x =- 120 THEN
            sigmoid_f := 994;
        ELSIF x =- 119 THEN
            sigmoid_f := 994;
        ELSIF x =- 118 THEN
            sigmoid_f := 994;
        ELSIF x =- 117 THEN
            sigmoid_f := 994;
        ELSIF x =- 116 THEN
            sigmoid_f := 995;
        ELSIF x =- 115 THEN
            sigmoid_f := 995;
        ELSIF x =- 114 THEN
            sigmoid_f := 995;
        ELSIF x =- 113 THEN
            sigmoid_f := 995;
        ELSIF x =- 112 THEN
            sigmoid_f := 996;
        ELSIF x =- 111 THEN
            sigmoid_f := 996;
        ELSIF x =- 110 THEN
            sigmoid_f := 996;
        ELSIF x =- 109 THEN
            sigmoid_f := 996;
        ELSIF x =- 108 THEN
            sigmoid_f := 997;
        ELSIF x =- 107 THEN
            sigmoid_f := 997;
        ELSIF x =- 106 THEN
            sigmoid_f := 997;
        ELSIF x =- 105 THEN
            sigmoid_f := 997;
        ELSIF x =- 104 THEN
            sigmoid_f := 998;
        ELSIF x =- 103 THEN
            sigmoid_f := 998;
        ELSIF x =- 102 THEN
            sigmoid_f := 998;
        ELSIF x =- 101 THEN
            sigmoid_f := 998;
        ELSIF x =- 100 THEN
            sigmoid_f := 999;
        ELSIF x =- 99 THEN
            sigmoid_f := 999;
        ELSIF x =- 98 THEN
            sigmoid_f := 999;
        ELSIF x =- 97 THEN
            sigmoid_f := 999;
        ELSIF x =- 96 THEN
            sigmoid_f := 1000;
        ELSIF x =- 95 THEN
            sigmoid_f := 1000;
        ELSIF x =- 94 THEN
            sigmoid_f := 1000;
        ELSIF x =- 93 THEN
            sigmoid_f := 1000;
        ELSIF x =- 92 THEN
            sigmoid_f := 1001;
        ELSIF x =- 91 THEN
            sigmoid_f := 1001;
        ELSIF x =- 90 THEN
            sigmoid_f := 1001;
        ELSIF x =- 89 THEN
            sigmoid_f := 1001;
        ELSIF x =- 88 THEN
            sigmoid_f := 1002;
        ELSIF x =- 87 THEN
            sigmoid_f := 1002;
        ELSIF x =- 86 THEN
            sigmoid_f := 1002;
        ELSIF x =- 85 THEN
            sigmoid_f := 1002;
        ELSIF x =- 84 THEN
            sigmoid_f := 1003;
        ELSIF x =- 83 THEN
            sigmoid_f := 1003;
        ELSIF x =- 82 THEN
            sigmoid_f := 1003;
        ELSIF x =- 81 THEN
            sigmoid_f := 1003;
        ELSIF x =- 80 THEN
            sigmoid_f := 1004;
        ELSIF x =- 79 THEN
            sigmoid_f := 1004;
        ELSIF x =- 78 THEN
            sigmoid_f := 1004;
        ELSIF x =- 77 THEN
            sigmoid_f := 1004;
        ELSIF x =- 76 THEN
            sigmoid_f := 1005;
        ELSIF x =- 75 THEN
            sigmoid_f := 1005;
        ELSIF x =- 74 THEN
            sigmoid_f := 1005;
        ELSIF x =- 73 THEN
            sigmoid_f := 1005;
        ELSIF x =- 72 THEN
            sigmoid_f := 1006;
        ELSIF x =- 71 THEN
            sigmoid_f := 1006;
        ELSIF x =- 70 THEN
            sigmoid_f := 1006;
        ELSIF x =- 69 THEN
            sigmoid_f := 1006;
        ELSIF x =- 68 THEN
            sigmoid_f := 1007;
        ELSIF x =- 67 THEN
            sigmoid_f := 1007;
        ELSIF x =- 66 THEN
            sigmoid_f := 1007;
        ELSIF x =- 65 THEN
            sigmoid_f := 1007;
        ELSIF x =- 64 THEN
            sigmoid_f := 1008;
        ELSIF x =- 63 THEN
            sigmoid_f := 1008;
        ELSIF x =- 62 THEN
            sigmoid_f := 1008;
        ELSIF x =- 61 THEN
            sigmoid_f := 1008;
        ELSIF x =- 60 THEN
            sigmoid_f := 1009;
        ELSIF x =- 59 THEN
            sigmoid_f := 1009;
        ELSIF x =- 58 THEN
            sigmoid_f := 1009;
        ELSIF x =- 57 THEN
            sigmoid_f := 1009;
        ELSIF x =- 56 THEN
            sigmoid_f := 1010;
        ELSIF x =- 55 THEN
            sigmoid_f := 1010;
        ELSIF x =- 54 THEN
            sigmoid_f := 1010;
        ELSIF x =- 53 THEN
            sigmoid_f := 1010;
        ELSIF x =- 52 THEN
            sigmoid_f := 1011;
        ELSIF x =- 51 THEN
            sigmoid_f := 1011;
        ELSIF x =- 50 THEN
            sigmoid_f := 1011;
        ELSIF x =- 49 THEN
            sigmoid_f := 1011;
        ELSIF x =- 48 THEN
            sigmoid_f := 1012;
        ELSIF x =- 47 THEN
            sigmoid_f := 1012;
        ELSIF x =- 46 THEN
            sigmoid_f := 1012;
        ELSIF x =- 45 THEN
            sigmoid_f := 1012;
        ELSIF x =- 44 THEN
            sigmoid_f := 1013;
        ELSIF x =- 43 THEN
            sigmoid_f := 1013;
        ELSIF x =- 42 THEN
            sigmoid_f := 1013;
        ELSIF x =- 41 THEN
            sigmoid_f := 1013;
        ELSIF x =- 40 THEN
            sigmoid_f := 1014;
        ELSIF x =- 39 THEN
            sigmoid_f := 1014;
        ELSIF x =- 38 THEN
            sigmoid_f := 1014;
        ELSIF x =- 37 THEN
            sigmoid_f := 1014;
        ELSIF x =- 36 THEN
            sigmoid_f := 1015;
        ELSIF x =- 35 THEN
            sigmoid_f := 1015;
        ELSIF x =- 34 THEN
            sigmoid_f := 1015;
        ELSIF x =- 33 THEN
            sigmoid_f := 1015;
        ELSIF x =- 32 THEN
            sigmoid_f := 1016;
        ELSIF x =- 31 THEN
            sigmoid_f := 1016;
        ELSIF x =- 30 THEN
            sigmoid_f := 1016;
        ELSIF x =- 29 THEN
            sigmoid_f := 1016;
        ELSIF x =- 28 THEN
            sigmoid_f := 1017;
        ELSIF x =- 27 THEN
            sigmoid_f := 1017;
        ELSIF x =- 26 THEN
            sigmoid_f := 1017;
        ELSIF x =- 25 THEN
            sigmoid_f := 1017;
        ELSIF x =- 24 THEN
            sigmoid_f := 1018;
        ELSIF x =- 23 THEN
            sigmoid_f := 1018;
        ELSIF x =- 22 THEN
            sigmoid_f := 1018;
        ELSIF x =- 21 THEN
            sigmoid_f := 1018;
        ELSIF x =- 20 THEN
            sigmoid_f := 1019;
        ELSIF x =- 19 THEN
            sigmoid_f := 1019;
        ELSIF x =- 18 THEN
            sigmoid_f := 1019;
        ELSIF x =- 17 THEN
            sigmoid_f := 1019;
        ELSIF x =- 16 THEN
            sigmoid_f := 1020;
        ELSIF x =- 15 THEN
            sigmoid_f := 1020;
        ELSIF x =- 14 THEN
            sigmoid_f := 1020;
        ELSIF x =- 13 THEN
            sigmoid_f := 1020;
        ELSIF x =- 12 THEN
            sigmoid_f := 1021;
        ELSIF x =- 11 THEN
            sigmoid_f := 1021;
        ELSIF x =- 10 THEN
            sigmoid_f := 1021;
        ELSIF x =- 9 THEN
            sigmoid_f := 1021;
        ELSIF x =- 8 THEN
            sigmoid_f := 1022;
        ELSIF x =- 7 THEN
            sigmoid_f := 1022;
        ELSIF x =- 6 THEN
            sigmoid_f := 1022;
        ELSIF x =- 5 THEN
            sigmoid_f := 1022;
        ELSIF x =- 4 THEN
            sigmoid_f := 1023;
        ELSIF x =- 3 THEN
            sigmoid_f := 1023;
        ELSIF x =- 2 THEN
            sigmoid_f := 1023;
        ELSIF x =- 1 THEN
            sigmoid_f := 1023;
        ELSIF x = 0 THEN
            sigmoid_f := 1024;
        ELSIF x = 1 THEN
            sigmoid_f := 1024;
        ELSIF x = 2 THEN
            sigmoid_f := 1024;
        ELSIF x = 3 THEN
            sigmoid_f := 1024;
        ELSIF x = 4 THEN
            sigmoid_f := 1025;
        ELSIF x = 5 THEN
            sigmoid_f := 1025;
        ELSIF x = 6 THEN
            sigmoid_f := 1025;
        ELSIF x = 7 THEN
            sigmoid_f := 1025;
        ELSIF x = 8 THEN
            sigmoid_f := 1026;
        ELSIF x = 9 THEN
            sigmoid_f := 1026;
        ELSIF x = 10 THEN
            sigmoid_f := 1026;
        ELSIF x = 11 THEN
            sigmoid_f := 1026;
        ELSIF x = 12 THEN
            sigmoid_f := 1027;
        ELSIF x = 13 THEN
            sigmoid_f := 1027;
        ELSIF x = 14 THEN
            sigmoid_f := 1027;
        ELSIF x = 15 THEN
            sigmoid_f := 1027;
        ELSIF x = 16 THEN
            sigmoid_f := 1028;
        ELSIF x = 17 THEN
            sigmoid_f := 1028;
        ELSIF x = 18 THEN
            sigmoid_f := 1028;
        ELSIF x = 19 THEN
            sigmoid_f := 1028;
        ELSIF x = 20 THEN
            sigmoid_f := 1029;
        ELSIF x = 21 THEN
            sigmoid_f := 1029;
        ELSIF x = 22 THEN
            sigmoid_f := 1029;
        ELSIF x = 23 THEN
            sigmoid_f := 1029;
        ELSIF x = 24 THEN
            sigmoid_f := 1030;
        ELSIF x = 25 THEN
            sigmoid_f := 1030;
        ELSIF x = 26 THEN
            sigmoid_f := 1030;
        ELSIF x = 27 THEN
            sigmoid_f := 1030;
        ELSIF x = 28 THEN
            sigmoid_f := 1031;
        ELSIF x = 29 THEN
            sigmoid_f := 1031;
        ELSIF x = 30 THEN
            sigmoid_f := 1031;
        ELSIF x = 31 THEN
            sigmoid_f := 1031;
        ELSIF x = 32 THEN
            sigmoid_f := 1032;
        ELSIF x = 33 THEN
            sigmoid_f := 1032;
        ELSIF x = 34 THEN
            sigmoid_f := 1032;
        ELSIF x = 35 THEN
            sigmoid_f := 1032;
        ELSIF x = 36 THEN
            sigmoid_f := 1033;
        ELSIF x = 37 THEN
            sigmoid_f := 1033;
        ELSIF x = 38 THEN
            sigmoid_f := 1033;
        ELSIF x = 39 THEN
            sigmoid_f := 1033;
        ELSIF x = 40 THEN
            sigmoid_f := 1034;
        ELSIF x = 41 THEN
            sigmoid_f := 1034;
        ELSIF x = 42 THEN
            sigmoid_f := 1034;
        ELSIF x = 43 THEN
            sigmoid_f := 1034;
        ELSIF x = 44 THEN
            sigmoid_f := 1035;
        ELSIF x = 45 THEN
            sigmoid_f := 1035;
        ELSIF x = 46 THEN
            sigmoid_f := 1035;
        ELSIF x = 47 THEN
            sigmoid_f := 1035;
        ELSIF x = 48 THEN
            sigmoid_f := 1036;
        ELSIF x = 49 THEN
            sigmoid_f := 1036;
        ELSIF x = 50 THEN
            sigmoid_f := 1036;
        ELSIF x = 51 THEN
            sigmoid_f := 1036;
        ELSIF x = 52 THEN
            sigmoid_f := 1037;
        ELSIF x = 53 THEN
            sigmoid_f := 1037;
        ELSIF x = 54 THEN
            sigmoid_f := 1037;
        ELSIF x = 55 THEN
            sigmoid_f := 1037;
        ELSIF x = 56 THEN
            sigmoid_f := 1038;
        ELSIF x = 57 THEN
            sigmoid_f := 1038;
        ELSIF x = 58 THEN
            sigmoid_f := 1038;
        ELSIF x = 59 THEN
            sigmoid_f := 1038;
        ELSIF x = 60 THEN
            sigmoid_f := 1039;
        ELSIF x = 61 THEN
            sigmoid_f := 1039;
        ELSIF x = 62 THEN
            sigmoid_f := 1039;
        ELSIF x = 63 THEN
            sigmoid_f := 1039;
        ELSIF x = 64 THEN
            sigmoid_f := 1040;
        ELSIF x = 65 THEN
            sigmoid_f := 1040;
        ELSIF x = 66 THEN
            sigmoid_f := 1040;
        ELSIF x = 67 THEN
            sigmoid_f := 1040;
        ELSIF x = 68 THEN
            sigmoid_f := 1041;
        ELSIF x = 69 THEN
            sigmoid_f := 1041;
        ELSIF x = 70 THEN
            sigmoid_f := 1041;
        ELSIF x = 71 THEN
            sigmoid_f := 1041;
        ELSIF x = 72 THEN
            sigmoid_f := 1042;
        ELSIF x = 73 THEN
            sigmoid_f := 1042;
        ELSIF x = 74 THEN
            sigmoid_f := 1042;
        ELSIF x = 75 THEN
            sigmoid_f := 1042;
        ELSIF x = 76 THEN
            sigmoid_f := 1043;
        ELSIF x = 77 THEN
            sigmoid_f := 1043;
        ELSIF x = 78 THEN
            sigmoid_f := 1043;
        ELSIF x = 79 THEN
            sigmoid_f := 1043;
        ELSIF x = 80 THEN
            sigmoid_f := 1044;
        ELSIF x = 81 THEN
            sigmoid_f := 1044;
        ELSIF x = 82 THEN
            sigmoid_f := 1044;
        ELSIF x = 83 THEN
            sigmoid_f := 1044;
        ELSIF x = 84 THEN
            sigmoid_f := 1045;
        ELSIF x = 85 THEN
            sigmoid_f := 1045;
        ELSIF x = 86 THEN
            sigmoid_f := 1045;
        ELSIF x = 87 THEN
            sigmoid_f := 1045;
        ELSIF x = 88 THEN
            sigmoid_f := 1046;
        ELSIF x = 89 THEN
            sigmoid_f := 1046;
        ELSIF x = 90 THEN
            sigmoid_f := 1046;
        ELSIF x = 91 THEN
            sigmoid_f := 1046;
        ELSIF x = 92 THEN
            sigmoid_f := 1047;
        ELSIF x = 93 THEN
            sigmoid_f := 1047;
        ELSIF x = 94 THEN
            sigmoid_f := 1047;
        ELSIF x = 95 THEN
            sigmoid_f := 1047;
        ELSIF x = 96 THEN
            sigmoid_f := 1048;
        ELSIF x = 97 THEN
            sigmoid_f := 1048;
        ELSIF x = 98 THEN
            sigmoid_f := 1048;
        ELSIF x = 99 THEN
            sigmoid_f := 1048;
        ELSIF x = 100 THEN
            sigmoid_f := 1049;
        ELSIF x = 101 THEN
            sigmoid_f := 1049;
        ELSIF x = 102 THEN
            sigmoid_f := 1049;
        ELSIF x = 103 THEN
            sigmoid_f := 1049;
        ELSIF x = 104 THEN
            sigmoid_f := 1050;
        ELSIF x = 105 THEN
            sigmoid_f := 1050;
        ELSIF x = 106 THEN
            sigmoid_f := 1050;
        ELSIF x = 107 THEN
            sigmoid_f := 1050;
        ELSIF x = 108 THEN
            sigmoid_f := 1051;
        ELSIF x = 109 THEN
            sigmoid_f := 1051;
        ELSIF x = 110 THEN
            sigmoid_f := 1051;
        ELSIF x = 111 THEN
            sigmoid_f := 1051;
        ELSIF x = 112 THEN
            sigmoid_f := 1052;
        ELSIF x = 113 THEN
            sigmoid_f := 1052;
        ELSIF x = 114 THEN
            sigmoid_f := 1052;
        ELSIF x = 115 THEN
            sigmoid_f := 1052;
        ELSIF x = 116 THEN
            sigmoid_f := 1053;
        ELSIF x = 117 THEN
            sigmoid_f := 1053;
        ELSIF x = 118 THEN
            sigmoid_f := 1053;
        ELSIF x = 119 THEN
            sigmoid_f := 1053;
        ELSIF x = 120 THEN
            sigmoid_f := 1054;
        ELSIF x = 121 THEN
            sigmoid_f := 1054;
        ELSIF x = 122 THEN
            sigmoid_f := 1054;
        ELSIF x = 123 THEN
            sigmoid_f := 1054;
        ELSIF x = 124 THEN
            sigmoid_f := 1055;
        ELSIF x = 125 THEN
            sigmoid_f := 1055;
        ELSIF x = 126 THEN
            sigmoid_f := 1055;
        ELSIF x = 127 THEN
            sigmoid_f := 1055;
        ELSIF x = 128 THEN
            sigmoid_f := 1056;
        ELSIF x = 129 THEN
            sigmoid_f := 1056;
        ELSIF x = 130 THEN
            sigmoid_f := 1056;
        ELSIF x = 131 THEN
            sigmoid_f := 1056;
        ELSIF x = 132 THEN
            sigmoid_f := 1057;
        ELSIF x = 133 THEN
            sigmoid_f := 1057;
        ELSIF x = 134 THEN
            sigmoid_f := 1057;
        ELSIF x = 135 THEN
            sigmoid_f := 1057;
        ELSIF x = 136 THEN
            sigmoid_f := 1058;
        ELSIF x = 137 THEN
            sigmoid_f := 1058;
        ELSIF x = 138 THEN
            sigmoid_f := 1058;
        ELSIF x = 139 THEN
            sigmoid_f := 1058;
        ELSIF x = 140 THEN
            sigmoid_f := 1059;
        ELSIF x = 141 THEN
            sigmoid_f := 1059;
        ELSIF x = 142 THEN
            sigmoid_f := 1059;
        ELSIF x = 143 THEN
            sigmoid_f := 1059;
        ELSIF x = 144 THEN
            sigmoid_f := 1060;
        ELSIF x = 145 THEN
            sigmoid_f := 1060;
        ELSIF x = 146 THEN
            sigmoid_f := 1060;
        ELSIF x = 147 THEN
            sigmoid_f := 1060;
        ELSIF x = 148 THEN
            sigmoid_f := 1061;
        ELSIF x = 149 THEN
            sigmoid_f := 1061;
        ELSIF x = 150 THEN
            sigmoid_f := 1061;
        ELSIF x = 151 THEN
            sigmoid_f := 1061;
        ELSIF x = 152 THEN
            sigmoid_f := 1062;
        ELSIF x = 153 THEN
            sigmoid_f := 1062;
        ELSIF x = 154 THEN
            sigmoid_f := 1062;
        ELSIF x = 155 THEN
            sigmoid_f := 1062;
        ELSIF x = 156 THEN
            sigmoid_f := 1063;
        ELSIF x = 157 THEN
            sigmoid_f := 1063;
        ELSIF x = 158 THEN
            sigmoid_f := 1063;
        ELSIF x = 159 THEN
            sigmoid_f := 1063;
        ELSIF x = 160 THEN
            sigmoid_f := 1064;
        ELSIF x = 161 THEN
            sigmoid_f := 1064;
        ELSIF x = 162 THEN
            sigmoid_f := 1064;
        ELSIF x = 163 THEN
            sigmoid_f := 1064;
        ELSIF x = 164 THEN
            sigmoid_f := 1065;
        ELSIF x = 165 THEN
            sigmoid_f := 1065;
        ELSIF x = 166 THEN
            sigmoid_f := 1065;
        ELSIF x = 167 THEN
            sigmoid_f := 1065;
        ELSIF x = 168 THEN
            sigmoid_f := 1066;
        ELSIF x = 169 THEN
            sigmoid_f := 1066;
        ELSIF x = 170 THEN
            sigmoid_f := 1066;
        ELSIF x = 171 THEN
            sigmoid_f := 1066;
        ELSIF x = 172 THEN
            sigmoid_f := 1067;
        ELSIF x = 173 THEN
            sigmoid_f := 1067;
        ELSIF x = 174 THEN
            sigmoid_f := 1067;
        ELSIF x = 175 THEN
            sigmoid_f := 1067;
        ELSIF x = 176 THEN
            sigmoid_f := 1068;
        ELSIF x = 177 THEN
            sigmoid_f := 1068;
        ELSIF x = 178 THEN
            sigmoid_f := 1068;
        ELSIF x = 179 THEN
            sigmoid_f := 1068;
        ELSIF x = 180 THEN
            sigmoid_f := 1069;
        ELSIF x = 181 THEN
            sigmoid_f := 1069;
        ELSIF x = 182 THEN
            sigmoid_f := 1069;
        ELSIF x = 183 THEN
            sigmoid_f := 1069;
        ELSIF x = 184 THEN
            sigmoid_f := 1070;
        ELSIF x = 185 THEN
            sigmoid_f := 1070;
        ELSIF x = 186 THEN
            sigmoid_f := 1070;
        ELSIF x = 187 THEN
            sigmoid_f := 1070;
        ELSIF x = 188 THEN
            sigmoid_f := 1071;
        ELSIF x = 189 THEN
            sigmoid_f := 1071;
        ELSIF x = 190 THEN
            sigmoid_f := 1071;
        ELSIF x = 191 THEN
            sigmoid_f := 1071;
        ELSIF x = 192 THEN
            sigmoid_f := 1072;
        ELSIF x = 193 THEN
            sigmoid_f := 1072;
        ELSIF x = 194 THEN
            sigmoid_f := 1072;
        ELSIF x = 195 THEN
            sigmoid_f := 1072;
        ELSIF x = 196 THEN
            sigmoid_f := 1073;
        ELSIF x = 197 THEN
            sigmoid_f := 1073;
        ELSIF x = 198 THEN
            sigmoid_f := 1073;
        ELSIF x = 199 THEN
            sigmoid_f := 1073;
        ELSIF x = 200 THEN
            sigmoid_f := 1074;
        ELSIF x = 201 THEN
            sigmoid_f := 1074;
        ELSIF x = 202 THEN
            sigmoid_f := 1074;
        ELSIF x = 203 THEN
            sigmoid_f := 1074;
        ELSIF x = 204 THEN
            sigmoid_f := 1075;
        ELSIF x = 205 THEN
            sigmoid_f := 1075;
        ELSIF x = 206 THEN
            sigmoid_f := 1075;
        ELSIF x = 207 THEN
            sigmoid_f := 1075;
        ELSIF x = 208 THEN
            sigmoid_f := 1076;
        ELSIF x = 209 THEN
            sigmoid_f := 1076;
        ELSIF x = 210 THEN
            sigmoid_f := 1076;
        ELSIF x = 211 THEN
            sigmoid_f := 1076;
        ELSIF x = 212 THEN
            sigmoid_f := 1077;
        ELSIF x = 213 THEN
            sigmoid_f := 1077;
        ELSIF x = 214 THEN
            sigmoid_f := 1077;
        ELSIF x = 215 THEN
            sigmoid_f := 1077;
        ELSIF x = 216 THEN
            sigmoid_f := 1078;
        ELSIF x = 217 THEN
            sigmoid_f := 1078;
        ELSIF x = 218 THEN
            sigmoid_f := 1078;
        ELSIF x = 219 THEN
            sigmoid_f := 1078;
        ELSIF x = 220 THEN
            sigmoid_f := 1079;
        ELSIF x = 221 THEN
            sigmoid_f := 1079;
        ELSIF x = 222 THEN
            sigmoid_f := 1079;
        ELSIF x = 223 THEN
            sigmoid_f := 1079;
        ELSIF x = 224 THEN
            sigmoid_f := 1080;
        ELSIF x = 225 THEN
            sigmoid_f := 1080;
        ELSIF x = 226 THEN
            sigmoid_f := 1080;
        ELSIF x = 227 THEN
            sigmoid_f := 1080;
        ELSIF x = 228 THEN
            sigmoid_f := 1081;
        ELSIF x = 229 THEN
            sigmoid_f := 1081;
        ELSIF x = 230 THEN
            sigmoid_f := 1081;
        ELSIF x = 231 THEN
            sigmoid_f := 1081;
        ELSIF x = 232 THEN
            sigmoid_f := 1082;
        ELSIF x = 233 THEN
            sigmoid_f := 1082;
        ELSIF x = 234 THEN
            sigmoid_f := 1082;
        ELSIF x = 235 THEN
            sigmoid_f := 1082;
        ELSIF x = 236 THEN
            sigmoid_f := 1083;
        ELSIF x = 237 THEN
            sigmoid_f := 1083;
        ELSIF x = 238 THEN
            sigmoid_f := 1083;
        ELSIF x = 239 THEN
            sigmoid_f := 1083;
        ELSIF x = 240 THEN
            sigmoid_f := 1084;
        ELSIF x = 241 THEN
            sigmoid_f := 1084;
        ELSIF x = 242 THEN
            sigmoid_f := 1084;
        ELSIF x = 243 THEN
            sigmoid_f := 1084;
        ELSIF x = 244 THEN
            sigmoid_f := 1085;
        ELSIF x = 245 THEN
            sigmoid_f := 1085;
        ELSIF x = 246 THEN
            sigmoid_f := 1085;
        ELSIF x = 247 THEN
            sigmoid_f := 1085;
        ELSIF x = 248 THEN
            sigmoid_f := 1086;
        ELSIF x = 249 THEN
            sigmoid_f := 1086;
        ELSIF x = 250 THEN
            sigmoid_f := 1086;
        ELSIF x = 251 THEN
            sigmoid_f := 1086;
        ELSIF x = 252 THEN
            sigmoid_f := 1087;
        ELSIF x = 253 THEN
            sigmoid_f := 1087;
        ELSIF x = 254 THEN
            sigmoid_f := 1087;
        ELSIF x = 255 THEN
            sigmoid_f := 1087;
        ELSIF x = 256 THEN
            sigmoid_f := 1088;
        ELSIF x = 257 THEN
            sigmoid_f := 1088;
        ELSIF x = 258 THEN
            sigmoid_f := 1088;
        ELSIF x = 259 THEN
            sigmoid_f := 1088;
        ELSIF x = 260 THEN
            sigmoid_f := 1089;
        ELSIF x = 261 THEN
            sigmoid_f := 1089;
        ELSIF x = 262 THEN
            sigmoid_f := 1089;
        ELSIF x = 263 THEN
            sigmoid_f := 1089;
        ELSIF x = 264 THEN
            sigmoid_f := 1090;
        ELSIF x = 265 THEN
            sigmoid_f := 1090;
        ELSIF x = 266 THEN
            sigmoid_f := 1090;
        ELSIF x = 267 THEN
            sigmoid_f := 1090;
        ELSIF x = 268 THEN
            sigmoid_f := 1091;
        ELSIF x = 269 THEN
            sigmoid_f := 1091;
        ELSIF x = 270 THEN
            sigmoid_f := 1091;
        ELSIF x = 271 THEN
            sigmoid_f := 1091;
        ELSIF x = 272 THEN
            sigmoid_f := 1092;
        ELSIF x = 273 THEN
            sigmoid_f := 1092;
        ELSIF x = 274 THEN
            sigmoid_f := 1092;
        ELSIF x = 275 THEN
            sigmoid_f := 1092;
        ELSIF x = 276 THEN
            sigmoid_f := 1093;
        ELSIF x = 277 THEN
            sigmoid_f := 1093;
        ELSIF x = 278 THEN
            sigmoid_f := 1093;
        ELSIF x = 279 THEN
            sigmoid_f := 1093;
        ELSIF x = 280 THEN
            sigmoid_f := 1094;
        ELSIF x = 281 THEN
            sigmoid_f := 1094;
        ELSIF x = 282 THEN
            sigmoid_f := 1094;
        ELSIF x = 283 THEN
            sigmoid_f := 1094;
        ELSIF x = 284 THEN
            sigmoid_f := 1095;
        ELSIF x = 285 THEN
            sigmoid_f := 1095;
        ELSIF x = 286 THEN
            sigmoid_f := 1095;
        ELSIF x = 287 THEN
            sigmoid_f := 1095;
        ELSIF x = 288 THEN
            sigmoid_f := 1096;
        ELSIF x = 289 THEN
            sigmoid_f := 1096;
        ELSIF x = 290 THEN
            sigmoid_f := 1096;
        ELSIF x = 291 THEN
            sigmoid_f := 1096;
        ELSIF x = 292 THEN
            sigmoid_f := 1097;
        ELSIF x = 293 THEN
            sigmoid_f := 1097;
        ELSIF x = 294 THEN
            sigmoid_f := 1097;
        ELSIF x = 295 THEN
            sigmoid_f := 1097;
        ELSIF x = 296 THEN
            sigmoid_f := 1098;
        ELSIF x = 297 THEN
            sigmoid_f := 1098;
        ELSIF x = 298 THEN
            sigmoid_f := 1098;
        ELSIF x = 299 THEN
            sigmoid_f := 1098;
        ELSIF x = 300 THEN
            sigmoid_f := 1099;
        ELSIF x = 301 THEN
            sigmoid_f := 1099;
        ELSIF x = 302 THEN
            sigmoid_f := 1099;
        ELSIF x = 303 THEN
            sigmoid_f := 1099;
        ELSIF x = 304 THEN
            sigmoid_f := 1100;
        ELSIF x = 305 THEN
            sigmoid_f := 1100;
        ELSIF x = 306 THEN
            sigmoid_f := 1100;
        ELSIF x = 307 THEN
            sigmoid_f := 1100;
        ELSIF x = 308 THEN
            sigmoid_f := 1101;
        ELSIF x = 309 THEN
            sigmoid_f := 1101;
        ELSIF x = 310 THEN
            sigmoid_f := 1101;
        ELSIF x = 311 THEN
            sigmoid_f := 1101;
        ELSIF x = 312 THEN
            sigmoid_f := 1102;
        ELSIF x = 313 THEN
            sigmoid_f := 1102;
        ELSIF x = 314 THEN
            sigmoid_f := 1102;
        ELSIF x = 315 THEN
            sigmoid_f := 1102;
        ELSIF x = 316 THEN
            sigmoid_f := 1103;
        ELSIF x = 317 THEN
            sigmoid_f := 1103;
        ELSIF x = 318 THEN
            sigmoid_f := 1103;
        ELSIF x = 319 THEN
            sigmoid_f := 1103;
        ELSIF x = 320 THEN
            sigmoid_f := 1104;
        ELSIF x = 321 THEN
            sigmoid_f := 1104;
        ELSIF x = 322 THEN
            sigmoid_f := 1104;
        ELSIF x = 323 THEN
            sigmoid_f := 1104;
        ELSIF x = 324 THEN
            sigmoid_f := 1105;
        ELSIF x = 325 THEN
            sigmoid_f := 1105;
        ELSIF x = 326 THEN
            sigmoid_f := 1105;
        ELSIF x = 327 THEN
            sigmoid_f := 1105;
        ELSIF x = 328 THEN
            sigmoid_f := 1106;
        ELSIF x = 329 THEN
            sigmoid_f := 1106;
        ELSIF x = 330 THEN
            sigmoid_f := 1106;
        ELSIF x = 331 THEN
            sigmoid_f := 1106;
        ELSIF x = 332 THEN
            sigmoid_f := 1107;
        ELSIF x = 333 THEN
            sigmoid_f := 1107;
        ELSIF x = 334 THEN
            sigmoid_f := 1107;
        ELSIF x = 335 THEN
            sigmoid_f := 1107;
        ELSIF x = 336 THEN
            sigmoid_f := 1108;
        ELSIF x = 337 THEN
            sigmoid_f := 1108;
        ELSIF x = 338 THEN
            sigmoid_f := 1108;
        ELSIF x = 339 THEN
            sigmoid_f := 1108;
        ELSIF x = 340 THEN
            sigmoid_f := 1109;
        ELSIF x = 341 THEN
            sigmoid_f := 1109;
        ELSIF x = 342 THEN
            sigmoid_f := 1109;
        ELSIF x = 343 THEN
            sigmoid_f := 1109;
        ELSIF x = 344 THEN
            sigmoid_f := 1110;
        ELSIF x = 345 THEN
            sigmoid_f := 1110;
        ELSIF x = 346 THEN
            sigmoid_f := 1110;
        ELSIF x = 347 THEN
            sigmoid_f := 1110;
        ELSIF x = 348 THEN
            sigmoid_f := 1111;
        ELSIF x = 349 THEN
            sigmoid_f := 1111;
        ELSIF x = 350 THEN
            sigmoid_f := 1111;
        ELSIF x = 351 THEN
            sigmoid_f := 1111;
        ELSIF x = 352 THEN
            sigmoid_f := 1112;
        ELSIF x = 353 THEN
            sigmoid_f := 1112;
        ELSIF x = 354 THEN
            sigmoid_f := 1112;
        ELSIF x = 355 THEN
            sigmoid_f := 1112;
        ELSIF x = 356 THEN
            sigmoid_f := 1113;
        ELSIF x = 357 THEN
            sigmoid_f := 1113;
        ELSIF x = 358 THEN
            sigmoid_f := 1113;
        ELSIF x = 359 THEN
            sigmoid_f := 1113;
        ELSIF x = 360 THEN
            sigmoid_f := 1114;
        ELSIF x = 361 THEN
            sigmoid_f := 1114;
        ELSIF x = 362 THEN
            sigmoid_f := 1114;
        ELSIF x = 363 THEN
            sigmoid_f := 1114;
        ELSIF x = 364 THEN
            sigmoid_f := 1115;
        ELSIF x = 365 THEN
            sigmoid_f := 1115;
        ELSIF x = 366 THEN
            sigmoid_f := 1115;
        ELSIF x = 367 THEN
            sigmoid_f := 1115;
        ELSIF x = 368 THEN
            sigmoid_f := 1116;
        ELSIF x = 369 THEN
            sigmoid_f := 1116;
        ELSIF x = 370 THEN
            sigmoid_f := 1116;
        ELSIF x = 371 THEN
            sigmoid_f := 1116;
        ELSIF x = 372 THEN
            sigmoid_f := 1117;
        ELSIF x = 373 THEN
            sigmoid_f := 1117;
        ELSIF x = 374 THEN
            sigmoid_f := 1117;
        ELSIF x = 375 THEN
            sigmoid_f := 1117;
        ELSIF x = 376 THEN
            sigmoid_f := 1118;
        ELSIF x = 377 THEN
            sigmoid_f := 1118;
        ELSIF x = 378 THEN
            sigmoid_f := 1118;
        ELSIF x = 379 THEN
            sigmoid_f := 1118;
        ELSIF x = 380 THEN
            sigmoid_f := 1119;
        ELSIF x = 381 THEN
            sigmoid_f := 1119;
        ELSIF x = 382 THEN
            sigmoid_f := 1119;
        ELSIF x = 383 THEN
            sigmoid_f := 1119;
        ELSIF x = 384 THEN
            sigmoid_f := 1120;
        ELSIF x = 385 THEN
            sigmoid_f := 1120;
        ELSIF x = 386 THEN
            sigmoid_f := 1120;
        ELSIF x = 387 THEN
            sigmoid_f := 1120;
        ELSIF x = 388 THEN
            sigmoid_f := 1121;
        ELSIF x = 389 THEN
            sigmoid_f := 1121;
        ELSIF x = 390 THEN
            sigmoid_f := 1121;
        ELSIF x = 391 THEN
            sigmoid_f := 1121;
        ELSIF x = 392 THEN
            sigmoid_f := 1122;
        ELSIF x = 393 THEN
            sigmoid_f := 1122;
        ELSIF x = 394 THEN
            sigmoid_f := 1122;
        ELSIF x = 395 THEN
            sigmoid_f := 1122;
        ELSIF x = 396 THEN
            sigmoid_f := 1123;
        ELSIF x = 397 THEN
            sigmoid_f := 1123;
        ELSIF x = 398 THEN
            sigmoid_f := 1123;
        ELSIF x = 399 THEN
            sigmoid_f := 1123;
        ELSIF x = 400 THEN
            sigmoid_f := 1124;
        ELSIF x = 401 THEN
            sigmoid_f := 1124;
        ELSIF x = 402 THEN
            sigmoid_f := 1124;
        ELSIF x = 403 THEN
            sigmoid_f := 1124;
        ELSIF x = 404 THEN
            sigmoid_f := 1125;
        ELSIF x = 405 THEN
            sigmoid_f := 1125;
        ELSIF x = 406 THEN
            sigmoid_f := 1125;
        ELSIF x = 407 THEN
            sigmoid_f := 1125;
        ELSIF x = 408 THEN
            sigmoid_f := 1126;
        ELSIF x = 409 THEN
            sigmoid_f := 1126;
        ELSIF x = 410 THEN
            sigmoid_f := 1126;
        ELSIF x = 411 THEN
            sigmoid_f := 1126;
        ELSIF x = 412 THEN
            sigmoid_f := 1127;
        ELSIF x = 413 THEN
            sigmoid_f := 1127;
        ELSIF x = 414 THEN
            sigmoid_f := 1127;
        ELSIF x = 415 THEN
            sigmoid_f := 1127;
        ELSIF x = 416 THEN
            sigmoid_f := 1128;
        ELSIF x = 417 THEN
            sigmoid_f := 1128;
        ELSIF x = 418 THEN
            sigmoid_f := 1128;
        ELSIF x = 419 THEN
            sigmoid_f := 1128;
        ELSIF x = 420 THEN
            sigmoid_f := 1129;
        ELSIF x = 421 THEN
            sigmoid_f := 1129;
        ELSIF x = 422 THEN
            sigmoid_f := 1129;
        ELSIF x = 423 THEN
            sigmoid_f := 1129;
        ELSIF x = 424 THEN
            sigmoid_f := 1130;
        ELSIF x = 425 THEN
            sigmoid_f := 1130;
        ELSIF x = 426 THEN
            sigmoid_f := 1130;
        ELSIF x = 427 THEN
            sigmoid_f := 1130;
        ELSIF x = 428 THEN
            sigmoid_f := 1131;
        ELSIF x = 429 THEN
            sigmoid_f := 1131;
        ELSIF x = 430 THEN
            sigmoid_f := 1131;
        ELSIF x = 431 THEN
            sigmoid_f := 1131;
        ELSIF x = 432 THEN
            sigmoid_f := 1132;
        ELSIF x = 433 THEN
            sigmoid_f := 1132;
        ELSIF x = 434 THEN
            sigmoid_f := 1132;
        ELSIF x = 435 THEN
            sigmoid_f := 1132;
        ELSIF x = 436 THEN
            sigmoid_f := 1133;
        ELSIF x = 437 THEN
            sigmoid_f := 1133;
        ELSIF x = 438 THEN
            sigmoid_f := 1133;
        ELSIF x = 439 THEN
            sigmoid_f := 1133;
        ELSIF x = 440 THEN
            sigmoid_f := 1134;
        ELSIF x = 441 THEN
            sigmoid_f := 1134;
        ELSIF x = 442 THEN
            sigmoid_f := 1134;
        ELSIF x = 443 THEN
            sigmoid_f := 1134;
        ELSIF x = 444 THEN
            sigmoid_f := 1135;
        ELSIF x = 445 THEN
            sigmoid_f := 1135;
        ELSIF x = 446 THEN
            sigmoid_f := 1135;
        ELSIF x = 447 THEN
            sigmoid_f := 1135;
        ELSIF x = 448 THEN
            sigmoid_f := 1136;
        ELSIF x = 449 THEN
            sigmoid_f := 1136;
        ELSIF x = 450 THEN
            sigmoid_f := 1136;
        ELSIF x = 451 THEN
            sigmoid_f := 1136;
        ELSIF x = 452 THEN
            sigmoid_f := 1137;
        ELSIF x = 453 THEN
            sigmoid_f := 1137;
        ELSIF x = 454 THEN
            sigmoid_f := 1137;
        ELSIF x = 455 THEN
            sigmoid_f := 1137;
        ELSIF x = 456 THEN
            sigmoid_f := 1138;
        ELSIF x = 457 THEN
            sigmoid_f := 1138;
        ELSIF x = 458 THEN
            sigmoid_f := 1138;
        ELSIF x = 459 THEN
            sigmoid_f := 1138;
        ELSIF x = 460 THEN
            sigmoid_f := 1139;
        ELSIF x = 461 THEN
            sigmoid_f := 1139;
        ELSIF x = 462 THEN
            sigmoid_f := 1139;
        ELSIF x = 463 THEN
            sigmoid_f := 1139;
        ELSIF x = 464 THEN
            sigmoid_f := 1140;
        ELSIF x = 465 THEN
            sigmoid_f := 1140;
        ELSIF x = 466 THEN
            sigmoid_f := 1140;
        ELSIF x = 467 THEN
            sigmoid_f := 1140;
        ELSIF x = 468 THEN
            sigmoid_f := 1141;
        ELSIF x = 469 THEN
            sigmoid_f := 1141;
        ELSIF x = 470 THEN
            sigmoid_f := 1141;
        ELSIF x = 471 THEN
            sigmoid_f := 1141;
        ELSIF x = 472 THEN
            sigmoid_f := 1142;
        ELSIF x = 473 THEN
            sigmoid_f := 1142;
        ELSIF x = 474 THEN
            sigmoid_f := 1142;
        ELSIF x = 475 THEN
            sigmoid_f := 1142;
        ELSIF x = 476 THEN
            sigmoid_f := 1143;
        ELSIF x = 477 THEN
            sigmoid_f := 1143;
        ELSIF x = 478 THEN
            sigmoid_f := 1143;
        ELSIF x = 479 THEN
            sigmoid_f := 1143;
        ELSIF x = 480 THEN
            sigmoid_f := 1144;
        ELSIF x = 481 THEN
            sigmoid_f := 1144;
        ELSIF x = 482 THEN
            sigmoid_f := 1144;
        ELSIF x = 483 THEN
            sigmoid_f := 1144;
        ELSIF x = 484 THEN
            sigmoid_f := 1145;
        ELSIF x = 485 THEN
            sigmoid_f := 1145;
        ELSIF x = 486 THEN
            sigmoid_f := 1145;
        ELSIF x = 487 THEN
            sigmoid_f := 1145;
        ELSIF x = 488 THEN
            sigmoid_f := 1146;
        ELSIF x = 489 THEN
            sigmoid_f := 1146;
        ELSIF x = 490 THEN
            sigmoid_f := 1146;
        ELSIF x = 491 THEN
            sigmoid_f := 1146;
        ELSIF x = 492 THEN
            sigmoid_f := 1147;
        ELSIF x = 493 THEN
            sigmoid_f := 1147;
        ELSIF x = 494 THEN
            sigmoid_f := 1147;
        ELSIF x = 495 THEN
            sigmoid_f := 1147;
        ELSIF x = 496 THEN
            sigmoid_f := 1148;
        ELSIF x = 497 THEN
            sigmoid_f := 1148;
        ELSIF x = 498 THEN
            sigmoid_f := 1148;
        ELSIF x = 499 THEN
            sigmoid_f := 1148;
        ELSIF x = 500 THEN
            sigmoid_f := 1149;
        ELSIF x = 501 THEN
            sigmoid_f := 1149;
        ELSIF x = 502 THEN
            sigmoid_f := 1149;
        ELSIF x = 503 THEN
            sigmoid_f := 1149;
        ELSIF x = 504 THEN
            sigmoid_f := 1150;
        ELSIF x = 505 THEN
            sigmoid_f := 1150;
        ELSIF x = 506 THEN
            sigmoid_f := 1150;
        ELSIF x = 507 THEN
            sigmoid_f := 1150;
        ELSIF x = 508 THEN
            sigmoid_f := 1151;
        ELSIF x = 509 THEN
            sigmoid_f := 1151;
        ELSIF x = 510 THEN
            sigmoid_f := 1151;
        ELSIF x = 511 THEN
            sigmoid_f := 1151;
        ELSIF x = 512 THEN
            sigmoid_f := 1151;
        ELSIF x = 513 THEN
            sigmoid_f := 1151;
        ELSIF x = 514 THEN
            sigmoid_f := 1152;
        ELSIF x = 515 THEN
            sigmoid_f := 1152;
        ELSIF x = 516 THEN
            sigmoid_f := 1152;
        ELSIF x = 517 THEN
            sigmoid_f := 1152;
        ELSIF x = 518 THEN
            sigmoid_f := 1153;
        ELSIF x = 519 THEN
            sigmoid_f := 1153;
        ELSIF x = 520 THEN
            sigmoid_f := 1153;
        ELSIF x = 521 THEN
            sigmoid_f := 1153;
        ELSIF x = 522 THEN
            sigmoid_f := 1154;
        ELSIF x = 523 THEN
            sigmoid_f := 1154;
        ELSIF x = 524 THEN
            sigmoid_f := 1154;
        ELSIF x = 525 THEN
            sigmoid_f := 1154;
        ELSIF x = 526 THEN
            sigmoid_f := 1155;
        ELSIF x = 527 THEN
            sigmoid_f := 1155;
        ELSIF x = 528 THEN
            sigmoid_f := 1155;
        ELSIF x = 529 THEN
            sigmoid_f := 1155;
        ELSIF x = 530 THEN
            sigmoid_f := 1156;
        ELSIF x = 531 THEN
            sigmoid_f := 1156;
        ELSIF x = 532 THEN
            sigmoid_f := 1156;
        ELSIF x = 533 THEN
            sigmoid_f := 1156;
        ELSIF x = 534 THEN
            sigmoid_f := 1157;
        ELSIF x = 535 THEN
            sigmoid_f := 1157;
        ELSIF x = 536 THEN
            sigmoid_f := 1157;
        ELSIF x = 537 THEN
            sigmoid_f := 1157;
        ELSIF x = 538 THEN
            sigmoid_f := 1158;
        ELSIF x = 539 THEN
            sigmoid_f := 1158;
        ELSIF x = 540 THEN
            sigmoid_f := 1158;
        ELSIF x = 541 THEN
            sigmoid_f := 1158;
        ELSIF x = 542 THEN
            sigmoid_f := 1159;
        ELSIF x = 543 THEN
            sigmoid_f := 1159;
        ELSIF x = 544 THEN
            sigmoid_f := 1159;
        ELSIF x = 545 THEN
            sigmoid_f := 1159;
        ELSIF x = 546 THEN
            sigmoid_f := 1159;
        ELSIF x = 547 THEN
            sigmoid_f := 1160;
        ELSIF x = 548 THEN
            sigmoid_f := 1160;
        ELSIF x = 549 THEN
            sigmoid_f := 1160;
        ELSIF x = 550 THEN
            sigmoid_f := 1160;
        ELSIF x = 551 THEN
            sigmoid_f := 1161;
        ELSIF x = 552 THEN
            sigmoid_f := 1161;
        ELSIF x = 553 THEN
            sigmoid_f := 1161;
        ELSIF x = 554 THEN
            sigmoid_f := 1161;
        ELSIF x = 555 THEN
            sigmoid_f := 1162;
        ELSIF x = 556 THEN
            sigmoid_f := 1162;
        ELSIF x = 557 THEN
            sigmoid_f := 1162;
        ELSIF x = 558 THEN
            sigmoid_f := 1162;
        ELSIF x = 559 THEN
            sigmoid_f := 1163;
        ELSIF x = 560 THEN
            sigmoid_f := 1163;
        ELSIF x = 561 THEN
            sigmoid_f := 1163;
        ELSIF x = 562 THEN
            sigmoid_f := 1163;
        ELSIF x = 563 THEN
            sigmoid_f := 1164;
        ELSIF x = 564 THEN
            sigmoid_f := 1164;
        ELSIF x = 565 THEN
            sigmoid_f := 1164;
        ELSIF x = 566 THEN
            sigmoid_f := 1164;
        ELSIF x = 567 THEN
            sigmoid_f := 1165;
        ELSIF x = 568 THEN
            sigmoid_f := 1165;
        ELSIF x = 569 THEN
            sigmoid_f := 1165;
        ELSIF x = 570 THEN
            sigmoid_f := 1165;
        ELSIF x = 571 THEN
            sigmoid_f := 1166;
        ELSIF x = 572 THEN
            sigmoid_f := 1166;
        ELSIF x = 573 THEN
            sigmoid_f := 1166;
        ELSIF x = 574 THEN
            sigmoid_f := 1166;
        ELSIF x = 575 THEN
            sigmoid_f := 1166;
        ELSIF x = 576 THEN
            sigmoid_f := 1167;
        ELSIF x = 577 THEN
            sigmoid_f := 1167;
        ELSIF x = 578 THEN
            sigmoid_f := 1167;
        ELSIF x = 579 THEN
            sigmoid_f := 1167;
        ELSIF x = 580 THEN
            sigmoid_f := 1168;
        ELSIF x = 581 THEN
            sigmoid_f := 1168;
        ELSIF x = 582 THEN
            sigmoid_f := 1168;
        ELSIF x = 583 THEN
            sigmoid_f := 1168;
        ELSIF x = 584 THEN
            sigmoid_f := 1169;
        ELSIF x = 585 THEN
            sigmoid_f := 1169;
        ELSIF x = 586 THEN
            sigmoid_f := 1169;
        ELSIF x = 587 THEN
            sigmoid_f := 1169;
        ELSIF x = 588 THEN
            sigmoid_f := 1170;
        ELSIF x = 589 THEN
            sigmoid_f := 1170;
        ELSIF x = 590 THEN
            sigmoid_f := 1170;
        ELSIF x = 591 THEN
            sigmoid_f := 1170;
        ELSIF x = 592 THEN
            sigmoid_f := 1171;
        ELSIF x = 593 THEN
            sigmoid_f := 1171;
        ELSIF x = 594 THEN
            sigmoid_f := 1171;
        ELSIF x = 595 THEN
            sigmoid_f := 1171;
        ELSIF x = 596 THEN
            sigmoid_f := 1172;
        ELSIF x = 597 THEN
            sigmoid_f := 1172;
        ELSIF x = 598 THEN
            sigmoid_f := 1172;
        ELSIF x = 599 THEN
            sigmoid_f := 1172;
        ELSIF x = 600 THEN
            sigmoid_f := 1173;
        ELSIF x = 601 THEN
            sigmoid_f := 1173;
        ELSIF x = 602 THEN
            sigmoid_f := 1173;
        ELSIF x = 603 THEN
            sigmoid_f := 1173;
        ELSIF x = 604 THEN
            sigmoid_f := 1173;
        ELSIF x = 605 THEN
            sigmoid_f := 1174;
        ELSIF x = 606 THEN
            sigmoid_f := 1174;
        ELSIF x = 607 THEN
            sigmoid_f := 1174;
        ELSIF x = 608 THEN
            sigmoid_f := 1174;
        ELSIF x = 609 THEN
            sigmoid_f := 1175;
        ELSIF x = 610 THEN
            sigmoid_f := 1175;
        ELSIF x = 611 THEN
            sigmoid_f := 1175;
        ELSIF x = 612 THEN
            sigmoid_f := 1175;
        ELSIF x = 613 THEN
            sigmoid_f := 1176;
        ELSIF x = 614 THEN
            sigmoid_f := 1176;
        ELSIF x = 615 THEN
            sigmoid_f := 1176;
        ELSIF x = 616 THEN
            sigmoid_f := 1176;
        ELSIF x = 617 THEN
            sigmoid_f := 1177;
        ELSIF x = 618 THEN
            sigmoid_f := 1177;
        ELSIF x = 619 THEN
            sigmoid_f := 1177;
        ELSIF x = 620 THEN
            sigmoid_f := 1177;
        ELSIF x = 621 THEN
            sigmoid_f := 1178;
        ELSIF x = 622 THEN
            sigmoid_f := 1178;
        ELSIF x = 623 THEN
            sigmoid_f := 1178;
        ELSIF x = 624 THEN
            sigmoid_f := 1178;
        ELSIF x = 625 THEN
            sigmoid_f := 1179;
        ELSIF x = 626 THEN
            sigmoid_f := 1179;
        ELSIF x = 627 THEN
            sigmoid_f := 1179;
        ELSIF x = 628 THEN
            sigmoid_f := 1179;
        ELSIF x = 629 THEN
            sigmoid_f := 1180;
        ELSIF x = 630 THEN
            sigmoid_f := 1180;
        ELSIF x = 631 THEN
            sigmoid_f := 1180;
        ELSIF x = 632 THEN
            sigmoid_f := 1180;
        ELSIF x = 633 THEN
            sigmoid_f := 1180;
        ELSIF x = 634 THEN
            sigmoid_f := 1181;
        ELSIF x = 635 THEN
            sigmoid_f := 1181;
        ELSIF x = 636 THEN
            sigmoid_f := 1181;
        ELSIF x = 637 THEN
            sigmoid_f := 1181;
        ELSIF x = 638 THEN
            sigmoid_f := 1182;
        ELSIF x = 639 THEN
            sigmoid_f := 1182;
        ELSIF x = 640 THEN
            sigmoid_f := 1182;
        ELSIF x = 641 THEN
            sigmoid_f := 1182;
        ELSIF x = 642 THEN
            sigmoid_f := 1183;
        ELSIF x = 643 THEN
            sigmoid_f := 1183;
        ELSIF x = 644 THEN
            sigmoid_f := 1183;
        ELSIF x = 645 THEN
            sigmoid_f := 1183;
        ELSIF x = 646 THEN
            sigmoid_f := 1184;
        ELSIF x = 647 THEN
            sigmoid_f := 1184;
        ELSIF x = 648 THEN
            sigmoid_f := 1184;
        ELSIF x = 649 THEN
            sigmoid_f := 1184;
        ELSIF x = 650 THEN
            sigmoid_f := 1185;
        ELSIF x = 651 THEN
            sigmoid_f := 1185;
        ELSIF x = 652 THEN
            sigmoid_f := 1185;
        ELSIF x = 653 THEN
            sigmoid_f := 1185;
        ELSIF x = 654 THEN
            sigmoid_f := 1186;
        ELSIF x = 655 THEN
            sigmoid_f := 1186;
        ELSIF x = 656 THEN
            sigmoid_f := 1186;
        ELSIF x = 657 THEN
            sigmoid_f := 1186;
        ELSIF x = 658 THEN
            sigmoid_f := 1187;
        ELSIF x = 659 THEN
            sigmoid_f := 1187;
        ELSIF x = 660 THEN
            sigmoid_f := 1187;
        ELSIF x = 661 THEN
            sigmoid_f := 1187;
        ELSIF x = 662 THEN
            sigmoid_f := 1188;
        ELSIF x = 663 THEN
            sigmoid_f := 1188;
        ELSIF x = 664 THEN
            sigmoid_f := 1188;
        ELSIF x = 665 THEN
            sigmoid_f := 1188;
        ELSIF x = 666 THEN
            sigmoid_f := 1188;
        ELSIF x = 667 THEN
            sigmoid_f := 1189;
        ELSIF x = 668 THEN
            sigmoid_f := 1189;
        ELSIF x = 669 THEN
            sigmoid_f := 1189;
        ELSIF x = 670 THEN
            sigmoid_f := 1189;
        ELSIF x = 671 THEN
            sigmoid_f := 1190;
        ELSIF x = 672 THEN
            sigmoid_f := 1190;
        ELSIF x = 673 THEN
            sigmoid_f := 1190;
        ELSIF x = 674 THEN
            sigmoid_f := 1190;
        ELSIF x = 675 THEN
            sigmoid_f := 1191;
        ELSIF x = 676 THEN
            sigmoid_f := 1191;
        ELSIF x = 677 THEN
            sigmoid_f := 1191;
        ELSIF x = 678 THEN
            sigmoid_f := 1191;
        ELSIF x = 679 THEN
            sigmoid_f := 1192;
        ELSIF x = 680 THEN
            sigmoid_f := 1192;
        ELSIF x = 681 THEN
            sigmoid_f := 1192;
        ELSIF x = 682 THEN
            sigmoid_f := 1192;
        ELSIF x = 683 THEN
            sigmoid_f := 1193;
        ELSIF x = 684 THEN
            sigmoid_f := 1193;
        ELSIF x = 685 THEN
            sigmoid_f := 1193;
        ELSIF x = 686 THEN
            sigmoid_f := 1193;
        ELSIF x = 687 THEN
            sigmoid_f := 1194;
        ELSIF x = 688 THEN
            sigmoid_f := 1194;
        ELSIF x = 689 THEN
            sigmoid_f := 1194;
        ELSIF x = 690 THEN
            sigmoid_f := 1194;
        ELSIF x = 691 THEN
            sigmoid_f := 1195;
        ELSIF x = 692 THEN
            sigmoid_f := 1195;
        ELSIF x = 693 THEN
            sigmoid_f := 1195;
        ELSIF x = 694 THEN
            sigmoid_f := 1195;
        ELSIF x = 695 THEN
            sigmoid_f := 1195;
        ELSIF x = 696 THEN
            sigmoid_f := 1196;
        ELSIF x = 697 THEN
            sigmoid_f := 1196;
        ELSIF x = 698 THEN
            sigmoid_f := 1196;
        ELSIF x = 699 THEN
            sigmoid_f := 1196;
        ELSIF x = 700 THEN
            sigmoid_f := 1197;
        ELSIF x = 701 THEN
            sigmoid_f := 1197;
        ELSIF x = 702 THEN
            sigmoid_f := 1197;
        ELSIF x = 703 THEN
            sigmoid_f := 1197;
        ELSIF x = 704 THEN
            sigmoid_f := 1198;
        ELSIF x = 705 THEN
            sigmoid_f := 1198;
        ELSIF x = 706 THEN
            sigmoid_f := 1198;
        ELSIF x = 707 THEN
            sigmoid_f := 1198;
        ELSIF x = 708 THEN
            sigmoid_f := 1199;
        ELSIF x = 709 THEN
            sigmoid_f := 1199;
        ELSIF x = 710 THEN
            sigmoid_f := 1199;
        ELSIF x = 711 THEN
            sigmoid_f := 1199;
        ELSIF x = 712 THEN
            sigmoid_f := 1200;
        ELSIF x = 713 THEN
            sigmoid_f := 1200;
        ELSIF x = 714 THEN
            sigmoid_f := 1200;
        ELSIF x = 715 THEN
            sigmoid_f := 1200;
        ELSIF x = 716 THEN
            sigmoid_f := 1201;
        ELSIF x = 717 THEN
            sigmoid_f := 1201;
        ELSIF x = 718 THEN
            sigmoid_f := 1201;
        ELSIF x = 719 THEN
            sigmoid_f := 1201;
        ELSIF x = 720 THEN
            sigmoid_f := 1202;
        ELSIF x = 721 THEN
            sigmoid_f := 1202;
        ELSIF x = 722 THEN
            sigmoid_f := 1202;
        ELSIF x = 723 THEN
            sigmoid_f := 1202;
        ELSIF x = 724 THEN
            sigmoid_f := 1202;
        ELSIF x = 725 THEN
            sigmoid_f := 1203;
        ELSIF x = 726 THEN
            sigmoid_f := 1203;
        ELSIF x = 727 THEN
            sigmoid_f := 1203;
        ELSIF x = 728 THEN
            sigmoid_f := 1203;
        ELSIF x = 729 THEN
            sigmoid_f := 1204;
        ELSIF x = 730 THEN
            sigmoid_f := 1204;
        ELSIF x = 731 THEN
            sigmoid_f := 1204;
        ELSIF x = 732 THEN
            sigmoid_f := 1204;
        ELSIF x = 733 THEN
            sigmoid_f := 1205;
        ELSIF x = 734 THEN
            sigmoid_f := 1205;
        ELSIF x = 735 THEN
            sigmoid_f := 1205;
        ELSIF x = 736 THEN
            sigmoid_f := 1205;
        ELSIF x = 737 THEN
            sigmoid_f := 1206;
        ELSIF x = 738 THEN
            sigmoid_f := 1206;
        ELSIF x = 739 THEN
            sigmoid_f := 1206;
        ELSIF x = 740 THEN
            sigmoid_f := 1206;
        ELSIF x = 741 THEN
            sigmoid_f := 1207;
        ELSIF x = 742 THEN
            sigmoid_f := 1207;
        ELSIF x = 743 THEN
            sigmoid_f := 1207;
        ELSIF x = 744 THEN
            sigmoid_f := 1207;
        ELSIF x = 745 THEN
            sigmoid_f := 1208;
        ELSIF x = 746 THEN
            sigmoid_f := 1208;
        ELSIF x = 747 THEN
            sigmoid_f := 1208;
        ELSIF x = 748 THEN
            sigmoid_f := 1208;
        ELSIF x = 749 THEN
            sigmoid_f := 1209;
        ELSIF x = 750 THEN
            sigmoid_f := 1209;
        ELSIF x = 751 THEN
            sigmoid_f := 1209;
        ELSIF x = 752 THEN
            sigmoid_f := 1209;
        ELSIF x = 753 THEN
            sigmoid_f := 1209;
        ELSIF x = 754 THEN
            sigmoid_f := 1210;
        ELSIF x = 755 THEN
            sigmoid_f := 1210;
        ELSIF x = 756 THEN
            sigmoid_f := 1210;
        ELSIF x = 757 THEN
            sigmoid_f := 1210;
        ELSIF x = 758 THEN
            sigmoid_f := 1211;
        ELSIF x = 759 THEN
            sigmoid_f := 1211;
        ELSIF x = 760 THEN
            sigmoid_f := 1211;
        ELSIF x = 761 THEN
            sigmoid_f := 1211;
        ELSIF x = 762 THEN
            sigmoid_f := 1212;
        ELSIF x = 763 THEN
            sigmoid_f := 1212;
        ELSIF x = 764 THEN
            sigmoid_f := 1212;
        ELSIF x = 765 THEN
            sigmoid_f := 1212;
        ELSIF x = 766 THEN
            sigmoid_f := 1213;
        ELSIF x = 767 THEN
            sigmoid_f := 1213;
        ELSIF x = 768 THEN
            sigmoid_f := 1213;
        ELSIF x = 769 THEN
            sigmoid_f := 1213;
        ELSIF x = 770 THEN
            sigmoid_f := 1214;
        ELSIF x = 771 THEN
            sigmoid_f := 1214;
        ELSIF x = 772 THEN
            sigmoid_f := 1214;
        ELSIF x = 773 THEN
            sigmoid_f := 1214;
        ELSIF x = 774 THEN
            sigmoid_f := 1215;
        ELSIF x = 775 THEN
            sigmoid_f := 1215;
        ELSIF x = 776 THEN
            sigmoid_f := 1215;
        ELSIF x = 777 THEN
            sigmoid_f := 1215;
        ELSIF x = 778 THEN
            sigmoid_f := 1216;
        ELSIF x = 779 THEN
            sigmoid_f := 1216;
        ELSIF x = 780 THEN
            sigmoid_f := 1216;
        ELSIF x = 781 THEN
            sigmoid_f := 1216;
        ELSIF x = 782 THEN
            sigmoid_f := 1217;
        ELSIF x = 783 THEN
            sigmoid_f := 1217;
        ELSIF x = 784 THEN
            sigmoid_f := 1217;
        ELSIF x = 785 THEN
            sigmoid_f := 1217;
        ELSIF x = 786 THEN
            sigmoid_f := 1217;
        ELSIF x = 787 THEN
            sigmoid_f := 1218;
        ELSIF x = 788 THEN
            sigmoid_f := 1218;
        ELSIF x = 789 THEN
            sigmoid_f := 1218;
        ELSIF x = 790 THEN
            sigmoid_f := 1218;
        ELSIF x = 791 THEN
            sigmoid_f := 1219;
        ELSIF x = 792 THEN
            sigmoid_f := 1219;
        ELSIF x = 793 THEN
            sigmoid_f := 1219;
        ELSIF x = 794 THEN
            sigmoid_f := 1219;
        ELSIF x = 795 THEN
            sigmoid_f := 1220;
        ELSIF x = 796 THEN
            sigmoid_f := 1220;
        ELSIF x = 797 THEN
            sigmoid_f := 1220;
        ELSIF x = 798 THEN
            sigmoid_f := 1220;
        ELSIF x = 799 THEN
            sigmoid_f := 1221;
        ELSIF x = 800 THEN
            sigmoid_f := 1221;
        ELSIF x = 801 THEN
            sigmoid_f := 1221;
        ELSIF x = 802 THEN
            sigmoid_f := 1221;
        ELSIF x = 803 THEN
            sigmoid_f := 1222;
        ELSIF x = 804 THEN
            sigmoid_f := 1222;
        ELSIF x = 805 THEN
            sigmoid_f := 1222;
        ELSIF x = 806 THEN
            sigmoid_f := 1222;
        ELSIF x = 807 THEN
            sigmoid_f := 1223;
        ELSIF x = 808 THEN
            sigmoid_f := 1223;
        ELSIF x = 809 THEN
            sigmoid_f := 1223;
        ELSIF x = 810 THEN
            sigmoid_f := 1223;
        ELSIF x = 811 THEN
            sigmoid_f := 1224;
        ELSIF x = 812 THEN
            sigmoid_f := 1224;
        ELSIF x = 813 THEN
            sigmoid_f := 1224;
        ELSIF x = 814 THEN
            sigmoid_f := 1224;
        ELSIF x = 815 THEN
            sigmoid_f := 1224;
        ELSIF x = 816 THEN
            sigmoid_f := 1225;
        ELSIF x = 817 THEN
            sigmoid_f := 1225;
        ELSIF x = 818 THEN
            sigmoid_f := 1225;
        ELSIF x = 819 THEN
            sigmoid_f := 1225;
        ELSIF x = 820 THEN
            sigmoid_f := 1226;
        ELSIF x = 821 THEN
            sigmoid_f := 1226;
        ELSIF x = 822 THEN
            sigmoid_f := 1226;
        ELSIF x = 823 THEN
            sigmoid_f := 1226;
        ELSIF x = 824 THEN
            sigmoid_f := 1227;
        ELSIF x = 825 THEN
            sigmoid_f := 1227;
        ELSIF x = 826 THEN
            sigmoid_f := 1227;
        ELSIF x = 827 THEN
            sigmoid_f := 1227;
        ELSIF x = 828 THEN
            sigmoid_f := 1228;
        ELSIF x = 829 THEN
            sigmoid_f := 1228;
        ELSIF x = 830 THEN
            sigmoid_f := 1228;
        ELSIF x = 831 THEN
            sigmoid_f := 1228;
        ELSIF x = 832 THEN
            sigmoid_f := 1229;
        ELSIF x = 833 THEN
            sigmoid_f := 1229;
        ELSIF x = 834 THEN
            sigmoid_f := 1229;
        ELSIF x = 835 THEN
            sigmoid_f := 1229;
        ELSIF x = 836 THEN
            sigmoid_f := 1230;
        ELSIF x = 837 THEN
            sigmoid_f := 1230;
        ELSIF x = 838 THEN
            sigmoid_f := 1230;
        ELSIF x = 839 THEN
            sigmoid_f := 1230;
        ELSIF x = 840 THEN
            sigmoid_f := 1231;
        ELSIF x = 841 THEN
            sigmoid_f := 1231;
        ELSIF x = 842 THEN
            sigmoid_f := 1231;
        ELSIF x = 843 THEN
            sigmoid_f := 1231;
        ELSIF x = 844 THEN
            sigmoid_f := 1231;
        ELSIF x = 845 THEN
            sigmoid_f := 1232;
        ELSIF x = 846 THEN
            sigmoid_f := 1232;
        ELSIF x = 847 THEN
            sigmoid_f := 1232;
        ELSIF x = 848 THEN
            sigmoid_f := 1232;
        ELSIF x = 849 THEN
            sigmoid_f := 1233;
        ELSIF x = 850 THEN
            sigmoid_f := 1233;
        ELSIF x = 851 THEN
            sigmoid_f := 1233;
        ELSIF x = 852 THEN
            sigmoid_f := 1233;
        ELSIF x = 853 THEN
            sigmoid_f := 1234;
        ELSIF x = 854 THEN
            sigmoid_f := 1234;
        ELSIF x = 855 THEN
            sigmoid_f := 1234;
        ELSIF x = 856 THEN
            sigmoid_f := 1234;
        ELSIF x = 857 THEN
            sigmoid_f := 1235;
        ELSIF x = 858 THEN
            sigmoid_f := 1235;
        ELSIF x = 859 THEN
            sigmoid_f := 1235;
        ELSIF x = 860 THEN
            sigmoid_f := 1235;
        ELSIF x = 861 THEN
            sigmoid_f := 1236;
        ELSIF x = 862 THEN
            sigmoid_f := 1236;
        ELSIF x = 863 THEN
            sigmoid_f := 1236;
        ELSIF x = 864 THEN
            sigmoid_f := 1236;
        ELSIF x = 865 THEN
            sigmoid_f := 1237;
        ELSIF x = 866 THEN
            sigmoid_f := 1237;
        ELSIF x = 867 THEN
            sigmoid_f := 1237;
        ELSIF x = 868 THEN
            sigmoid_f := 1237;
        ELSIF x = 869 THEN
            sigmoid_f := 1238;
        ELSIF x = 870 THEN
            sigmoid_f := 1238;
        ELSIF x = 871 THEN
            sigmoid_f := 1238;
        ELSIF x = 872 THEN
            sigmoid_f := 1238;
        ELSIF x = 873 THEN
            sigmoid_f := 1239;
        ELSIF x = 874 THEN
            sigmoid_f := 1239;
        ELSIF x = 875 THEN
            sigmoid_f := 1239;
        ELSIF x = 876 THEN
            sigmoid_f := 1239;
        ELSIF x = 877 THEN
            sigmoid_f := 1239;
        ELSIF x = 878 THEN
            sigmoid_f := 1240;
        ELSIF x = 879 THEN
            sigmoid_f := 1240;
        ELSIF x = 880 THEN
            sigmoid_f := 1240;
        ELSIF x = 881 THEN
            sigmoid_f := 1240;
        ELSIF x = 882 THEN
            sigmoid_f := 1241;
        ELSIF x = 883 THEN
            sigmoid_f := 1241;
        ELSIF x = 884 THEN
            sigmoid_f := 1241;
        ELSIF x = 885 THEN
            sigmoid_f := 1241;
        ELSIF x = 886 THEN
            sigmoid_f := 1242;
        ELSIF x = 887 THEN
            sigmoid_f := 1242;
        ELSIF x = 888 THEN
            sigmoid_f := 1242;
        ELSIF x = 889 THEN
            sigmoid_f := 1242;
        ELSIF x = 890 THEN
            sigmoid_f := 1243;
        ELSIF x = 891 THEN
            sigmoid_f := 1243;
        ELSIF x = 892 THEN
            sigmoid_f := 1243;
        ELSIF x = 893 THEN
            sigmoid_f := 1243;
        ELSIF x = 894 THEN
            sigmoid_f := 1244;
        ELSIF x = 895 THEN
            sigmoid_f := 1244;
        ELSIF x = 896 THEN
            sigmoid_f := 1244;
        ELSIF x = 897 THEN
            sigmoid_f := 1244;
        ELSIF x = 898 THEN
            sigmoid_f := 1245;
        ELSIF x = 899 THEN
            sigmoid_f := 1245;
        ELSIF x = 900 THEN
            sigmoid_f := 1245;
        ELSIF x = 901 THEN
            sigmoid_f := 1245;
        ELSIF x = 902 THEN
            sigmoid_f := 1246;
        ELSIF x = 903 THEN
            sigmoid_f := 1246;
        ELSIF x = 904 THEN
            sigmoid_f := 1246;
        ELSIF x = 905 THEN
            sigmoid_f := 1246;
        ELSIF x = 906 THEN
            sigmoid_f := 1246;
        ELSIF x = 907 THEN
            sigmoid_f := 1247;
        ELSIF x = 908 THEN
            sigmoid_f := 1247;
        ELSIF x = 909 THEN
            sigmoid_f := 1247;
        ELSIF x = 910 THEN
            sigmoid_f := 1247;
        ELSIF x = 911 THEN
            sigmoid_f := 1248;
        ELSIF x = 912 THEN
            sigmoid_f := 1248;
        ELSIF x = 913 THEN
            sigmoid_f := 1248;
        ELSIF x = 914 THEN
            sigmoid_f := 1248;
        ELSIF x = 915 THEN
            sigmoid_f := 1249;
        ELSIF x = 916 THEN
            sigmoid_f := 1249;
        ELSIF x = 917 THEN
            sigmoid_f := 1249;
        ELSIF x = 918 THEN
            sigmoid_f := 1249;
        ELSIF x = 919 THEN
            sigmoid_f := 1250;
        ELSIF x = 920 THEN
            sigmoid_f := 1250;
        ELSIF x = 921 THEN
            sigmoid_f := 1250;
        ELSIF x = 922 THEN
            sigmoid_f := 1250;
        ELSIF x = 923 THEN
            sigmoid_f := 1251;
        ELSIF x = 924 THEN
            sigmoid_f := 1251;
        ELSIF x = 925 THEN
            sigmoid_f := 1251;
        ELSIF x = 926 THEN
            sigmoid_f := 1251;
        ELSIF x = 927 THEN
            sigmoid_f := 1252;
        ELSIF x = 928 THEN
            sigmoid_f := 1252;
        ELSIF x = 929 THEN
            sigmoid_f := 1252;
        ELSIF x = 930 THEN
            sigmoid_f := 1252;
        ELSIF x = 931 THEN
            sigmoid_f := 1253;
        ELSIF x = 932 THEN
            sigmoid_f := 1253;
        ELSIF x = 933 THEN
            sigmoid_f := 1253;
        ELSIF x = 934 THEN
            sigmoid_f := 1253;
        ELSIF x = 935 THEN
            sigmoid_f := 1253;
        ELSIF x = 936 THEN
            sigmoid_f := 1254;
        ELSIF x = 937 THEN
            sigmoid_f := 1254;
        ELSIF x = 938 THEN
            sigmoid_f := 1254;
        ELSIF x = 939 THEN
            sigmoid_f := 1254;
        ELSIF x = 940 THEN
            sigmoid_f := 1255;
        ELSIF x = 941 THEN
            sigmoid_f := 1255;
        ELSIF x = 942 THEN
            sigmoid_f := 1255;
        ELSIF x = 943 THEN
            sigmoid_f := 1255;
        ELSIF x = 944 THEN
            sigmoid_f := 1256;
        ELSIF x = 945 THEN
            sigmoid_f := 1256;
        ELSIF x = 946 THEN
            sigmoid_f := 1256;
        ELSIF x = 947 THEN
            sigmoid_f := 1256;
        ELSIF x = 948 THEN
            sigmoid_f := 1257;
        ELSIF x = 949 THEN
            sigmoid_f := 1257;
        ELSIF x = 950 THEN
            sigmoid_f := 1257;
        ELSIF x = 951 THEN
            sigmoid_f := 1257;
        ELSIF x = 952 THEN
            sigmoid_f := 1258;
        ELSIF x = 953 THEN
            sigmoid_f := 1258;
        ELSIF x = 954 THEN
            sigmoid_f := 1258;
        ELSIF x = 955 THEN
            sigmoid_f := 1258;
        ELSIF x = 956 THEN
            sigmoid_f := 1259;
        ELSIF x = 957 THEN
            sigmoid_f := 1259;
        ELSIF x = 958 THEN
            sigmoid_f := 1259;
        ELSIF x = 959 THEN
            sigmoid_f := 1259;
        ELSIF x = 960 THEN
            sigmoid_f := 1260;
        ELSIF x = 961 THEN
            sigmoid_f := 1260;
        ELSIF x = 962 THEN
            sigmoid_f := 1260;
        ELSIF x = 963 THEN
            sigmoid_f := 1260;
        ELSIF x = 964 THEN
            sigmoid_f := 1260;
        ELSIF x = 965 THEN
            sigmoid_f := 1261;
        ELSIF x = 966 THEN
            sigmoid_f := 1261;
        ELSIF x = 967 THEN
            sigmoid_f := 1261;
        ELSIF x = 968 THEN
            sigmoid_f := 1261;
        ELSIF x = 969 THEN
            sigmoid_f := 1262;
        ELSIF x = 970 THEN
            sigmoid_f := 1262;
        ELSIF x = 971 THEN
            sigmoid_f := 1262;
        ELSIF x = 972 THEN
            sigmoid_f := 1262;
        ELSIF x = 973 THEN
            sigmoid_f := 1263;
        ELSIF x = 974 THEN
            sigmoid_f := 1263;
        ELSIF x = 975 THEN
            sigmoid_f := 1263;
        ELSIF x = 976 THEN
            sigmoid_f := 1263;
        ELSIF x = 977 THEN
            sigmoid_f := 1264;
        ELSIF x = 978 THEN
            sigmoid_f := 1264;
        ELSIF x = 979 THEN
            sigmoid_f := 1264;
        ELSIF x = 980 THEN
            sigmoid_f := 1264;
        ELSIF x = 981 THEN
            sigmoid_f := 1265;
        ELSIF x = 982 THEN
            sigmoid_f := 1265;
        ELSIF x = 983 THEN
            sigmoid_f := 1265;
        ELSIF x = 984 THEN
            sigmoid_f := 1265;
        ELSIF x = 985 THEN
            sigmoid_f := 1266;
        ELSIF x = 986 THEN
            sigmoid_f := 1266;
        ELSIF x = 987 THEN
            sigmoid_f := 1266;
        ELSIF x = 988 THEN
            sigmoid_f := 1266;
        ELSIF x = 989 THEN
            sigmoid_f := 1267;
        ELSIF x = 990 THEN
            sigmoid_f := 1267;
        ELSIF x = 991 THEN
            sigmoid_f := 1267;
        ELSIF x = 992 THEN
            sigmoid_f := 1267;
        ELSIF x = 993 THEN
            sigmoid_f := 1268;
        ELSIF x = 994 THEN
            sigmoid_f := 1268;
        ELSIF x = 995 THEN
            sigmoid_f := 1268;
        ELSIF x = 996 THEN
            sigmoid_f := 1268;
        ELSIF x = 997 THEN
            sigmoid_f := 1268;
        ELSIF x = 998 THEN
            sigmoid_f := 1269;
        ELSIF x = 999 THEN
            sigmoid_f := 1269;
        ELSIF x = 1000 THEN
            sigmoid_f := 1269;
        ELSIF x = 1001 THEN
            sigmoid_f := 1269;
        ELSIF x = 1002 THEN
            sigmoid_f := 1270;
        ELSIF x = 1003 THEN
            sigmoid_f := 1270;
        ELSIF x = 1004 THEN
            sigmoid_f := 1270;
        ELSIF x = 1005 THEN
            sigmoid_f := 1270;
        ELSIF x = 1006 THEN
            sigmoid_f := 1271;
        ELSIF x = 1007 THEN
            sigmoid_f := 1271;
        ELSIF x = 1008 THEN
            sigmoid_f := 1271;
        ELSIF x = 1009 THEN
            sigmoid_f := 1271;
        ELSIF x = 1010 THEN
            sigmoid_f := 1272;
        ELSIF x = 1011 THEN
            sigmoid_f := 1272;
        ELSIF x = 1012 THEN
            sigmoid_f := 1272;
        ELSIF x = 1013 THEN
            sigmoid_f := 1272;
        ELSIF x = 1014 THEN
            sigmoid_f := 1273;
        ELSIF x = 1015 THEN
            sigmoid_f := 1273;
        ELSIF x = 1016 THEN
            sigmoid_f := 1273;
        ELSIF x = 1017 THEN
            sigmoid_f := 1273;
        ELSIF x = 1018 THEN
            sigmoid_f := 1274;
        ELSIF x = 1019 THEN
            sigmoid_f := 1274;
        ELSIF x = 1020 THEN
            sigmoid_f := 1274;
        ELSIF x = 1021 THEN
            sigmoid_f := 1274;
        ELSIF x = 1022 THEN
            sigmoid_f := 1275;
        ELSIF x = 1023 THEN
            sigmoid_f := 1275;
        ELSIF x = 1024 THEN
            sigmoid_f := 1275;
        ELSIF x = 1025 THEN
            sigmoid_f := 1275;
        ELSIF x = 1026 THEN
            sigmoid_f := 1275;
        ELSIF x = 1027 THEN
            sigmoid_f := 1276;
        ELSIF x = 1028 THEN
            sigmoid_f := 1276;
        ELSIF x = 1029 THEN
            sigmoid_f := 1276;
        ELSIF x = 1030 THEN
            sigmoid_f := 1276;
        ELSIF x = 1031 THEN
            sigmoid_f := 1277;
        ELSIF x = 1032 THEN
            sigmoid_f := 1277;
        ELSIF x = 1033 THEN
            sigmoid_f := 1277;
        ELSIF x = 1034 THEN
            sigmoid_f := 1277;
        ELSIF x = 1035 THEN
            sigmoid_f := 1277;
        ELSIF x = 1036 THEN
            sigmoid_f := 1278;
        ELSIF x = 1037 THEN
            sigmoid_f := 1278;
        ELSIF x = 1038 THEN
            sigmoid_f := 1278;
        ELSIF x = 1039 THEN
            sigmoid_f := 1278;
        ELSIF x = 1040 THEN
            sigmoid_f := 1279;
        ELSIF x = 1041 THEN
            sigmoid_f := 1279;
        ELSIF x = 1042 THEN
            sigmoid_f := 1279;
        ELSIF x = 1043 THEN
            sigmoid_f := 1279;
        ELSIF x = 1044 THEN
            sigmoid_f := 1280;
        ELSIF x = 1045 THEN
            sigmoid_f := 1280;
        ELSIF x = 1046 THEN
            sigmoid_f := 1280;
        ELSIF x = 1047 THEN
            sigmoid_f := 1280;
        ELSIF x = 1048 THEN
            sigmoid_f := 1280;
        ELSIF x = 1049 THEN
            sigmoid_f := 1281;
        ELSIF x = 1050 THEN
            sigmoid_f := 1281;
        ELSIF x = 1051 THEN
            sigmoid_f := 1281;
        ELSIF x = 1052 THEN
            sigmoid_f := 1281;
        ELSIF x = 1053 THEN
            sigmoid_f := 1282;
        ELSIF x = 1054 THEN
            sigmoid_f := 1282;
        ELSIF x = 1055 THEN
            sigmoid_f := 1282;
        ELSIF x = 1056 THEN
            sigmoid_f := 1282;
        ELSIF x = 1057 THEN
            sigmoid_f := 1282;
        ELSIF x = 1058 THEN
            sigmoid_f := 1283;
        ELSIF x = 1059 THEN
            sigmoid_f := 1283;
        ELSIF x = 1060 THEN
            sigmoid_f := 1283;
        ELSIF x = 1061 THEN
            sigmoid_f := 1283;
        ELSIF x = 1062 THEN
            sigmoid_f := 1284;
        ELSIF x = 1063 THEN
            sigmoid_f := 1284;
        ELSIF x = 1064 THEN
            sigmoid_f := 1284;
        ELSIF x = 1065 THEN
            sigmoid_f := 1284;
        ELSIF x = 1066 THEN
            sigmoid_f := 1285;
        ELSIF x = 1067 THEN
            sigmoid_f := 1285;
        ELSIF x = 1068 THEN
            sigmoid_f := 1285;
        ELSIF x = 1069 THEN
            sigmoid_f := 1285;
        ELSIF x = 1070 THEN
            sigmoid_f := 1285;
        ELSIF x = 1071 THEN
            sigmoid_f := 1286;
        ELSIF x = 1072 THEN
            sigmoid_f := 1286;
        ELSIF x = 1073 THEN
            sigmoid_f := 1286;
        ELSIF x = 1074 THEN
            sigmoid_f := 1286;
        ELSIF x = 1075 THEN
            sigmoid_f := 1287;
        ELSIF x = 1076 THEN
            sigmoid_f := 1287;
        ELSIF x = 1077 THEN
            sigmoid_f := 1287;
        ELSIF x = 1078 THEN
            sigmoid_f := 1287;
        ELSIF x = 1079 THEN
            sigmoid_f := 1287;
        ELSIF x = 1080 THEN
            sigmoid_f := 1288;
        ELSIF x = 1081 THEN
            sigmoid_f := 1288;
        ELSIF x = 1082 THEN
            sigmoid_f := 1288;
        ELSIF x = 1083 THEN
            sigmoid_f := 1288;
        ELSIF x = 1084 THEN
            sigmoid_f := 1289;
        ELSIF x = 1085 THEN
            sigmoid_f := 1289;
        ELSIF x = 1086 THEN
            sigmoid_f := 1289;
        ELSIF x = 1087 THEN
            sigmoid_f := 1289;
        ELSIF x = 1088 THEN
            sigmoid_f := 1290;
        ELSIF x = 1089 THEN
            sigmoid_f := 1290;
        ELSIF x = 1090 THEN
            sigmoid_f := 1290;
        ELSIF x = 1091 THEN
            sigmoid_f := 1290;
        ELSIF x = 1092 THEN
            sigmoid_f := 1290;
        ELSIF x = 1093 THEN
            sigmoid_f := 1291;
        ELSIF x = 1094 THEN
            sigmoid_f := 1291;
        ELSIF x = 1095 THEN
            sigmoid_f := 1291;
        ELSIF x = 1096 THEN
            sigmoid_f := 1291;
        ELSIF x = 1097 THEN
            sigmoid_f := 1292;
        ELSIF x = 1098 THEN
            sigmoid_f := 1292;
        ELSIF x = 1099 THEN
            sigmoid_f := 1292;
        ELSIF x = 1100 THEN
            sigmoid_f := 1292;
        ELSIF x = 1101 THEN
            sigmoid_f := 1292;
        ELSIF x = 1102 THEN
            sigmoid_f := 1293;
        ELSIF x = 1103 THEN
            sigmoid_f := 1293;
        ELSIF x = 1104 THEN
            sigmoid_f := 1293;
        ELSIF x = 1105 THEN
            sigmoid_f := 1293;
        ELSIF x = 1106 THEN
            sigmoid_f := 1294;
        ELSIF x = 1107 THEN
            sigmoid_f := 1294;
        ELSIF x = 1108 THEN
            sigmoid_f := 1294;
        ELSIF x = 1109 THEN
            sigmoid_f := 1294;
        ELSIF x = 1110 THEN
            sigmoid_f := 1295;
        ELSIF x = 1111 THEN
            sigmoid_f := 1295;
        ELSIF x = 1112 THEN
            sigmoid_f := 1295;
        ELSIF x = 1113 THEN
            sigmoid_f := 1295;
        ELSIF x = 1114 THEN
            sigmoid_f := 1295;
        ELSIF x = 1115 THEN
            sigmoid_f := 1296;
        ELSIF x = 1116 THEN
            sigmoid_f := 1296;
        ELSIF x = 1117 THEN
            sigmoid_f := 1296;
        ELSIF x = 1118 THEN
            sigmoid_f := 1296;
        ELSIF x = 1119 THEN
            sigmoid_f := 1297;
        ELSIF x = 1120 THEN
            sigmoid_f := 1297;
        ELSIF x = 1121 THEN
            sigmoid_f := 1297;
        ELSIF x = 1122 THEN
            sigmoid_f := 1297;
        ELSIF x = 1123 THEN
            sigmoid_f := 1297;
        ELSIF x = 1124 THEN
            sigmoid_f := 1298;
        ELSIF x = 1125 THEN
            sigmoid_f := 1298;
        ELSIF x = 1126 THEN
            sigmoid_f := 1298;
        ELSIF x = 1127 THEN
            sigmoid_f := 1298;
        ELSIF x = 1128 THEN
            sigmoid_f := 1299;
        ELSIF x = 1129 THEN
            sigmoid_f := 1299;
        ELSIF x = 1130 THEN
            sigmoid_f := 1299;
        ELSIF x = 1131 THEN
            sigmoid_f := 1299;
        ELSIF x = 1132 THEN
            sigmoid_f := 1300;
        ELSIF x = 1133 THEN
            sigmoid_f := 1300;
        ELSIF x = 1134 THEN
            sigmoid_f := 1300;
        ELSIF x = 1135 THEN
            sigmoid_f := 1300;
        ELSIF x = 1136 THEN
            sigmoid_f := 1300;
        ELSIF x = 1137 THEN
            sigmoid_f := 1301;
        ELSIF x = 1138 THEN
            sigmoid_f := 1301;
        ELSIF x = 1139 THEN
            sigmoid_f := 1301;
        ELSIF x = 1140 THEN
            sigmoid_f := 1301;
        ELSIF x = 1141 THEN
            sigmoid_f := 1302;
        ELSIF x = 1142 THEN
            sigmoid_f := 1302;
        ELSIF x = 1143 THEN
            sigmoid_f := 1302;
        ELSIF x = 1144 THEN
            sigmoid_f := 1302;
        ELSIF x = 1145 THEN
            sigmoid_f := 1302;
        ELSIF x = 1146 THEN
            sigmoid_f := 1303;
        ELSIF x = 1147 THEN
            sigmoid_f := 1303;
        ELSIF x = 1148 THEN
            sigmoid_f := 1303;
        ELSIF x = 1149 THEN
            sigmoid_f := 1303;
        ELSIF x = 1150 THEN
            sigmoid_f := 1304;
        ELSIF x = 1151 THEN
            sigmoid_f := 1304;
        ELSIF x = 1152 THEN
            sigmoid_f := 1304;
        ELSIF x = 1153 THEN
            sigmoid_f := 1304;
        ELSIF x = 1154 THEN
            sigmoid_f := 1305;
        ELSIF x = 1155 THEN
            sigmoid_f := 1305;
        ELSIF x = 1156 THEN
            sigmoid_f := 1305;
        ELSIF x = 1157 THEN
            sigmoid_f := 1305;
        ELSIF x = 1158 THEN
            sigmoid_f := 1305;
        ELSIF x = 1159 THEN
            sigmoid_f := 1306;
        ELSIF x = 1160 THEN
            sigmoid_f := 1306;
        ELSIF x = 1161 THEN
            sigmoid_f := 1306;
        ELSIF x = 1162 THEN
            sigmoid_f := 1306;
        ELSIF x = 1163 THEN
            sigmoid_f := 1307;
        ELSIF x = 1164 THEN
            sigmoid_f := 1307;
        ELSIF x = 1165 THEN
            sigmoid_f := 1307;
        ELSIF x = 1166 THEN
            sigmoid_f := 1307;
        ELSIF x = 1167 THEN
            sigmoid_f := 1307;
        ELSIF x = 1168 THEN
            sigmoid_f := 1308;
        ELSIF x = 1169 THEN
            sigmoid_f := 1308;
        ELSIF x = 1170 THEN
            sigmoid_f := 1308;
        ELSIF x = 1171 THEN
            sigmoid_f := 1308;
        ELSIF x = 1172 THEN
            sigmoid_f := 1309;
        ELSIF x = 1173 THEN
            sigmoid_f := 1309;
        ELSIF x = 1174 THEN
            sigmoid_f := 1309;
        ELSIF x = 1175 THEN
            sigmoid_f := 1309;
        ELSIF x = 1176 THEN
            sigmoid_f := 1310;
        ELSIF x = 1177 THEN
            sigmoid_f := 1310;
        ELSIF x = 1178 THEN
            sigmoid_f := 1310;
        ELSIF x = 1179 THEN
            sigmoid_f := 1310;
        ELSIF x = 1180 THEN
            sigmoid_f := 1310;
        ELSIF x = 1181 THEN
            sigmoid_f := 1311;
        ELSIF x = 1182 THEN
            sigmoid_f := 1311;
        ELSIF x = 1183 THEN
            sigmoid_f := 1311;
        ELSIF x = 1184 THEN
            sigmoid_f := 1311;
        ELSIF x = 1185 THEN
            sigmoid_f := 1312;
        ELSIF x = 1186 THEN
            sigmoid_f := 1312;
        ELSIF x = 1187 THEN
            sigmoid_f := 1312;
        ELSIF x = 1188 THEN
            sigmoid_f := 1312;
        ELSIF x = 1189 THEN
            sigmoid_f := 1312;
        ELSIF x = 1190 THEN
            sigmoid_f := 1313;
        ELSIF x = 1191 THEN
            sigmoid_f := 1313;
        ELSIF x = 1192 THEN
            sigmoid_f := 1313;
        ELSIF x = 1193 THEN
            sigmoid_f := 1313;
        ELSIF x = 1194 THEN
            sigmoid_f := 1314;
        ELSIF x = 1195 THEN
            sigmoid_f := 1314;
        ELSIF x = 1196 THEN
            sigmoid_f := 1314;
        ELSIF x = 1197 THEN
            sigmoid_f := 1314;
        ELSIF x = 1198 THEN
            sigmoid_f := 1315;
        ELSIF x = 1199 THEN
            sigmoid_f := 1315;
        ELSIF x = 1200 THEN
            sigmoid_f := 1315;
        ELSIF x = 1201 THEN
            sigmoid_f := 1315;
        ELSIF x = 1202 THEN
            sigmoid_f := 1315;
        ELSIF x = 1203 THEN
            sigmoid_f := 1316;
        ELSIF x = 1204 THEN
            sigmoid_f := 1316;
        ELSIF x = 1205 THEN
            sigmoid_f := 1316;
        ELSIF x = 1206 THEN
            sigmoid_f := 1316;
        ELSIF x = 1207 THEN
            sigmoid_f := 1317;
        ELSIF x = 1208 THEN
            sigmoid_f := 1317;
        ELSIF x = 1209 THEN
            sigmoid_f := 1317;
        ELSIF x = 1210 THEN
            sigmoid_f := 1317;
        ELSIF x = 1211 THEN
            sigmoid_f := 1317;
        ELSIF x = 1212 THEN
            sigmoid_f := 1318;
        ELSIF x = 1213 THEN
            sigmoid_f := 1318;
        ELSIF x = 1214 THEN
            sigmoid_f := 1318;
        ELSIF x = 1215 THEN
            sigmoid_f := 1318;
        ELSIF x = 1216 THEN
            sigmoid_f := 1319;
        ELSIF x = 1217 THEN
            sigmoid_f := 1319;
        ELSIF x = 1218 THEN
            sigmoid_f := 1319;
        ELSIF x = 1219 THEN
            sigmoid_f := 1319;
        ELSIF x = 1220 THEN
            sigmoid_f := 1320;
        ELSIF x = 1221 THEN
            sigmoid_f := 1320;
        ELSIF x = 1222 THEN
            sigmoid_f := 1320;
        ELSIF x = 1223 THEN
            sigmoid_f := 1320;
        ELSIF x = 1224 THEN
            sigmoid_f := 1320;
        ELSIF x = 1225 THEN
            sigmoid_f := 1321;
        ELSIF x = 1226 THEN
            sigmoid_f := 1321;
        ELSIF x = 1227 THEN
            sigmoid_f := 1321;
        ELSIF x = 1228 THEN
            sigmoid_f := 1321;
        ELSIF x = 1229 THEN
            sigmoid_f := 1322;
        ELSIF x = 1230 THEN
            sigmoid_f := 1322;
        ELSIF x = 1231 THEN
            sigmoid_f := 1322;
        ELSIF x = 1232 THEN
            sigmoid_f := 1322;
        ELSIF x = 1233 THEN
            sigmoid_f := 1322;
        ELSIF x = 1234 THEN
            sigmoid_f := 1323;
        ELSIF x = 1235 THEN
            sigmoid_f := 1323;
        ELSIF x = 1236 THEN
            sigmoid_f := 1323;
        ELSIF x = 1237 THEN
            sigmoid_f := 1323;
        ELSIF x = 1238 THEN
            sigmoid_f := 1324;
        ELSIF x = 1239 THEN
            sigmoid_f := 1324;
        ELSIF x = 1240 THEN
            sigmoid_f := 1324;
        ELSIF x = 1241 THEN
            sigmoid_f := 1324;
        ELSIF x = 1242 THEN
            sigmoid_f := 1324;
        ELSIF x = 1243 THEN
            sigmoid_f := 1325;
        ELSIF x = 1244 THEN
            sigmoid_f := 1325;
        ELSIF x = 1245 THEN
            sigmoid_f := 1325;
        ELSIF x = 1246 THEN
            sigmoid_f := 1325;
        ELSIF x = 1247 THEN
            sigmoid_f := 1326;
        ELSIF x = 1248 THEN
            sigmoid_f := 1326;
        ELSIF x = 1249 THEN
            sigmoid_f := 1326;
        ELSIF x = 1250 THEN
            sigmoid_f := 1326;
        ELSIF x = 1251 THEN
            sigmoid_f := 1327;
        ELSIF x = 1252 THEN
            sigmoid_f := 1327;
        ELSIF x = 1253 THEN
            sigmoid_f := 1327;
        ELSIF x = 1254 THEN
            sigmoid_f := 1327;
        ELSIF x = 1255 THEN
            sigmoid_f := 1327;
        ELSIF x = 1256 THEN
            sigmoid_f := 1328;
        ELSIF x = 1257 THEN
            sigmoid_f := 1328;
        ELSIF x = 1258 THEN
            sigmoid_f := 1328;
        ELSIF x = 1259 THEN
            sigmoid_f := 1328;
        ELSIF x = 1260 THEN
            sigmoid_f := 1329;
        ELSIF x = 1261 THEN
            sigmoid_f := 1329;
        ELSIF x = 1262 THEN
            sigmoid_f := 1329;
        ELSIF x = 1263 THEN
            sigmoid_f := 1329;
        ELSIF x = 1264 THEN
            sigmoid_f := 1329;
        ELSIF x = 1265 THEN
            sigmoid_f := 1330;
        ELSIF x = 1266 THEN
            sigmoid_f := 1330;
        ELSIF x = 1267 THEN
            sigmoid_f := 1330;
        ELSIF x = 1268 THEN
            sigmoid_f := 1330;
        ELSIF x = 1269 THEN
            sigmoid_f := 1331;
        ELSIF x = 1270 THEN
            sigmoid_f := 1331;
        ELSIF x = 1271 THEN
            sigmoid_f := 1331;
        ELSIF x = 1272 THEN
            sigmoid_f := 1331;
        ELSIF x = 1273 THEN
            sigmoid_f := 1332;
        ELSIF x = 1274 THEN
            sigmoid_f := 1332;
        ELSIF x = 1275 THEN
            sigmoid_f := 1332;
        ELSIF x = 1276 THEN
            sigmoid_f := 1332;
        ELSIF x = 1277 THEN
            sigmoid_f := 1332;
        ELSIF x = 1278 THEN
            sigmoid_f := 1333;
        ELSIF x = 1279 THEN
            sigmoid_f := 1333;
        ELSIF x = 1280 THEN
            sigmoid_f := 1333;
        ELSIF x = 1281 THEN
            sigmoid_f := 1333;
        ELSIF x = 1282 THEN
            sigmoid_f := 1334;
        ELSIF x = 1283 THEN
            sigmoid_f := 1334;
        ELSIF x = 1284 THEN
            sigmoid_f := 1334;
        ELSIF x = 1285 THEN
            sigmoid_f := 1334;
        ELSIF x = 1286 THEN
            sigmoid_f := 1334;
        ELSIF x = 1287 THEN
            sigmoid_f := 1335;
        ELSIF x = 1288 THEN
            sigmoid_f := 1335;
        ELSIF x = 1289 THEN
            sigmoid_f := 1335;
        ELSIF x = 1290 THEN
            sigmoid_f := 1335;
        ELSIF x = 1291 THEN
            sigmoid_f := 1336;
        ELSIF x = 1292 THEN
            sigmoid_f := 1336;
        ELSIF x = 1293 THEN
            sigmoid_f := 1336;
        ELSIF x = 1294 THEN
            sigmoid_f := 1336;
        ELSIF x = 1295 THEN
            sigmoid_f := 1337;
        ELSIF x = 1296 THEN
            sigmoid_f := 1337;
        ELSIF x = 1297 THEN
            sigmoid_f := 1337;
        ELSIF x = 1298 THEN
            sigmoid_f := 1337;
        ELSIF x = 1299 THEN
            sigmoid_f := 1337;
        ELSIF x = 1300 THEN
            sigmoid_f := 1338;
        ELSIF x = 1301 THEN
            sigmoid_f := 1338;
        ELSIF x = 1302 THEN
            sigmoid_f := 1338;
        ELSIF x = 1303 THEN
            sigmoid_f := 1338;
        ELSIF x = 1304 THEN
            sigmoid_f := 1339;
        ELSIF x = 1305 THEN
            sigmoid_f := 1339;
        ELSIF x = 1306 THEN
            sigmoid_f := 1339;
        ELSIF x = 1307 THEN
            sigmoid_f := 1339;
        ELSIF x = 1308 THEN
            sigmoid_f := 1339;
        ELSIF x = 1309 THEN
            sigmoid_f := 1340;
        ELSIF x = 1310 THEN
            sigmoid_f := 1340;
        ELSIF x = 1311 THEN
            sigmoid_f := 1340;
        ELSIF x = 1312 THEN
            sigmoid_f := 1340;
        ELSIF x = 1313 THEN
            sigmoid_f := 1341;
        ELSIF x = 1314 THEN
            sigmoid_f := 1341;
        ELSIF x = 1315 THEN
            sigmoid_f := 1341;
        ELSIF x = 1316 THEN
            sigmoid_f := 1341;
        ELSIF x = 1317 THEN
            sigmoid_f := 1342;
        ELSIF x = 1318 THEN
            sigmoid_f := 1342;
        ELSIF x = 1319 THEN
            sigmoid_f := 1342;
        ELSIF x = 1320 THEN
            sigmoid_f := 1342;
        ELSIF x = 1321 THEN
            sigmoid_f := 1342;
        ELSIF x = 1322 THEN
            sigmoid_f := 1343;
        ELSIF x = 1323 THEN
            sigmoid_f := 1343;
        ELSIF x = 1324 THEN
            sigmoid_f := 1343;
        ELSIF x = 1325 THEN
            sigmoid_f := 1343;
        ELSIF x = 1326 THEN
            sigmoid_f := 1344;
        ELSIF x = 1327 THEN
            sigmoid_f := 1344;
        ELSIF x = 1328 THEN
            sigmoid_f := 1344;
        ELSIF x = 1329 THEN
            sigmoid_f := 1344;
        ELSIF x = 1330 THEN
            sigmoid_f := 1344;
        ELSIF x = 1331 THEN
            sigmoid_f := 1345;
        ELSIF x = 1332 THEN
            sigmoid_f := 1345;
        ELSIF x = 1333 THEN
            sigmoid_f := 1345;
        ELSIF x = 1334 THEN
            sigmoid_f := 1345;
        ELSIF x = 1335 THEN
            sigmoid_f := 1346;
        ELSIF x = 1336 THEN
            sigmoid_f := 1346;
        ELSIF x = 1337 THEN
            sigmoid_f := 1346;
        ELSIF x = 1338 THEN
            sigmoid_f := 1346;
        ELSIF x = 1339 THEN
            sigmoid_f := 1347;
        ELSIF x = 1340 THEN
            sigmoid_f := 1347;
        ELSIF x = 1341 THEN
            sigmoid_f := 1347;
        ELSIF x = 1342 THEN
            sigmoid_f := 1347;
        ELSIF x = 1343 THEN
            sigmoid_f := 1347;
        ELSIF x = 1344 THEN
            sigmoid_f := 1348;
        ELSIF x = 1345 THEN
            sigmoid_f := 1348;
        ELSIF x = 1346 THEN
            sigmoid_f := 1348;
        ELSIF x = 1347 THEN
            sigmoid_f := 1348;
        ELSIF x = 1348 THEN
            sigmoid_f := 1349;
        ELSIF x = 1349 THEN
            sigmoid_f := 1349;
        ELSIF x = 1350 THEN
            sigmoid_f := 1349;
        ELSIF x = 1351 THEN
            sigmoid_f := 1349;
        ELSIF x = 1352 THEN
            sigmoid_f := 1349;
        ELSIF x = 1353 THEN
            sigmoid_f := 1350;
        ELSIF x = 1354 THEN
            sigmoid_f := 1350;
        ELSIF x = 1355 THEN
            sigmoid_f := 1350;
        ELSIF x = 1356 THEN
            sigmoid_f := 1350;
        ELSIF x = 1357 THEN
            sigmoid_f := 1351;
        ELSIF x = 1358 THEN
            sigmoid_f := 1351;
        ELSIF x = 1359 THEN
            sigmoid_f := 1351;
        ELSIF x = 1360 THEN
            sigmoid_f := 1351;
        ELSIF x = 1361 THEN
            sigmoid_f := 1352;
        ELSIF x = 1362 THEN
            sigmoid_f := 1352;
        ELSIF x = 1363 THEN
            sigmoid_f := 1352;
        ELSIF x = 1364 THEN
            sigmoid_f := 1352;
        ELSIF x = 1365 THEN
            sigmoid_f := 1352;
        ELSIF x = 1366 THEN
            sigmoid_f := 1353;
        ELSIF x = 1367 THEN
            sigmoid_f := 1353;
        ELSIF x = 1368 THEN
            sigmoid_f := 1353;
        ELSIF x = 1369 THEN
            sigmoid_f := 1353;
        ELSIF x = 1370 THEN
            sigmoid_f := 1354;
        ELSIF x = 1371 THEN
            sigmoid_f := 1354;
        ELSIF x = 1372 THEN
            sigmoid_f := 1354;
        ELSIF x = 1373 THEN
            sigmoid_f := 1354;
        ELSIF x = 1374 THEN
            sigmoid_f := 1354;
        ELSIF x = 1375 THEN
            sigmoid_f := 1355;
        ELSIF x = 1376 THEN
            sigmoid_f := 1355;
        ELSIF x = 1377 THEN
            sigmoid_f := 1355;
        ELSIF x = 1378 THEN
            sigmoid_f := 1355;
        ELSIF x = 1379 THEN
            sigmoid_f := 1356;
        ELSIF x = 1380 THEN
            sigmoid_f := 1356;
        ELSIF x = 1381 THEN
            sigmoid_f := 1356;
        ELSIF x = 1382 THEN
            sigmoid_f := 1356;
        ELSIF x = 1383 THEN
            sigmoid_f := 1357;
        ELSIF x = 1384 THEN
            sigmoid_f := 1357;
        ELSIF x = 1385 THEN
            sigmoid_f := 1357;
        ELSIF x = 1386 THEN
            sigmoid_f := 1357;
        ELSIF x = 1387 THEN
            sigmoid_f := 1357;
        ELSIF x = 1388 THEN
            sigmoid_f := 1358;
        ELSIF x = 1389 THEN
            sigmoid_f := 1358;
        ELSIF x = 1390 THEN
            sigmoid_f := 1358;
        ELSIF x = 1391 THEN
            sigmoid_f := 1358;
        ELSIF x = 1392 THEN
            sigmoid_f := 1359;
        ELSIF x = 1393 THEN
            sigmoid_f := 1359;
        ELSIF x = 1394 THEN
            sigmoid_f := 1359;
        ELSIF x = 1395 THEN
            sigmoid_f := 1359;
        ELSIF x = 1396 THEN
            sigmoid_f := 1359;
        ELSIF x = 1397 THEN
            sigmoid_f := 1360;
        ELSIF x = 1398 THEN
            sigmoid_f := 1360;
        ELSIF x = 1399 THEN
            sigmoid_f := 1360;
        ELSIF x = 1400 THEN
            sigmoid_f := 1360;
        ELSIF x = 1401 THEN
            sigmoid_f := 1361;
        ELSIF x = 1402 THEN
            sigmoid_f := 1361;
        ELSIF x = 1403 THEN
            sigmoid_f := 1361;
        ELSIF x = 1404 THEN
            sigmoid_f := 1361;
        ELSIF x = 1405 THEN
            sigmoid_f := 1362;
        ELSIF x = 1406 THEN
            sigmoid_f := 1362;
        ELSIF x = 1407 THEN
            sigmoid_f := 1362;
        ELSIF x = 1408 THEN
            sigmoid_f := 1362;
        ELSIF x = 1409 THEN
            sigmoid_f := 1362;
        ELSIF x = 1410 THEN
            sigmoid_f := 1363;
        ELSIF x = 1411 THEN
            sigmoid_f := 1363;
        ELSIF x = 1412 THEN
            sigmoid_f := 1363;
        ELSIF x = 1413 THEN
            sigmoid_f := 1363;
        ELSIF x = 1414 THEN
            sigmoid_f := 1364;
        ELSIF x = 1415 THEN
            sigmoid_f := 1364;
        ELSIF x = 1416 THEN
            sigmoid_f := 1364;
        ELSIF x = 1417 THEN
            sigmoid_f := 1364;
        ELSIF x = 1418 THEN
            sigmoid_f := 1364;
        ELSIF x = 1419 THEN
            sigmoid_f := 1365;
        ELSIF x = 1420 THEN
            sigmoid_f := 1365;
        ELSIF x = 1421 THEN
            sigmoid_f := 1365;
        ELSIF x = 1422 THEN
            sigmoid_f := 1365;
        ELSIF x = 1423 THEN
            sigmoid_f := 1366;
        ELSIF x = 1424 THEN
            sigmoid_f := 1366;
        ELSIF x = 1425 THEN
            sigmoid_f := 1366;
        ELSIF x = 1426 THEN
            sigmoid_f := 1366;
        ELSIF x = 1427 THEN
            sigmoid_f := 1367;
        ELSIF x = 1428 THEN
            sigmoid_f := 1367;
        ELSIF x = 1429 THEN
            sigmoid_f := 1367;
        ELSIF x = 1430 THEN
            sigmoid_f := 1367;
        ELSIF x = 1431 THEN
            sigmoid_f := 1367;
        ELSIF x = 1432 THEN
            sigmoid_f := 1368;
        ELSIF x = 1433 THEN
            sigmoid_f := 1368;
        ELSIF x = 1434 THEN
            sigmoid_f := 1368;
        ELSIF x = 1435 THEN
            sigmoid_f := 1368;
        ELSIF x = 1436 THEN
            sigmoid_f := 1369;
        ELSIF x = 1437 THEN
            sigmoid_f := 1369;
        ELSIF x = 1438 THEN
            sigmoid_f := 1369;
        ELSIF x = 1439 THEN
            sigmoid_f := 1369;
        ELSIF x = 1440 THEN
            sigmoid_f := 1369;
        ELSIF x = 1441 THEN
            sigmoid_f := 1370;
        ELSIF x = 1442 THEN
            sigmoid_f := 1370;
        ELSIF x = 1443 THEN
            sigmoid_f := 1370;
        ELSIF x = 1444 THEN
            sigmoid_f := 1370;
        ELSIF x = 1445 THEN
            sigmoid_f := 1371;
        ELSIF x = 1446 THEN
            sigmoid_f := 1371;
        ELSIF x = 1447 THEN
            sigmoid_f := 1371;
        ELSIF x = 1448 THEN
            sigmoid_f := 1371;
        ELSIF x = 1449 THEN
            sigmoid_f := 1371;
        ELSIF x = 1450 THEN
            sigmoid_f := 1372;
        ELSIF x = 1451 THEN
            sigmoid_f := 1372;
        ELSIF x = 1452 THEN
            sigmoid_f := 1372;
        ELSIF x = 1453 THEN
            sigmoid_f := 1372;
        ELSIF x = 1454 THEN
            sigmoid_f := 1373;
        ELSIF x = 1455 THEN
            sigmoid_f := 1373;
        ELSIF x = 1456 THEN
            sigmoid_f := 1373;
        ELSIF x = 1457 THEN
            sigmoid_f := 1373;
        ELSIF x = 1458 THEN
            sigmoid_f := 1374;
        ELSIF x = 1459 THEN
            sigmoid_f := 1374;
        ELSIF x = 1460 THEN
            sigmoid_f := 1374;
        ELSIF x = 1461 THEN
            sigmoid_f := 1374;
        ELSIF x = 1462 THEN
            sigmoid_f := 1374;
        ELSIF x = 1463 THEN
            sigmoid_f := 1375;
        ELSIF x = 1464 THEN
            sigmoid_f := 1375;
        ELSIF x = 1465 THEN
            sigmoid_f := 1375;
        ELSIF x = 1466 THEN
            sigmoid_f := 1375;
        ELSIF x = 1467 THEN
            sigmoid_f := 1376;
        ELSIF x = 1468 THEN
            sigmoid_f := 1376;
        ELSIF x = 1469 THEN
            sigmoid_f := 1376;
        ELSIF x = 1470 THEN
            sigmoid_f := 1376;
        ELSIF x = 1471 THEN
            sigmoid_f := 1376;
        ELSIF x = 1472 THEN
            sigmoid_f := 1377;
        ELSIF x = 1473 THEN
            sigmoid_f := 1377;
        ELSIF x = 1474 THEN
            sigmoid_f := 1377;
        ELSIF x = 1475 THEN
            sigmoid_f := 1377;
        ELSIF x = 1476 THEN
            sigmoid_f := 1378;
        ELSIF x = 1477 THEN
            sigmoid_f := 1378;
        ELSIF x = 1478 THEN
            sigmoid_f := 1378;
        ELSIF x = 1479 THEN
            sigmoid_f := 1378;
        ELSIF x = 1480 THEN
            sigmoid_f := 1379;
        ELSIF x = 1481 THEN
            sigmoid_f := 1379;
        ELSIF x = 1482 THEN
            sigmoid_f := 1379;
        ELSIF x = 1483 THEN
            sigmoid_f := 1379;
        ELSIF x = 1484 THEN
            sigmoid_f := 1379;
        ELSIF x = 1485 THEN
            sigmoid_f := 1380;
        ELSIF x = 1486 THEN
            sigmoid_f := 1380;
        ELSIF x = 1487 THEN
            sigmoid_f := 1380;
        ELSIF x = 1488 THEN
            sigmoid_f := 1380;
        ELSIF x = 1489 THEN
            sigmoid_f := 1381;
        ELSIF x = 1490 THEN
            sigmoid_f := 1381;
        ELSIF x = 1491 THEN
            sigmoid_f := 1381;
        ELSIF x = 1492 THEN
            sigmoid_f := 1381;
        ELSIF x = 1493 THEN
            sigmoid_f := 1381;
        ELSIF x = 1494 THEN
            sigmoid_f := 1382;
        ELSIF x = 1495 THEN
            sigmoid_f := 1382;
        ELSIF x = 1496 THEN
            sigmoid_f := 1382;
        ELSIF x = 1497 THEN
            sigmoid_f := 1382;
        ELSIF x = 1498 THEN
            sigmoid_f := 1383;
        ELSIF x = 1499 THEN
            sigmoid_f := 1383;
        ELSIF x = 1500 THEN
            sigmoid_f := 1383;
        ELSIF x = 1501 THEN
            sigmoid_f := 1383;
        ELSIF x = 1502 THEN
            sigmoid_f := 1384;
        ELSIF x = 1503 THEN
            sigmoid_f := 1384;
        ELSIF x = 1504 THEN
            sigmoid_f := 1384;
        ELSIF x = 1505 THEN
            sigmoid_f := 1384;
        ELSIF x = 1506 THEN
            sigmoid_f := 1384;
        ELSIF x = 1507 THEN
            sigmoid_f := 1385;
        ELSIF x = 1508 THEN
            sigmoid_f := 1385;
        ELSIF x = 1509 THEN
            sigmoid_f := 1385;
        ELSIF x = 1510 THEN
            sigmoid_f := 1385;
        ELSIF x = 1511 THEN
            sigmoid_f := 1386;
        ELSIF x = 1512 THEN
            sigmoid_f := 1386;
        ELSIF x = 1513 THEN
            sigmoid_f := 1386;
        ELSIF x = 1514 THEN
            sigmoid_f := 1386;
        ELSIF x = 1515 THEN
            sigmoid_f := 1386;
        ELSIF x = 1516 THEN
            sigmoid_f := 1387;
        ELSIF x = 1517 THEN
            sigmoid_f := 1387;
        ELSIF x = 1518 THEN
            sigmoid_f := 1387;
        ELSIF x = 1519 THEN
            sigmoid_f := 1387;
        ELSIF x = 1520 THEN
            sigmoid_f := 1388;
        ELSIF x = 1521 THEN
            sigmoid_f := 1388;
        ELSIF x = 1522 THEN
            sigmoid_f := 1388;
        ELSIF x = 1523 THEN
            sigmoid_f := 1388;
        ELSIF x = 1524 THEN
            sigmoid_f := 1389;
        ELSIF x = 1525 THEN
            sigmoid_f := 1389;
        ELSIF x = 1526 THEN
            sigmoid_f := 1389;
        ELSIF x = 1527 THEN
            sigmoid_f := 1389;
        ELSIF x = 1528 THEN
            sigmoid_f := 1389;
        ELSIF x = 1529 THEN
            sigmoid_f := 1390;
        ELSIF x = 1530 THEN
            sigmoid_f := 1390;
        ELSIF x = 1531 THEN
            sigmoid_f := 1390;
        ELSIF x = 1532 THEN
            sigmoid_f := 1390;
        ELSIF x = 1533 THEN
            sigmoid_f := 1391;
        ELSIF x = 1534 THEN
            sigmoid_f := 1391;
        ELSIF x = 1535 THEN
            sigmoid_f := 1391;
        ELSIF x = 1536 THEN
            sigmoid_f := 1392;
        ELSIF x = 1537 THEN
            sigmoid_f := 1392;
        ELSIF x = 1538 THEN
            sigmoid_f := 1392;
        ELSIF x = 1539 THEN
            sigmoid_f := 1392;
        ELSIF x = 1540 THEN
            sigmoid_f := 1392;
        ELSIF x = 1541 THEN
            sigmoid_f := 1393;
        ELSIF x = 1542 THEN
            sigmoid_f := 1393;
        ELSIF x = 1543 THEN
            sigmoid_f := 1393;
        ELSIF x = 1544 THEN
            sigmoid_f := 1393;
        ELSIF x = 1545 THEN
            sigmoid_f := 1393;
        ELSIF x = 1546 THEN
            sigmoid_f := 1394;
        ELSIF x = 1547 THEN
            sigmoid_f := 1394;
        ELSIF x = 1548 THEN
            sigmoid_f := 1394;
        ELSIF x = 1549 THEN
            sigmoid_f := 1394;
        ELSIF x = 1550 THEN
            sigmoid_f := 1394;
        ELSIF x = 1551 THEN
            sigmoid_f := 1395;
        ELSIF x = 1552 THEN
            sigmoid_f := 1395;
        ELSIF x = 1553 THEN
            sigmoid_f := 1395;
        ELSIF x = 1554 THEN
            sigmoid_f := 1395;
        ELSIF x = 1555 THEN
            sigmoid_f := 1395;
        ELSIF x = 1556 THEN
            sigmoid_f := 1396;
        ELSIF x = 1557 THEN
            sigmoid_f := 1396;
        ELSIF x = 1558 THEN
            sigmoid_f := 1396;
        ELSIF x = 1559 THEN
            sigmoid_f := 1396;
        ELSIF x = 1560 THEN
            sigmoid_f := 1396;
        ELSIF x = 1561 THEN
            sigmoid_f := 1397;
        ELSIF x = 1562 THEN
            sigmoid_f := 1397;
        ELSIF x = 1563 THEN
            sigmoid_f := 1397;
        ELSIF x = 1564 THEN
            sigmoid_f := 1397;
        ELSIF x = 1565 THEN
            sigmoid_f := 1398;
        ELSIF x = 1566 THEN
            sigmoid_f := 1398;
        ELSIF x = 1567 THEN
            sigmoid_f := 1398;
        ELSIF x = 1568 THEN
            sigmoid_f := 1398;
        ELSIF x = 1569 THEN
            sigmoid_f := 1398;
        ELSIF x = 1570 THEN
            sigmoid_f := 1399;
        ELSIF x = 1571 THEN
            sigmoid_f := 1399;
        ELSIF x = 1572 THEN
            sigmoid_f := 1399;
        ELSIF x = 1573 THEN
            sigmoid_f := 1399;
        ELSIF x = 1574 THEN
            sigmoid_f := 1399;
        ELSIF x = 1575 THEN
            sigmoid_f := 1400;
        ELSIF x = 1576 THEN
            sigmoid_f := 1400;
        ELSIF x = 1577 THEN
            sigmoid_f := 1400;
        ELSIF x = 1578 THEN
            sigmoid_f := 1400;
        ELSIF x = 1579 THEN
            sigmoid_f := 1400;
        ELSIF x = 1580 THEN
            sigmoid_f := 1401;
        ELSIF x = 1581 THEN
            sigmoid_f := 1401;
        ELSIF x = 1582 THEN
            sigmoid_f := 1401;
        ELSIF x = 1583 THEN
            sigmoid_f := 1401;
        ELSIF x = 1584 THEN
            sigmoid_f := 1401;
        ELSIF x = 1585 THEN
            sigmoid_f := 1402;
        ELSIF x = 1586 THEN
            sigmoid_f := 1402;
        ELSIF x = 1587 THEN
            sigmoid_f := 1402;
        ELSIF x = 1588 THEN
            sigmoid_f := 1402;
        ELSIF x = 1589 THEN
            sigmoid_f := 1402;
        ELSIF x = 1590 THEN
            sigmoid_f := 1403;
        ELSIF x = 1591 THEN
            sigmoid_f := 1403;
        ELSIF x = 1592 THEN
            sigmoid_f := 1403;
        ELSIF x = 1593 THEN
            sigmoid_f := 1403;
        ELSIF x = 1594 THEN
            sigmoid_f := 1404;
        ELSIF x = 1595 THEN
            sigmoid_f := 1404;
        ELSIF x = 1596 THEN
            sigmoid_f := 1404;
        ELSIF x = 1597 THEN
            sigmoid_f := 1404;
        ELSIF x = 1598 THEN
            sigmoid_f := 1404;
        ELSIF x = 1599 THEN
            sigmoid_f := 1405;
        ELSIF x = 1600 THEN
            sigmoid_f := 1405;
        ELSIF x = 1601 THEN
            sigmoid_f := 1405;
        ELSIF x = 1602 THEN
            sigmoid_f := 1405;
        ELSIF x = 1603 THEN
            sigmoid_f := 1405;
        ELSIF x = 1604 THEN
            sigmoid_f := 1406;
        ELSIF x = 1605 THEN
            sigmoid_f := 1406;
        ELSIF x = 1606 THEN
            sigmoid_f := 1406;
        ELSIF x = 1607 THEN
            sigmoid_f := 1406;
        ELSIF x = 1608 THEN
            sigmoid_f := 1406;
        ELSIF x = 1609 THEN
            sigmoid_f := 1407;
        ELSIF x = 1610 THEN
            sigmoid_f := 1407;
        ELSIF x = 1611 THEN
            sigmoid_f := 1407;
        ELSIF x = 1612 THEN
            sigmoid_f := 1407;
        ELSIF x = 1613 THEN
            sigmoid_f := 1407;
        ELSIF x = 1614 THEN
            sigmoid_f := 1408;
        ELSIF x = 1615 THEN
            sigmoid_f := 1408;
        ELSIF x = 1616 THEN
            sigmoid_f := 1408;
        ELSIF x = 1617 THEN
            sigmoid_f := 1408;
        ELSIF x = 1618 THEN
            sigmoid_f := 1408;
        ELSIF x = 1619 THEN
            sigmoid_f := 1409;
        ELSIF x = 1620 THEN
            sigmoid_f := 1409;
        ELSIF x = 1621 THEN
            sigmoid_f := 1409;
        ELSIF x = 1622 THEN
            sigmoid_f := 1409;
        ELSIF x = 1623 THEN
            sigmoid_f := 1410;
        ELSIF x = 1624 THEN
            sigmoid_f := 1410;
        ELSIF x = 1625 THEN
            sigmoid_f := 1410;
        ELSIF x = 1626 THEN
            sigmoid_f := 1410;
        ELSIF x = 1627 THEN
            sigmoid_f := 1410;
        ELSIF x = 1628 THEN
            sigmoid_f := 1411;
        ELSIF x = 1629 THEN
            sigmoid_f := 1411;
        ELSIF x = 1630 THEN
            sigmoid_f := 1411;
        ELSIF x = 1631 THEN
            sigmoid_f := 1411;
        ELSIF x = 1632 THEN
            sigmoid_f := 1411;
        ELSIF x = 1633 THEN
            sigmoid_f := 1412;
        ELSIF x = 1634 THEN
            sigmoid_f := 1412;
        ELSIF x = 1635 THEN
            sigmoid_f := 1412;
        ELSIF x = 1636 THEN
            sigmoid_f := 1412;
        ELSIF x = 1637 THEN
            sigmoid_f := 1412;
        ELSIF x = 1638 THEN
            sigmoid_f := 1413;
        ELSIF x = 1639 THEN
            sigmoid_f := 1413;
        ELSIF x = 1640 THEN
            sigmoid_f := 1413;
        ELSIF x = 1641 THEN
            sigmoid_f := 1413;
        ELSIF x = 1642 THEN
            sigmoid_f := 1413;
        ELSIF x = 1643 THEN
            sigmoid_f := 1414;
        ELSIF x = 1644 THEN
            sigmoid_f := 1414;
        ELSIF x = 1645 THEN
            sigmoid_f := 1414;
        ELSIF x = 1646 THEN
            sigmoid_f := 1414;
        ELSIF x = 1647 THEN
            sigmoid_f := 1414;
        ELSIF x = 1648 THEN
            sigmoid_f := 1415;
        ELSIF x = 1649 THEN
            sigmoid_f := 1415;
        ELSIF x = 1650 THEN
            sigmoid_f := 1415;
        ELSIF x = 1651 THEN
            sigmoid_f := 1415;
        ELSIF x = 1652 THEN
            sigmoid_f := 1416;
        ELSIF x = 1653 THEN
            sigmoid_f := 1416;
        ELSIF x = 1654 THEN
            sigmoid_f := 1416;
        ELSIF x = 1655 THEN
            sigmoid_f := 1416;
        ELSIF x = 1656 THEN
            sigmoid_f := 1416;
        ELSIF x = 1657 THEN
            sigmoid_f := 1417;
        ELSIF x = 1658 THEN
            sigmoid_f := 1417;
        ELSIF x = 1659 THEN
            sigmoid_f := 1417;
        ELSIF x = 1660 THEN
            sigmoid_f := 1417;
        ELSIF x = 1661 THEN
            sigmoid_f := 1417;
        ELSIF x = 1662 THEN
            sigmoid_f := 1418;
        ELSIF x = 1663 THEN
            sigmoid_f := 1418;
        ELSIF x = 1664 THEN
            sigmoid_f := 1418;
        ELSIF x = 1665 THEN
            sigmoid_f := 1418;
        ELSIF x = 1666 THEN
            sigmoid_f := 1418;
        ELSIF x = 1667 THEN
            sigmoid_f := 1419;
        ELSIF x = 1668 THEN
            sigmoid_f := 1419;
        ELSIF x = 1669 THEN
            sigmoid_f := 1419;
        ELSIF x = 1670 THEN
            sigmoid_f := 1419;
        ELSIF x = 1671 THEN
            sigmoid_f := 1419;
        ELSIF x = 1672 THEN
            sigmoid_f := 1420;
        ELSIF x = 1673 THEN
            sigmoid_f := 1420;
        ELSIF x = 1674 THEN
            sigmoid_f := 1420;
        ELSIF x = 1675 THEN
            sigmoid_f := 1420;
        ELSIF x = 1676 THEN
            sigmoid_f := 1420;
        ELSIF x = 1677 THEN
            sigmoid_f := 1421;
        ELSIF x = 1678 THEN
            sigmoid_f := 1421;
        ELSIF x = 1679 THEN
            sigmoid_f := 1421;
        ELSIF x = 1680 THEN
            sigmoid_f := 1421;
        ELSIF x = 1681 THEN
            sigmoid_f := 1422;
        ELSIF x = 1682 THEN
            sigmoid_f := 1422;
        ELSIF x = 1683 THEN
            sigmoid_f := 1422;
        ELSIF x = 1684 THEN
            sigmoid_f := 1422;
        ELSIF x = 1685 THEN
            sigmoid_f := 1422;
        ELSIF x = 1686 THEN
            sigmoid_f := 1423;
        ELSIF x = 1687 THEN
            sigmoid_f := 1423;
        ELSIF x = 1688 THEN
            sigmoid_f := 1423;
        ELSIF x = 1689 THEN
            sigmoid_f := 1423;
        ELSIF x = 1690 THEN
            sigmoid_f := 1423;
        ELSIF x = 1691 THEN
            sigmoid_f := 1424;
        ELSIF x = 1692 THEN
            sigmoid_f := 1424;
        ELSIF x = 1693 THEN
            sigmoid_f := 1424;
        ELSIF x = 1694 THEN
            sigmoid_f := 1424;
        ELSIF x = 1695 THEN
            sigmoid_f := 1424;
        ELSIF x = 1696 THEN
            sigmoid_f := 1425;
        ELSIF x = 1697 THEN
            sigmoid_f := 1425;
        ELSIF x = 1698 THEN
            sigmoid_f := 1425;
        ELSIF x = 1699 THEN
            sigmoid_f := 1425;
        ELSIF x = 1700 THEN
            sigmoid_f := 1425;
        ELSIF x = 1701 THEN
            sigmoid_f := 1426;
        ELSIF x = 1702 THEN
            sigmoid_f := 1426;
        ELSIF x = 1703 THEN
            sigmoid_f := 1426;
        ELSIF x = 1704 THEN
            sigmoid_f := 1426;
        ELSIF x = 1705 THEN
            sigmoid_f := 1426;
        ELSIF x = 1706 THEN
            sigmoid_f := 1427;
        ELSIF x = 1707 THEN
            sigmoid_f := 1427;
        ELSIF x = 1708 THEN
            sigmoid_f := 1427;
        ELSIF x = 1709 THEN
            sigmoid_f := 1427;
        ELSIF x = 1710 THEN
            sigmoid_f := 1428;
        ELSIF x = 1711 THEN
            sigmoid_f := 1428;
        ELSIF x = 1712 THEN
            sigmoid_f := 1428;
        ELSIF x = 1713 THEN
            sigmoid_f := 1428;
        ELSIF x = 1714 THEN
            sigmoid_f := 1428;
        ELSIF x = 1715 THEN
            sigmoid_f := 1429;
        ELSIF x = 1716 THEN
            sigmoid_f := 1429;
        ELSIF x = 1717 THEN
            sigmoid_f := 1429;
        ELSIF x = 1718 THEN
            sigmoid_f := 1429;
        ELSIF x = 1719 THEN
            sigmoid_f := 1429;
        ELSIF x = 1720 THEN
            sigmoid_f := 1430;
        ELSIF x = 1721 THEN
            sigmoid_f := 1430;
        ELSIF x = 1722 THEN
            sigmoid_f := 1430;
        ELSIF x = 1723 THEN
            sigmoid_f := 1430;
        ELSIF x = 1724 THEN
            sigmoid_f := 1430;
        ELSIF x = 1725 THEN
            sigmoid_f := 1431;
        ELSIF x = 1726 THEN
            sigmoid_f := 1431;
        ELSIF x = 1727 THEN
            sigmoid_f := 1431;
        ELSIF x = 1728 THEN
            sigmoid_f := 1431;
        ELSIF x = 1729 THEN
            sigmoid_f := 1431;
        ELSIF x = 1730 THEN
            sigmoid_f := 1432;
        ELSIF x = 1731 THEN
            sigmoid_f := 1432;
        ELSIF x = 1732 THEN
            sigmoid_f := 1432;
        ELSIF x = 1733 THEN
            sigmoid_f := 1432;
        ELSIF x = 1734 THEN
            sigmoid_f := 1432;
        ELSIF x = 1735 THEN
            sigmoid_f := 1433;
        ELSIF x = 1736 THEN
            sigmoid_f := 1433;
        ELSIF x = 1737 THEN
            sigmoid_f := 1433;
        ELSIF x = 1738 THEN
            sigmoid_f := 1433;
        ELSIF x = 1739 THEN
            sigmoid_f := 1434;
        ELSIF x = 1740 THEN
            sigmoid_f := 1434;
        ELSIF x = 1741 THEN
            sigmoid_f := 1434;
        ELSIF x = 1742 THEN
            sigmoid_f := 1434;
        ELSIF x = 1743 THEN
            sigmoid_f := 1434;
        ELSIF x = 1744 THEN
            sigmoid_f := 1435;
        ELSIF x = 1745 THEN
            sigmoid_f := 1435;
        ELSIF x = 1746 THEN
            sigmoid_f := 1435;
        ELSIF x = 1747 THEN
            sigmoid_f := 1435;
        ELSIF x = 1748 THEN
            sigmoid_f := 1435;
        ELSIF x = 1749 THEN
            sigmoid_f := 1436;
        ELSIF x = 1750 THEN
            sigmoid_f := 1436;
        ELSIF x = 1751 THEN
            sigmoid_f := 1436;
        ELSIF x = 1752 THEN
            sigmoid_f := 1436;
        ELSIF x = 1753 THEN
            sigmoid_f := 1436;
        ELSIF x = 1754 THEN
            sigmoid_f := 1437;
        ELSIF x = 1755 THEN
            sigmoid_f := 1437;
        ELSIF x = 1756 THEN
            sigmoid_f := 1437;
        ELSIF x = 1757 THEN
            sigmoid_f := 1437;
        ELSIF x = 1758 THEN
            sigmoid_f := 1437;
        ELSIF x = 1759 THEN
            sigmoid_f := 1438;
        ELSIF x = 1760 THEN
            sigmoid_f := 1438;
        ELSIF x = 1761 THEN
            sigmoid_f := 1438;
        ELSIF x = 1762 THEN
            sigmoid_f := 1438;
        ELSIF x = 1763 THEN
            sigmoid_f := 1438;
        ELSIF x = 1764 THEN
            sigmoid_f := 1439;
        ELSIF x = 1765 THEN
            sigmoid_f := 1439;
        ELSIF x = 1766 THEN
            sigmoid_f := 1439;
        ELSIF x = 1767 THEN
            sigmoid_f := 1439;
        ELSIF x = 1768 THEN
            sigmoid_f := 1440;
        ELSIF x = 1769 THEN
            sigmoid_f := 1440;
        ELSIF x = 1770 THEN
            sigmoid_f := 1440;
        ELSIF x = 1771 THEN
            sigmoid_f := 1440;
        ELSIF x = 1772 THEN
            sigmoid_f := 1440;
        ELSIF x = 1773 THEN
            sigmoid_f := 1441;
        ELSIF x = 1774 THEN
            sigmoid_f := 1441;
        ELSIF x = 1775 THEN
            sigmoid_f := 1441;
        ELSIF x = 1776 THEN
            sigmoid_f := 1441;
        ELSIF x = 1777 THEN
            sigmoid_f := 1441;
        ELSIF x = 1778 THEN
            sigmoid_f := 1442;
        ELSIF x = 1779 THEN
            sigmoid_f := 1442;
        ELSIF x = 1780 THEN
            sigmoid_f := 1442;
        ELSIF x = 1781 THEN
            sigmoid_f := 1442;
        ELSIF x = 1782 THEN
            sigmoid_f := 1442;
        ELSIF x = 1783 THEN
            sigmoid_f := 1443;
        ELSIF x = 1784 THEN
            sigmoid_f := 1443;
        ELSIF x = 1785 THEN
            sigmoid_f := 1443;
        ELSIF x = 1786 THEN
            sigmoid_f := 1443;
        ELSIF x = 1787 THEN
            sigmoid_f := 1443;
        ELSIF x = 1788 THEN
            sigmoid_f := 1444;
        ELSIF x = 1789 THEN
            sigmoid_f := 1444;
        ELSIF x = 1790 THEN
            sigmoid_f := 1444;
        ELSIF x = 1791 THEN
            sigmoid_f := 1444;
        ELSIF x = 1792 THEN
            sigmoid_f := 1445;
        ELSIF x = 1793 THEN
            sigmoid_f := 1445;
        ELSIF x = 1794 THEN
            sigmoid_f := 1445;
        ELSIF x = 1795 THEN
            sigmoid_f := 1445;
        ELSIF x = 1796 THEN
            sigmoid_f := 1445;
        ELSIF x = 1797 THEN
            sigmoid_f := 1446;
        ELSIF x = 1798 THEN
            sigmoid_f := 1446;
        ELSIF x = 1799 THEN
            sigmoid_f := 1446;
        ELSIF x = 1800 THEN
            sigmoid_f := 1446;
        ELSIF x = 1801 THEN
            sigmoid_f := 1446;
        ELSIF x = 1802 THEN
            sigmoid_f := 1447;
        ELSIF x = 1803 THEN
            sigmoid_f := 1447;
        ELSIF x = 1804 THEN
            sigmoid_f := 1447;
        ELSIF x = 1805 THEN
            sigmoid_f := 1447;
        ELSIF x = 1806 THEN
            sigmoid_f := 1447;
        ELSIF x = 1807 THEN
            sigmoid_f := 1448;
        ELSIF x = 1808 THEN
            sigmoid_f := 1448;
        ELSIF x = 1809 THEN
            sigmoid_f := 1448;
        ELSIF x = 1810 THEN
            sigmoid_f := 1448;
        ELSIF x = 1811 THEN
            sigmoid_f := 1448;
        ELSIF x = 1812 THEN
            sigmoid_f := 1449;
        ELSIF x = 1813 THEN
            sigmoid_f := 1449;
        ELSIF x = 1814 THEN
            sigmoid_f := 1449;
        ELSIF x = 1815 THEN
            sigmoid_f := 1449;
        ELSIF x = 1816 THEN
            sigmoid_f := 1449;
        ELSIF x = 1817 THEN
            sigmoid_f := 1450;
        ELSIF x = 1818 THEN
            sigmoid_f := 1450;
        ELSIF x = 1819 THEN
            sigmoid_f := 1450;
        ELSIF x = 1820 THEN
            sigmoid_f := 1450;
        ELSIF x = 1821 THEN
            sigmoid_f := 1451;
        ELSIF x = 1822 THEN
            sigmoid_f := 1451;
        ELSIF x = 1823 THEN
            sigmoid_f := 1451;
        ELSIF x = 1824 THEN
            sigmoid_f := 1451;
        ELSIF x = 1825 THEN
            sigmoid_f := 1451;
        ELSIF x = 1826 THEN
            sigmoid_f := 1452;
        ELSIF x = 1827 THEN
            sigmoid_f := 1452;
        ELSIF x = 1828 THEN
            sigmoid_f := 1452;
        ELSIF x = 1829 THEN
            sigmoid_f := 1452;
        ELSIF x = 1830 THEN
            sigmoid_f := 1452;
        ELSIF x = 1831 THEN
            sigmoid_f := 1453;
        ELSIF x = 1832 THEN
            sigmoid_f := 1453;
        ELSIF x = 1833 THEN
            sigmoid_f := 1453;
        ELSIF x = 1834 THEN
            sigmoid_f := 1453;
        ELSIF x = 1835 THEN
            sigmoid_f := 1453;
        ELSIF x = 1836 THEN
            sigmoid_f := 1454;
        ELSIF x = 1837 THEN
            sigmoid_f := 1454;
        ELSIF x = 1838 THEN
            sigmoid_f := 1454;
        ELSIF x = 1839 THEN
            sigmoid_f := 1454;
        ELSIF x = 1840 THEN
            sigmoid_f := 1454;
        ELSIF x = 1841 THEN
            sigmoid_f := 1455;
        ELSIF x = 1842 THEN
            sigmoid_f := 1455;
        ELSIF x = 1843 THEN
            sigmoid_f := 1455;
        ELSIF x = 1844 THEN
            sigmoid_f := 1455;
        ELSIF x = 1845 THEN
            sigmoid_f := 1455;
        ELSIF x = 1846 THEN
            sigmoid_f := 1456;
        ELSIF x = 1847 THEN
            sigmoid_f := 1456;
        ELSIF x = 1848 THEN
            sigmoid_f := 1456;
        ELSIF x = 1849 THEN
            sigmoid_f := 1456;
        ELSIF x = 1850 THEN
            sigmoid_f := 1457;
        ELSIF x = 1851 THEN
            sigmoid_f := 1457;
        ELSIF x = 1852 THEN
            sigmoid_f := 1457;
        ELSIF x = 1853 THEN
            sigmoid_f := 1457;
        ELSIF x = 1854 THEN
            sigmoid_f := 1457;
        ELSIF x = 1855 THEN
            sigmoid_f := 1458;
        ELSIF x = 1856 THEN
            sigmoid_f := 1458;
        ELSIF x = 1857 THEN
            sigmoid_f := 1458;
        ELSIF x = 1858 THEN
            sigmoid_f := 1458;
        ELSIF x = 1859 THEN
            sigmoid_f := 1458;
        ELSIF x = 1860 THEN
            sigmoid_f := 1459;
        ELSIF x = 1861 THEN
            sigmoid_f := 1459;
        ELSIF x = 1862 THEN
            sigmoid_f := 1459;
        ELSIF x = 1863 THEN
            sigmoid_f := 1459;
        ELSIF x = 1864 THEN
            sigmoid_f := 1459;
        ELSIF x = 1865 THEN
            sigmoid_f := 1460;
        ELSIF x = 1866 THEN
            sigmoid_f := 1460;
        ELSIF x = 1867 THEN
            sigmoid_f := 1460;
        ELSIF x = 1868 THEN
            sigmoid_f := 1460;
        ELSIF x = 1869 THEN
            sigmoid_f := 1460;
        ELSIF x = 1870 THEN
            sigmoid_f := 1461;
        ELSIF x = 1871 THEN
            sigmoid_f := 1461;
        ELSIF x = 1872 THEN
            sigmoid_f := 1461;
        ELSIF x = 1873 THEN
            sigmoid_f := 1461;
        ELSIF x = 1874 THEN
            sigmoid_f := 1461;
        ELSIF x = 1875 THEN
            sigmoid_f := 1462;
        ELSIF x = 1876 THEN
            sigmoid_f := 1462;
        ELSIF x = 1877 THEN
            sigmoid_f := 1462;
        ELSIF x = 1878 THEN
            sigmoid_f := 1462;
        ELSIF x = 1879 THEN
            sigmoid_f := 1463;
        ELSIF x = 1880 THEN
            sigmoid_f := 1463;
        ELSIF x = 1881 THEN
            sigmoid_f := 1463;
        ELSIF x = 1882 THEN
            sigmoid_f := 1463;
        ELSIF x = 1883 THEN
            sigmoid_f := 1463;
        ELSIF x = 1884 THEN
            sigmoid_f := 1464;
        ELSIF x = 1885 THEN
            sigmoid_f := 1464;
        ELSIF x = 1886 THEN
            sigmoid_f := 1464;
        ELSIF x = 1887 THEN
            sigmoid_f := 1464;
        ELSIF x = 1888 THEN
            sigmoid_f := 1464;
        ELSIF x = 1889 THEN
            sigmoid_f := 1465;
        ELSIF x = 1890 THEN
            sigmoid_f := 1465;
        ELSIF x = 1891 THEN
            sigmoid_f := 1465;
        ELSIF x = 1892 THEN
            sigmoid_f := 1465;
        ELSIF x = 1893 THEN
            sigmoid_f := 1465;
        ELSIF x = 1894 THEN
            sigmoid_f := 1466;
        ELSIF x = 1895 THEN
            sigmoid_f := 1466;
        ELSIF x = 1896 THEN
            sigmoid_f := 1466;
        ELSIF x = 1897 THEN
            sigmoid_f := 1466;
        ELSIF x = 1898 THEN
            sigmoid_f := 1466;
        ELSIF x = 1899 THEN
            sigmoid_f := 1467;
        ELSIF x = 1900 THEN
            sigmoid_f := 1467;
        ELSIF x = 1901 THEN
            sigmoid_f := 1467;
        ELSIF x = 1902 THEN
            sigmoid_f := 1467;
        ELSIF x = 1903 THEN
            sigmoid_f := 1467;
        ELSIF x = 1904 THEN
            sigmoid_f := 1468;
        ELSIF x = 1905 THEN
            sigmoid_f := 1468;
        ELSIF x = 1906 THEN
            sigmoid_f := 1468;
        ELSIF x = 1907 THEN
            sigmoid_f := 1468;
        ELSIF x = 1908 THEN
            sigmoid_f := 1469;
        ELSIF x = 1909 THEN
            sigmoid_f := 1469;
        ELSIF x = 1910 THEN
            sigmoid_f := 1469;
        ELSIF x = 1911 THEN
            sigmoid_f := 1469;
        ELSIF x = 1912 THEN
            sigmoid_f := 1469;
        ELSIF x = 1913 THEN
            sigmoid_f := 1470;
        ELSIF x = 1914 THEN
            sigmoid_f := 1470;
        ELSIF x = 1915 THEN
            sigmoid_f := 1470;
        ELSIF x = 1916 THEN
            sigmoid_f := 1470;
        ELSIF x = 1917 THEN
            sigmoid_f := 1470;
        ELSIF x = 1918 THEN
            sigmoid_f := 1471;
        ELSIF x = 1919 THEN
            sigmoid_f := 1471;
        ELSIF x = 1920 THEN
            sigmoid_f := 1471;
        ELSIF x = 1921 THEN
            sigmoid_f := 1471;
        ELSIF x = 1922 THEN
            sigmoid_f := 1471;
        ELSIF x = 1923 THEN
            sigmoid_f := 1472;
        ELSIF x = 1924 THEN
            sigmoid_f := 1472;
        ELSIF x = 1925 THEN
            sigmoid_f := 1472;
        ELSIF x = 1926 THEN
            sigmoid_f := 1472;
        ELSIF x = 1927 THEN
            sigmoid_f := 1472;
        ELSIF x = 1928 THEN
            sigmoid_f := 1473;
        ELSIF x = 1929 THEN
            sigmoid_f := 1473;
        ELSIF x = 1930 THEN
            sigmoid_f := 1473;
        ELSIF x = 1931 THEN
            sigmoid_f := 1473;
        ELSIF x = 1932 THEN
            sigmoid_f := 1473;
        ELSIF x = 1933 THEN
            sigmoid_f := 1474;
        ELSIF x = 1934 THEN
            sigmoid_f := 1474;
        ELSIF x = 1935 THEN
            sigmoid_f := 1474;
        ELSIF x = 1936 THEN
            sigmoid_f := 1474;
        ELSIF x = 1937 THEN
            sigmoid_f := 1475;
        ELSIF x = 1938 THEN
            sigmoid_f := 1475;
        ELSIF x = 1939 THEN
            sigmoid_f := 1475;
        ELSIF x = 1940 THEN
            sigmoid_f := 1475;
        ELSIF x = 1941 THEN
            sigmoid_f := 1475;
        ELSIF x = 1942 THEN
            sigmoid_f := 1476;
        ELSIF x = 1943 THEN
            sigmoid_f := 1476;
        ELSIF x = 1944 THEN
            sigmoid_f := 1476;
        ELSIF x = 1945 THEN
            sigmoid_f := 1476;
        ELSIF x = 1946 THEN
            sigmoid_f := 1476;
        ELSIF x = 1947 THEN
            sigmoid_f := 1477;
        ELSIF x = 1948 THEN
            sigmoid_f := 1477;
        ELSIF x = 1949 THEN
            sigmoid_f := 1477;
        ELSIF x = 1950 THEN
            sigmoid_f := 1477;
        ELSIF x = 1951 THEN
            sigmoid_f := 1477;
        ELSIF x = 1952 THEN
            sigmoid_f := 1478;
        ELSIF x = 1953 THEN
            sigmoid_f := 1478;
        ELSIF x = 1954 THEN
            sigmoid_f := 1478;
        ELSIF x = 1955 THEN
            sigmoid_f := 1478;
        ELSIF x = 1956 THEN
            sigmoid_f := 1478;
        ELSIF x = 1957 THEN
            sigmoid_f := 1479;
        ELSIF x = 1958 THEN
            sigmoid_f := 1479;
        ELSIF x = 1959 THEN
            sigmoid_f := 1479;
        ELSIF x = 1960 THEN
            sigmoid_f := 1479;
        ELSIF x = 1961 THEN
            sigmoid_f := 1479;
        ELSIF x = 1962 THEN
            sigmoid_f := 1480;
        ELSIF x = 1963 THEN
            sigmoid_f := 1480;
        ELSIF x = 1964 THEN
            sigmoid_f := 1480;
        ELSIF x = 1965 THEN
            sigmoid_f := 1480;
        ELSIF x = 1966 THEN
            sigmoid_f := 1481;
        ELSIF x = 1967 THEN
            sigmoid_f := 1481;
        ELSIF x = 1968 THEN
            sigmoid_f := 1481;
        ELSIF x = 1969 THEN
            sigmoid_f := 1481;
        ELSIF x = 1970 THEN
            sigmoid_f := 1481;
        ELSIF x = 1971 THEN
            sigmoid_f := 1482;
        ELSIF x = 1972 THEN
            sigmoid_f := 1482;
        ELSIF x = 1973 THEN
            sigmoid_f := 1482;
        ELSIF x = 1974 THEN
            sigmoid_f := 1482;
        ELSIF x = 1975 THEN
            sigmoid_f := 1482;
        ELSIF x = 1976 THEN
            sigmoid_f := 1483;
        ELSIF x = 1977 THEN
            sigmoid_f := 1483;
        ELSIF x = 1978 THEN
            sigmoid_f := 1483;
        ELSIF x = 1979 THEN
            sigmoid_f := 1483;
        ELSIF x = 1980 THEN
            sigmoid_f := 1483;
        ELSIF x = 1981 THEN
            sigmoid_f := 1484;
        ELSIF x = 1982 THEN
            sigmoid_f := 1484;
        ELSIF x = 1983 THEN
            sigmoid_f := 1484;
        ELSIF x = 1984 THEN
            sigmoid_f := 1484;
        ELSIF x = 1985 THEN
            sigmoid_f := 1484;
        ELSIF x = 1986 THEN
            sigmoid_f := 1485;
        ELSIF x = 1987 THEN
            sigmoid_f := 1485;
        ELSIF x = 1988 THEN
            sigmoid_f := 1485;
        ELSIF x = 1989 THEN
            sigmoid_f := 1485;
        ELSIF x = 1990 THEN
            sigmoid_f := 1485;
        ELSIF x = 1991 THEN
            sigmoid_f := 1486;
        ELSIF x = 1992 THEN
            sigmoid_f := 1486;
        ELSIF x = 1993 THEN
            sigmoid_f := 1486;
        ELSIF x = 1994 THEN
            sigmoid_f := 1486;
        ELSIF x = 1995 THEN
            sigmoid_f := 1487;
        ELSIF x = 1996 THEN
            sigmoid_f := 1487;
        ELSIF x = 1997 THEN
            sigmoid_f := 1487;
        ELSIF x = 1998 THEN
            sigmoid_f := 1487;
        ELSIF x = 1999 THEN
            sigmoid_f := 1487;
        ELSIF x = 2000 THEN
            sigmoid_f := 1488;
        ELSIF x = 2001 THEN
            sigmoid_f := 1488;
        ELSIF x = 2002 THEN
            sigmoid_f := 1488;
        ELSIF x = 2003 THEN
            sigmoid_f := 1488;
        ELSIF x = 2004 THEN
            sigmoid_f := 1488;
        ELSIF x = 2005 THEN
            sigmoid_f := 1489;
        ELSIF x = 2006 THEN
            sigmoid_f := 1489;
        ELSIF x = 2007 THEN
            sigmoid_f := 1489;
        ELSIF x = 2008 THEN
            sigmoid_f := 1489;
        ELSIF x = 2009 THEN
            sigmoid_f := 1489;
        ELSIF x = 2010 THEN
            sigmoid_f := 1490;
        ELSIF x = 2011 THEN
            sigmoid_f := 1490;
        ELSIF x = 2012 THEN
            sigmoid_f := 1490;
        ELSIF x = 2013 THEN
            sigmoid_f := 1490;
        ELSIF x = 2014 THEN
            sigmoid_f := 1490;
        ELSIF x = 2015 THEN
            sigmoid_f := 1491;
        ELSIF x = 2016 THEN
            sigmoid_f := 1491;
        ELSIF x = 2017 THEN
            sigmoid_f := 1491;
        ELSIF x = 2018 THEN
            sigmoid_f := 1491;
        ELSIF x = 2019 THEN
            sigmoid_f := 1491;
        ELSIF x = 2020 THEN
            sigmoid_f := 1492;
        ELSIF x = 2021 THEN
            sigmoid_f := 1492;
        ELSIF x = 2022 THEN
            sigmoid_f := 1492;
        ELSIF x = 2023 THEN
            sigmoid_f := 1492;
        ELSIF x = 2024 THEN
            sigmoid_f := 1493;
        ELSIF x = 2025 THEN
            sigmoid_f := 1493;
        ELSIF x = 2026 THEN
            sigmoid_f := 1493;
        ELSIF x = 2027 THEN
            sigmoid_f := 1493;
        ELSIF x = 2028 THEN
            sigmoid_f := 1493;
        ELSIF x = 2029 THEN
            sigmoid_f := 1494;
        ELSIF x = 2030 THEN
            sigmoid_f := 1494;
        ELSIF x = 2031 THEN
            sigmoid_f := 1494;
        ELSIF x = 2032 THEN
            sigmoid_f := 1494;
        ELSIF x = 2033 THEN
            sigmoid_f := 1494;
        ELSIF x = 2034 THEN
            sigmoid_f := 1495;
        ELSIF x = 2035 THEN
            sigmoid_f := 1495;
        ELSIF x = 2036 THEN
            sigmoid_f := 1495;
        ELSIF x = 2037 THEN
            sigmoid_f := 1495;
        ELSIF x = 2038 THEN
            sigmoid_f := 1495;
        ELSIF x = 2039 THEN
            sigmoid_f := 1496;
        ELSIF x = 2040 THEN
            sigmoid_f := 1496;
        ELSIF x = 2041 THEN
            sigmoid_f := 1496;
        ELSIF x = 2042 THEN
            sigmoid_f := 1496;
        ELSIF x = 2043 THEN
            sigmoid_f := 1496;
        ELSIF x = 2044 THEN
            sigmoid_f := 1497;
        ELSIF x = 2045 THEN
            sigmoid_f := 1497;
        ELSIF x = 2046 THEN
            sigmoid_f := 1497;
        ELSIF x = 2047 THEN
            sigmoid_f := 1497;
        ELSIF x = 2048 THEN
            sigmoid_f := 1498;
        ELSIF x = 2049 THEN
            sigmoid_f := 1498;
        ELSIF x = 2050 THEN
            sigmoid_f := 1498;
        ELSIF x = 2051 THEN
            sigmoid_f := 1498;
        ELSIF x = 2052 THEN
            sigmoid_f := 1498;
        ELSIF x = 2053 THEN
            sigmoid_f := 1498;
        ELSIF x = 2054 THEN
            sigmoid_f := 1499;
        ELSIF x = 2055 THEN
            sigmoid_f := 1499;
        ELSIF x = 2056 THEN
            sigmoid_f := 1499;
        ELSIF x = 2057 THEN
            sigmoid_f := 1499;
        ELSIF x = 2058 THEN
            sigmoid_f := 1499;
        ELSIF x = 2059 THEN
            sigmoid_f := 1500;
        ELSIF x = 2060 THEN
            sigmoid_f := 1500;
        ELSIF x = 2061 THEN
            sigmoid_f := 1500;
        ELSIF x = 2062 THEN
            sigmoid_f := 1500;
        ELSIF x = 2063 THEN
            sigmoid_f := 1500;
        ELSIF x = 2064 THEN
            sigmoid_f := 1500;
        ELSIF x = 2065 THEN
            sigmoid_f := 1501;
        ELSIF x = 2066 THEN
            sigmoid_f := 1501;
        ELSIF x = 2067 THEN
            sigmoid_f := 1501;
        ELSIF x = 2068 THEN
            sigmoid_f := 1501;
        ELSIF x = 2069 THEN
            sigmoid_f := 1501;
        ELSIF x = 2070 THEN
            sigmoid_f := 1502;
        ELSIF x = 2071 THEN
            sigmoid_f := 1502;
        ELSIF x = 2072 THEN
            sigmoid_f := 1502;
        ELSIF x = 2073 THEN
            sigmoid_f := 1502;
        ELSIF x = 2074 THEN
            sigmoid_f := 1502;
        ELSIF x = 2075 THEN
            sigmoid_f := 1503;
        ELSIF x = 2076 THEN
            sigmoid_f := 1503;
        ELSIF x = 2077 THEN
            sigmoid_f := 1503;
        ELSIF x = 2078 THEN
            sigmoid_f := 1503;
        ELSIF x = 2079 THEN
            sigmoid_f := 1503;
        ELSIF x = 2080 THEN
            sigmoid_f := 1503;
        ELSIF x = 2081 THEN
            sigmoid_f := 1504;
        ELSIF x = 2082 THEN
            sigmoid_f := 1504;
        ELSIF x = 2083 THEN
            sigmoid_f := 1504;
        ELSIF x = 2084 THEN
            sigmoid_f := 1504;
        ELSIF x = 2085 THEN
            sigmoid_f := 1504;
        ELSIF x = 2086 THEN
            sigmoid_f := 1505;
        ELSIF x = 2087 THEN
            sigmoid_f := 1505;
        ELSIF x = 2088 THEN
            sigmoid_f := 1505;
        ELSIF x = 2089 THEN
            sigmoid_f := 1505;
        ELSIF x = 2090 THEN
            sigmoid_f := 1505;
        ELSIF x = 2091 THEN
            sigmoid_f := 1505;
        ELSIF x = 2092 THEN
            sigmoid_f := 1506;
        ELSIF x = 2093 THEN
            sigmoid_f := 1506;
        ELSIF x = 2094 THEN
            sigmoid_f := 1506;
        ELSIF x = 2095 THEN
            sigmoid_f := 1506;
        ELSIF x = 2096 THEN
            sigmoid_f := 1506;
        ELSIF x = 2097 THEN
            sigmoid_f := 1507;
        ELSIF x = 2098 THEN
            sigmoid_f := 1507;
        ELSIF x = 2099 THEN
            sigmoid_f := 1507;
        ELSIF x = 2100 THEN
            sigmoid_f := 1507;
        ELSIF x = 2101 THEN
            sigmoid_f := 1507;
        ELSIF x = 2102 THEN
            sigmoid_f := 1508;
        ELSIF x = 2103 THEN
            sigmoid_f := 1508;
        ELSIF x = 2104 THEN
            sigmoid_f := 1508;
        ELSIF x = 2105 THEN
            sigmoid_f := 1508;
        ELSIF x = 2106 THEN
            sigmoid_f := 1508;
        ELSIF x = 2107 THEN
            sigmoid_f := 1508;
        ELSIF x = 2108 THEN
            sigmoid_f := 1509;
        ELSIF x = 2109 THEN
            sigmoid_f := 1509;
        ELSIF x = 2110 THEN
            sigmoid_f := 1509;
        ELSIF x = 2111 THEN
            sigmoid_f := 1509;
        ELSIF x = 2112 THEN
            sigmoid_f := 1509;
        ELSIF x = 2113 THEN
            sigmoid_f := 1510;
        ELSIF x = 2114 THEN
            sigmoid_f := 1510;
        ELSIF x = 2115 THEN
            sigmoid_f := 1510;
        ELSIF x = 2116 THEN
            sigmoid_f := 1510;
        ELSIF x = 2117 THEN
            sigmoid_f := 1510;
        ELSIF x = 2118 THEN
            sigmoid_f := 1511;
        ELSIF x = 2119 THEN
            sigmoid_f := 1511;
        ELSIF x = 2120 THEN
            sigmoid_f := 1511;
        ELSIF x = 2121 THEN
            sigmoid_f := 1511;
        ELSIF x = 2122 THEN
            sigmoid_f := 1511;
        ELSIF x = 2123 THEN
            sigmoid_f := 1511;
        ELSIF x = 2124 THEN
            sigmoid_f := 1512;
        ELSIF x = 2125 THEN
            sigmoid_f := 1512;
        ELSIF x = 2126 THEN
            sigmoid_f := 1512;
        ELSIF x = 2127 THEN
            sigmoid_f := 1512;
        ELSIF x = 2128 THEN
            sigmoid_f := 1512;
        ELSIF x = 2129 THEN
            sigmoid_f := 1513;
        ELSIF x = 2130 THEN
            sigmoid_f := 1513;
        ELSIF x = 2131 THEN
            sigmoid_f := 1513;
        ELSIF x = 2132 THEN
            sigmoid_f := 1513;
        ELSIF x = 2133 THEN
            sigmoid_f := 1513;
        ELSIF x = 2134 THEN
            sigmoid_f := 1513;
        ELSIF x = 2135 THEN
            sigmoid_f := 1514;
        ELSIF x = 2136 THEN
            sigmoid_f := 1514;
        ELSIF x = 2137 THEN
            sigmoid_f := 1514;
        ELSIF x = 2138 THEN
            sigmoid_f := 1514;
        ELSIF x = 2139 THEN
            sigmoid_f := 1514;
        ELSIF x = 2140 THEN
            sigmoid_f := 1515;
        ELSIF x = 2141 THEN
            sigmoid_f := 1515;
        ELSIF x = 2142 THEN
            sigmoid_f := 1515;
        ELSIF x = 2143 THEN
            sigmoid_f := 1515;
        ELSIF x = 2144 THEN
            sigmoid_f := 1515;
        ELSIF x = 2145 THEN
            sigmoid_f := 1516;
        ELSIF x = 2146 THEN
            sigmoid_f := 1516;
        ELSIF x = 2147 THEN
            sigmoid_f := 1516;
        ELSIF x = 2148 THEN
            sigmoid_f := 1516;
        ELSIF x = 2149 THEN
            sigmoid_f := 1516;
        ELSIF x = 2150 THEN
            sigmoid_f := 1516;
        ELSIF x = 2151 THEN
            sigmoid_f := 1517;
        ELSIF x = 2152 THEN
            sigmoid_f := 1517;
        ELSIF x = 2153 THEN
            sigmoid_f := 1517;
        ELSIF x = 2154 THEN
            sigmoid_f := 1517;
        ELSIF x = 2155 THEN
            sigmoid_f := 1517;
        ELSIF x = 2156 THEN
            sigmoid_f := 1518;
        ELSIF x = 2157 THEN
            sigmoid_f := 1518;
        ELSIF x = 2158 THEN
            sigmoid_f := 1518;
        ELSIF x = 2159 THEN
            sigmoid_f := 1518;
        ELSIF x = 2160 THEN
            sigmoid_f := 1518;
        ELSIF x = 2161 THEN
            sigmoid_f := 1519;
        ELSIF x = 2162 THEN
            sigmoid_f := 1519;
        ELSIF x = 2163 THEN
            sigmoid_f := 1519;
        ELSIF x = 2164 THEN
            sigmoid_f := 1519;
        ELSIF x = 2165 THEN
            sigmoid_f := 1519;
        ELSIF x = 2166 THEN
            sigmoid_f := 1519;
        ELSIF x = 2167 THEN
            sigmoid_f := 1520;
        ELSIF x = 2168 THEN
            sigmoid_f := 1520;
        ELSIF x = 2169 THEN
            sigmoid_f := 1520;
        ELSIF x = 2170 THEN
            sigmoid_f := 1520;
        ELSIF x = 2171 THEN
            sigmoid_f := 1520;
        ELSIF x = 2172 THEN
            sigmoid_f := 1521;
        ELSIF x = 2173 THEN
            sigmoid_f := 1521;
        ELSIF x = 2174 THEN
            sigmoid_f := 1521;
        ELSIF x = 2175 THEN
            sigmoid_f := 1521;
        ELSIF x = 2176 THEN
            sigmoid_f := 1521;
        ELSIF x = 2177 THEN
            sigmoid_f := 1521;
        ELSIF x = 2178 THEN
            sigmoid_f := 1522;
        ELSIF x = 2179 THEN
            sigmoid_f := 1522;
        ELSIF x = 2180 THEN
            sigmoid_f := 1522;
        ELSIF x = 2181 THEN
            sigmoid_f := 1522;
        ELSIF x = 2182 THEN
            sigmoid_f := 1522;
        ELSIF x = 2183 THEN
            sigmoid_f := 1523;
        ELSIF x = 2184 THEN
            sigmoid_f := 1523;
        ELSIF x = 2185 THEN
            sigmoid_f := 1523;
        ELSIF x = 2186 THEN
            sigmoid_f := 1523;
        ELSIF x = 2187 THEN
            sigmoid_f := 1523;
        ELSIF x = 2188 THEN
            sigmoid_f := 1524;
        ELSIF x = 2189 THEN
            sigmoid_f := 1524;
        ELSIF x = 2190 THEN
            sigmoid_f := 1524;
        ELSIF x = 2191 THEN
            sigmoid_f := 1524;
        ELSIF x = 2192 THEN
            sigmoid_f := 1524;
        ELSIF x = 2193 THEN
            sigmoid_f := 1524;
        ELSIF x = 2194 THEN
            sigmoid_f := 1525;
        ELSIF x = 2195 THEN
            sigmoid_f := 1525;
        ELSIF x = 2196 THEN
            sigmoid_f := 1525;
        ELSIF x = 2197 THEN
            sigmoid_f := 1525;
        ELSIF x = 2198 THEN
            sigmoid_f := 1525;
        ELSIF x = 2199 THEN
            sigmoid_f := 1526;
        ELSIF x = 2200 THEN
            sigmoid_f := 1526;
        ELSIF x = 2201 THEN
            sigmoid_f := 1526;
        ELSIF x = 2202 THEN
            sigmoid_f := 1526;
        ELSIF x = 2203 THEN
            sigmoid_f := 1526;
        ELSIF x = 2204 THEN
            sigmoid_f := 1527;
        ELSIF x = 2205 THEN
            sigmoid_f := 1527;
        ELSIF x = 2206 THEN
            sigmoid_f := 1527;
        ELSIF x = 2207 THEN
            sigmoid_f := 1527;
        ELSIF x = 2208 THEN
            sigmoid_f := 1527;
        ELSIF x = 2209 THEN
            sigmoid_f := 1527;
        ELSIF x = 2210 THEN
            sigmoid_f := 1528;
        ELSIF x = 2211 THEN
            sigmoid_f := 1528;
        ELSIF x = 2212 THEN
            sigmoid_f := 1528;
        ELSIF x = 2213 THEN
            sigmoid_f := 1528;
        ELSIF x = 2214 THEN
            sigmoid_f := 1528;
        ELSIF x = 2215 THEN
            sigmoid_f := 1529;
        ELSIF x = 2216 THEN
            sigmoid_f := 1529;
        ELSIF x = 2217 THEN
            sigmoid_f := 1529;
        ELSIF x = 2218 THEN
            sigmoid_f := 1529;
        ELSIF x = 2219 THEN
            sigmoid_f := 1529;
        ELSIF x = 2220 THEN
            sigmoid_f := 1529;
        ELSIF x = 2221 THEN
            sigmoid_f := 1530;
        ELSIF x = 2222 THEN
            sigmoid_f := 1530;
        ELSIF x = 2223 THEN
            sigmoid_f := 1530;
        ELSIF x = 2224 THEN
            sigmoid_f := 1530;
        ELSIF x = 2225 THEN
            sigmoid_f := 1530;
        ELSIF x = 2226 THEN
            sigmoid_f := 1531;
        ELSIF x = 2227 THEN
            sigmoid_f := 1531;
        ELSIF x = 2228 THEN
            sigmoid_f := 1531;
        ELSIF x = 2229 THEN
            sigmoid_f := 1531;
        ELSIF x = 2230 THEN
            sigmoid_f := 1531;
        ELSIF x = 2231 THEN
            sigmoid_f := 1532;
        ELSIF x = 2232 THEN
            sigmoid_f := 1532;
        ELSIF x = 2233 THEN
            sigmoid_f := 1532;
        ELSIF x = 2234 THEN
            sigmoid_f := 1532;
        ELSIF x = 2235 THEN
            sigmoid_f := 1532;
        ELSIF x = 2236 THEN
            sigmoid_f := 1532;
        ELSIF x = 2237 THEN
            sigmoid_f := 1533;
        ELSIF x = 2238 THEN
            sigmoid_f := 1533;
        ELSIF x = 2239 THEN
            sigmoid_f := 1533;
        ELSIF x = 2240 THEN
            sigmoid_f := 1533;
        ELSIF x = 2241 THEN
            sigmoid_f := 1533;
        ELSIF x = 2242 THEN
            sigmoid_f := 1534;
        ELSIF x = 2243 THEN
            sigmoid_f := 1534;
        ELSIF x = 2244 THEN
            sigmoid_f := 1534;
        ELSIF x = 2245 THEN
            sigmoid_f := 1534;
        ELSIF x = 2246 THEN
            sigmoid_f := 1534;
        ELSIF x = 2247 THEN
            sigmoid_f := 1535;
        ELSIF x = 2248 THEN
            sigmoid_f := 1535;
        ELSIF x = 2249 THEN
            sigmoid_f := 1535;
        ELSIF x = 2250 THEN
            sigmoid_f := 1535;
        ELSIF x = 2251 THEN
            sigmoid_f := 1535;
        ELSIF x = 2252 THEN
            sigmoid_f := 1535;
        ELSIF x = 2253 THEN
            sigmoid_f := 1536;
        ELSIF x = 2254 THEN
            sigmoid_f := 1536;
        ELSIF x = 2255 THEN
            sigmoid_f := 1536;
        ELSIF x = 2256 THEN
            sigmoid_f := 1536;
        ELSIF x = 2257 THEN
            sigmoid_f := 1536;
        ELSIF x = 2258 THEN
            sigmoid_f := 1537;
        ELSIF x = 2259 THEN
            sigmoid_f := 1537;
        ELSIF x = 2260 THEN
            sigmoid_f := 1537;
        ELSIF x = 2261 THEN
            sigmoid_f := 1537;
        ELSIF x = 2262 THEN
            sigmoid_f := 1537;
        ELSIF x = 2263 THEN
            sigmoid_f := 1537;
        ELSIF x = 2264 THEN
            sigmoid_f := 1538;
        ELSIF x = 2265 THEN
            sigmoid_f := 1538;
        ELSIF x = 2266 THEN
            sigmoid_f := 1538;
        ELSIF x = 2267 THEN
            sigmoid_f := 1538;
        ELSIF x = 2268 THEN
            sigmoid_f := 1538;
        ELSIF x = 2269 THEN
            sigmoid_f := 1539;
        ELSIF x = 2270 THEN
            sigmoid_f := 1539;
        ELSIF x = 2271 THEN
            sigmoid_f := 1539;
        ELSIF x = 2272 THEN
            sigmoid_f := 1539;
        ELSIF x = 2273 THEN
            sigmoid_f := 1539;
        ELSIF x = 2274 THEN
            sigmoid_f := 1540;
        ELSIF x = 2275 THEN
            sigmoid_f := 1540;
        ELSIF x = 2276 THEN
            sigmoid_f := 1540;
        ELSIF x = 2277 THEN
            sigmoid_f := 1540;
        ELSIF x = 2278 THEN
            sigmoid_f := 1540;
        ELSIF x = 2279 THEN
            sigmoid_f := 1540;
        ELSIF x = 2280 THEN
            sigmoid_f := 1541;
        ELSIF x = 2281 THEN
            sigmoid_f := 1541;
        ELSIF x = 2282 THEN
            sigmoid_f := 1541;
        ELSIF x = 2283 THEN
            sigmoid_f := 1541;
        ELSIF x = 2284 THEN
            sigmoid_f := 1541;
        ELSIF x = 2285 THEN
            sigmoid_f := 1542;
        ELSIF x = 2286 THEN
            sigmoid_f := 1542;
        ELSIF x = 2287 THEN
            sigmoid_f := 1542;
        ELSIF x = 2288 THEN
            sigmoid_f := 1542;
        ELSIF x = 2289 THEN
            sigmoid_f := 1542;
        ELSIF x = 2290 THEN
            sigmoid_f := 1543;
        ELSIF x = 2291 THEN
            sigmoid_f := 1543;
        ELSIF x = 2292 THEN
            sigmoid_f := 1543;
        ELSIF x = 2293 THEN
            sigmoid_f := 1543;
        ELSIF x = 2294 THEN
            sigmoid_f := 1543;
        ELSIF x = 2295 THEN
            sigmoid_f := 1543;
        ELSIF x = 2296 THEN
            sigmoid_f := 1544;
        ELSIF x = 2297 THEN
            sigmoid_f := 1544;
        ELSIF x = 2298 THEN
            sigmoid_f := 1544;
        ELSIF x = 2299 THEN
            sigmoid_f := 1544;
        ELSIF x = 2300 THEN
            sigmoid_f := 1544;
        ELSIF x = 2301 THEN
            sigmoid_f := 1545;
        ELSIF x = 2302 THEN
            sigmoid_f := 1545;
        ELSIF x = 2303 THEN
            sigmoid_f := 1545;
        ELSIF x = 2304 THEN
            sigmoid_f := 1545;
        ELSIF x = 2305 THEN
            sigmoid_f := 1545;
        ELSIF x = 2306 THEN
            sigmoid_f := 1545;
        ELSIF x = 2307 THEN
            sigmoid_f := 1546;
        ELSIF x = 2308 THEN
            sigmoid_f := 1546;
        ELSIF x = 2309 THEN
            sigmoid_f := 1546;
        ELSIF x = 2310 THEN
            sigmoid_f := 1546;
        ELSIF x = 2311 THEN
            sigmoid_f := 1546;
        ELSIF x = 2312 THEN
            sigmoid_f := 1547;
        ELSIF x = 2313 THEN
            sigmoid_f := 1547;
        ELSIF x = 2314 THEN
            sigmoid_f := 1547;
        ELSIF x = 2315 THEN
            sigmoid_f := 1547;
        ELSIF x = 2316 THEN
            sigmoid_f := 1547;
        ELSIF x = 2317 THEN
            sigmoid_f := 1548;
        ELSIF x = 2318 THEN
            sigmoid_f := 1548;
        ELSIF x = 2319 THEN
            sigmoid_f := 1548;
        ELSIF x = 2320 THEN
            sigmoid_f := 1548;
        ELSIF x = 2321 THEN
            sigmoid_f := 1548;
        ELSIF x = 2322 THEN
            sigmoid_f := 1548;
        ELSIF x = 2323 THEN
            sigmoid_f := 1549;
        ELSIF x = 2324 THEN
            sigmoid_f := 1549;
        ELSIF x = 2325 THEN
            sigmoid_f := 1549;
        ELSIF x = 2326 THEN
            sigmoid_f := 1549;
        ELSIF x = 2327 THEN
            sigmoid_f := 1549;
        ELSIF x = 2328 THEN
            sigmoid_f := 1550;
        ELSIF x = 2329 THEN
            sigmoid_f := 1550;
        ELSIF x = 2330 THEN
            sigmoid_f := 1550;
        ELSIF x = 2331 THEN
            sigmoid_f := 1550;
        ELSIF x = 2332 THEN
            sigmoid_f := 1550;
        ELSIF x = 2333 THEN
            sigmoid_f := 1551;
        ELSIF x = 2334 THEN
            sigmoid_f := 1551;
        ELSIF x = 2335 THEN
            sigmoid_f := 1551;
        ELSIF x = 2336 THEN
            sigmoid_f := 1551;
        ELSIF x = 2337 THEN
            sigmoid_f := 1551;
        ELSIF x = 2338 THEN
            sigmoid_f := 1551;
        ELSIF x = 2339 THEN
            sigmoid_f := 1552;
        ELSIF x = 2340 THEN
            sigmoid_f := 1552;
        ELSIF x = 2341 THEN
            sigmoid_f := 1552;
        ELSIF x = 2342 THEN
            sigmoid_f := 1552;
        ELSIF x = 2343 THEN
            sigmoid_f := 1552;
        ELSIF x = 2344 THEN
            sigmoid_f := 1553;
        ELSIF x = 2345 THEN
            sigmoid_f := 1553;
        ELSIF x = 2346 THEN
            sigmoid_f := 1553;
        ELSIF x = 2347 THEN
            sigmoid_f := 1553;
        ELSIF x = 2348 THEN
            sigmoid_f := 1553;
        ELSIF x = 2349 THEN
            sigmoid_f := 1553;
        ELSIF x = 2350 THEN
            sigmoid_f := 1554;
        ELSIF x = 2351 THEN
            sigmoid_f := 1554;
        ELSIF x = 2352 THEN
            sigmoid_f := 1554;
        ELSIF x = 2353 THEN
            sigmoid_f := 1554;
        ELSIF x = 2354 THEN
            sigmoid_f := 1554;
        ELSIF x = 2355 THEN
            sigmoid_f := 1555;
        ELSIF x = 2356 THEN
            sigmoid_f := 1555;
        ELSIF x = 2357 THEN
            sigmoid_f := 1555;
        ELSIF x = 2358 THEN
            sigmoid_f := 1555;
        ELSIF x = 2359 THEN
            sigmoid_f := 1555;
        ELSIF x = 2360 THEN
            sigmoid_f := 1556;
        ELSIF x = 2361 THEN
            sigmoid_f := 1556;
        ELSIF x = 2362 THEN
            sigmoid_f := 1556;
        ELSIF x = 2363 THEN
            sigmoid_f := 1556;
        ELSIF x = 2364 THEN
            sigmoid_f := 1556;
        ELSIF x = 2365 THEN
            sigmoid_f := 1556;
        ELSIF x = 2366 THEN
            sigmoid_f := 1557;
        ELSIF x = 2367 THEN
            sigmoid_f := 1557;
        ELSIF x = 2368 THEN
            sigmoid_f := 1557;
        ELSIF x = 2369 THEN
            sigmoid_f := 1557;
        ELSIF x = 2370 THEN
            sigmoid_f := 1557;
        ELSIF x = 2371 THEN
            sigmoid_f := 1558;
        ELSIF x = 2372 THEN
            sigmoid_f := 1558;
        ELSIF x = 2373 THEN
            sigmoid_f := 1558;
        ELSIF x = 2374 THEN
            sigmoid_f := 1558;
        ELSIF x = 2375 THEN
            sigmoid_f := 1558;
        ELSIF x = 2376 THEN
            sigmoid_f := 1559;
        ELSIF x = 2377 THEN
            sigmoid_f := 1559;
        ELSIF x = 2378 THEN
            sigmoid_f := 1559;
        ELSIF x = 2379 THEN
            sigmoid_f := 1559;
        ELSIF x = 2380 THEN
            sigmoid_f := 1559;
        ELSIF x = 2381 THEN
            sigmoid_f := 1559;
        ELSIF x = 2382 THEN
            sigmoid_f := 1560;
        ELSIF x = 2383 THEN
            sigmoid_f := 1560;
        ELSIF x = 2384 THEN
            sigmoid_f := 1560;
        ELSIF x = 2385 THEN
            sigmoid_f := 1560;
        ELSIF x = 2386 THEN
            sigmoid_f := 1560;
        ELSIF x = 2387 THEN
            sigmoid_f := 1561;
        ELSIF x = 2388 THEN
            sigmoid_f := 1561;
        ELSIF x = 2389 THEN
            sigmoid_f := 1561;
        ELSIF x = 2390 THEN
            sigmoid_f := 1561;
        ELSIF x = 2391 THEN
            sigmoid_f := 1561;
        ELSIF x = 2392 THEN
            sigmoid_f := 1561;
        ELSIF x = 2393 THEN
            sigmoid_f := 1562;
        ELSIF x = 2394 THEN
            sigmoid_f := 1562;
        ELSIF x = 2395 THEN
            sigmoid_f := 1562;
        ELSIF x = 2396 THEN
            sigmoid_f := 1562;
        ELSIF x = 2397 THEN
            sigmoid_f := 1562;
        ELSIF x = 2398 THEN
            sigmoid_f := 1563;
        ELSIF x = 2399 THEN
            sigmoid_f := 1563;
        ELSIF x = 2400 THEN
            sigmoid_f := 1563;
        ELSIF x = 2401 THEN
            sigmoid_f := 1563;
        ELSIF x = 2402 THEN
            sigmoid_f := 1563;
        ELSIF x = 2403 THEN
            sigmoid_f := 1564;
        ELSIF x = 2404 THEN
            sigmoid_f := 1564;
        ELSIF x = 2405 THEN
            sigmoid_f := 1564;
        ELSIF x = 2406 THEN
            sigmoid_f := 1564;
        ELSIF x = 2407 THEN
            sigmoid_f := 1564;
        ELSIF x = 2408 THEN
            sigmoid_f := 1564;
        ELSIF x = 2409 THEN
            sigmoid_f := 1565;
        ELSIF x = 2410 THEN
            sigmoid_f := 1565;
        ELSIF x = 2411 THEN
            sigmoid_f := 1565;
        ELSIF x = 2412 THEN
            sigmoid_f := 1565;
        ELSIF x = 2413 THEN
            sigmoid_f := 1565;
        ELSIF x = 2414 THEN
            sigmoid_f := 1566;
        ELSIF x = 2415 THEN
            sigmoid_f := 1566;
        ELSIF x = 2416 THEN
            sigmoid_f := 1566;
        ELSIF x = 2417 THEN
            sigmoid_f := 1566;
        ELSIF x = 2418 THEN
            sigmoid_f := 1566;
        ELSIF x = 2419 THEN
            sigmoid_f := 1567;
        ELSIF x = 2420 THEN
            sigmoid_f := 1567;
        ELSIF x = 2421 THEN
            sigmoid_f := 1567;
        ELSIF x = 2422 THEN
            sigmoid_f := 1567;
        ELSIF x = 2423 THEN
            sigmoid_f := 1567;
        ELSIF x = 2424 THEN
            sigmoid_f := 1567;
        ELSIF x = 2425 THEN
            sigmoid_f := 1568;
        ELSIF x = 2426 THEN
            sigmoid_f := 1568;
        ELSIF x = 2427 THEN
            sigmoid_f := 1568;
        ELSIF x = 2428 THEN
            sigmoid_f := 1568;
        ELSIF x = 2429 THEN
            sigmoid_f := 1568;
        ELSIF x = 2430 THEN
            sigmoid_f := 1569;
        ELSIF x = 2431 THEN
            sigmoid_f := 1569;
        ELSIF x = 2432 THEN
            sigmoid_f := 1569;
        ELSIF x = 2433 THEN
            sigmoid_f := 1569;
        ELSIF x = 2434 THEN
            sigmoid_f := 1569;
        ELSIF x = 2435 THEN
            sigmoid_f := 1569;
        ELSIF x = 2436 THEN
            sigmoid_f := 1570;
        ELSIF x = 2437 THEN
            sigmoid_f := 1570;
        ELSIF x = 2438 THEN
            sigmoid_f := 1570;
        ELSIF x = 2439 THEN
            sigmoid_f := 1570;
        ELSIF x = 2440 THEN
            sigmoid_f := 1570;
        ELSIF x = 2441 THEN
            sigmoid_f := 1571;
        ELSIF x = 2442 THEN
            sigmoid_f := 1571;
        ELSIF x = 2443 THEN
            sigmoid_f := 1571;
        ELSIF x = 2444 THEN
            sigmoid_f := 1571;
        ELSIF x = 2445 THEN
            sigmoid_f := 1571;
        ELSIF x = 2446 THEN
            sigmoid_f := 1572;
        ELSIF x = 2447 THEN
            sigmoid_f := 1572;
        ELSIF x = 2448 THEN
            sigmoid_f := 1572;
        ELSIF x = 2449 THEN
            sigmoid_f := 1572;
        ELSIF x = 2450 THEN
            sigmoid_f := 1572;
        ELSIF x = 2451 THEN
            sigmoid_f := 1572;
        ELSIF x = 2452 THEN
            sigmoid_f := 1573;
        ELSIF x = 2453 THEN
            sigmoid_f := 1573;
        ELSIF x = 2454 THEN
            sigmoid_f := 1573;
        ELSIF x = 2455 THEN
            sigmoid_f := 1573;
        ELSIF x = 2456 THEN
            sigmoid_f := 1573;
        ELSIF x = 2457 THEN
            sigmoid_f := 1574;
        ELSIF x = 2458 THEN
            sigmoid_f := 1574;
        ELSIF x = 2459 THEN
            sigmoid_f := 1574;
        ELSIF x = 2460 THEN
            sigmoid_f := 1574;
        ELSIF x = 2461 THEN
            sigmoid_f := 1574;
        ELSIF x = 2462 THEN
            sigmoid_f := 1575;
        ELSIF x = 2463 THEN
            sigmoid_f := 1575;
        ELSIF x = 2464 THEN
            sigmoid_f := 1575;
        ELSIF x = 2465 THEN
            sigmoid_f := 1575;
        ELSIF x = 2466 THEN
            sigmoid_f := 1575;
        ELSIF x = 2467 THEN
            sigmoid_f := 1575;
        ELSIF x = 2468 THEN
            sigmoid_f := 1576;
        ELSIF x = 2469 THEN
            sigmoid_f := 1576;
        ELSIF x = 2470 THEN
            sigmoid_f := 1576;
        ELSIF x = 2471 THEN
            sigmoid_f := 1576;
        ELSIF x = 2472 THEN
            sigmoid_f := 1576;
        ELSIF x = 2473 THEN
            sigmoid_f := 1577;
        ELSIF x = 2474 THEN
            sigmoid_f := 1577;
        ELSIF x = 2475 THEN
            sigmoid_f := 1577;
        ELSIF x = 2476 THEN
            sigmoid_f := 1577;
        ELSIF x = 2477 THEN
            sigmoid_f := 1577;
        ELSIF x = 2478 THEN
            sigmoid_f := 1577;
        ELSIF x = 2479 THEN
            sigmoid_f := 1578;
        ELSIF x = 2480 THEN
            sigmoid_f := 1578;
        ELSIF x = 2481 THEN
            sigmoid_f := 1578;
        ELSIF x = 2482 THEN
            sigmoid_f := 1578;
        ELSIF x = 2483 THEN
            sigmoid_f := 1578;
        ELSIF x = 2484 THEN
            sigmoid_f := 1579;
        ELSIF x = 2485 THEN
            sigmoid_f := 1579;
        ELSIF x = 2486 THEN
            sigmoid_f := 1579;
        ELSIF x = 2487 THEN
            sigmoid_f := 1579;
        ELSIF x = 2488 THEN
            sigmoid_f := 1579;
        ELSIF x = 2489 THEN
            sigmoid_f := 1580;
        ELSIF x = 2490 THEN
            sigmoid_f := 1580;
        ELSIF x = 2491 THEN
            sigmoid_f := 1580;
        ELSIF x = 2492 THEN
            sigmoid_f := 1580;
        ELSIF x = 2493 THEN
            sigmoid_f := 1580;
        ELSIF x = 2494 THEN
            sigmoid_f := 1580;
        ELSIF x = 2495 THEN
            sigmoid_f := 1581;
        ELSIF x = 2496 THEN
            sigmoid_f := 1581;
        ELSIF x = 2497 THEN
            sigmoid_f := 1581;
        ELSIF x = 2498 THEN
            sigmoid_f := 1581;
        ELSIF x = 2499 THEN
            sigmoid_f := 1581;
        ELSIF x = 2500 THEN
            sigmoid_f := 1582;
        ELSIF x = 2501 THEN
            sigmoid_f := 1582;
        ELSIF x = 2502 THEN
            sigmoid_f := 1582;
        ELSIF x = 2503 THEN
            sigmoid_f := 1582;
        ELSIF x = 2504 THEN
            sigmoid_f := 1582;
        ELSIF x = 2505 THEN
            sigmoid_f := 1583;
        ELSIF x = 2506 THEN
            sigmoid_f := 1583;
        ELSIF x = 2507 THEN
            sigmoid_f := 1583;
        ELSIF x = 2508 THEN
            sigmoid_f := 1583;
        ELSIF x = 2509 THEN
            sigmoid_f := 1583;
        ELSIF x = 2510 THEN
            sigmoid_f := 1583;
        ELSIF x = 2511 THEN
            sigmoid_f := 1584;
        ELSIF x = 2512 THEN
            sigmoid_f := 1584;
        ELSIF x = 2513 THEN
            sigmoid_f := 1584;
        ELSIF x = 2514 THEN
            sigmoid_f := 1584;
        ELSIF x = 2515 THEN
            sigmoid_f := 1584;
        ELSIF x = 2516 THEN
            sigmoid_f := 1585;
        ELSIF x = 2517 THEN
            sigmoid_f := 1585;
        ELSIF x = 2518 THEN
            sigmoid_f := 1585;
        ELSIF x = 2519 THEN
            sigmoid_f := 1585;
        ELSIF x = 2520 THEN
            sigmoid_f := 1585;
        ELSIF x = 2521 THEN
            sigmoid_f := 1585;
        ELSIF x = 2522 THEN
            sigmoid_f := 1586;
        ELSIF x = 2523 THEN
            sigmoid_f := 1586;
        ELSIF x = 2524 THEN
            sigmoid_f := 1586;
        ELSIF x = 2525 THEN
            sigmoid_f := 1586;
        ELSIF x = 2526 THEN
            sigmoid_f := 1586;
        ELSIF x = 2527 THEN
            sigmoid_f := 1587;
        ELSIF x = 2528 THEN
            sigmoid_f := 1587;
        ELSIF x = 2529 THEN
            sigmoid_f := 1587;
        ELSIF x = 2530 THEN
            sigmoid_f := 1587;
        ELSIF x = 2531 THEN
            sigmoid_f := 1587;
        ELSIF x = 2532 THEN
            sigmoid_f := 1588;
        ELSIF x = 2533 THEN
            sigmoid_f := 1588;
        ELSIF x = 2534 THEN
            sigmoid_f := 1588;
        ELSIF x = 2535 THEN
            sigmoid_f := 1588;
        ELSIF x = 2536 THEN
            sigmoid_f := 1588;
        ELSIF x = 2537 THEN
            sigmoid_f := 1588;
        ELSIF x = 2538 THEN
            sigmoid_f := 1589;
        ELSIF x = 2539 THEN
            sigmoid_f := 1589;
        ELSIF x = 2540 THEN
            sigmoid_f := 1589;
        ELSIF x = 2541 THEN
            sigmoid_f := 1589;
        ELSIF x = 2542 THEN
            sigmoid_f := 1589;
        ELSIF x = 2543 THEN
            sigmoid_f := 1590;
        ELSIF x = 2544 THEN
            sigmoid_f := 1590;
        ELSIF x = 2545 THEN
            sigmoid_f := 1590;
        ELSIF x = 2546 THEN
            sigmoid_f := 1590;
        ELSIF x = 2547 THEN
            sigmoid_f := 1590;
        ELSIF x = 2548 THEN
            sigmoid_f := 1591;
        ELSIF x = 2549 THEN
            sigmoid_f := 1591;
        ELSIF x = 2550 THEN
            sigmoid_f := 1591;
        ELSIF x = 2551 THEN
            sigmoid_f := 1591;
        ELSIF x = 2552 THEN
            sigmoid_f := 1591;
        ELSIF x = 2553 THEN
            sigmoid_f := 1591;
        ELSIF x = 2554 THEN
            sigmoid_f := 1592;
        ELSIF x = 2555 THEN
            sigmoid_f := 1592;
        ELSIF x = 2556 THEN
            sigmoid_f := 1592;
        ELSIF x = 2557 THEN
            sigmoid_f := 1592;
        ELSIF x = 2558 THEN
            sigmoid_f := 1592;
        ELSIF x = 2559 THEN
            sigmoid_f := 1593;
        ELSIF x = 2560 THEN
            sigmoid_f := 1593;
        ELSIF x = 2561 THEN
            sigmoid_f := 1593;
        ELSIF x = 2562 THEN
            sigmoid_f := 1593;
        ELSIF x = 2563 THEN
            sigmoid_f := 1593;
        ELSIF x = 2564 THEN
            sigmoid_f := 1593;
        ELSIF x = 2565 THEN
            sigmoid_f := 1594;
        ELSIF x = 2566 THEN
            sigmoid_f := 1594;
        ELSIF x = 2567 THEN
            sigmoid_f := 1594;
        ELSIF x = 2568 THEN
            sigmoid_f := 1594;
        ELSIF x = 2569 THEN
            sigmoid_f := 1594;
        ELSIF x = 2570 THEN
            sigmoid_f := 1594;
        ELSIF x = 2571 THEN
            sigmoid_f := 1595;
        ELSIF x = 2572 THEN
            sigmoid_f := 1595;
        ELSIF x = 2573 THEN
            sigmoid_f := 1595;
        ELSIF x = 2574 THEN
            sigmoid_f := 1595;
        ELSIF x = 2575 THEN
            sigmoid_f := 1595;
        ELSIF x = 2576 THEN
            sigmoid_f := 1595;
        ELSIF x = 2577 THEN
            sigmoid_f := 1595;
        ELSIF x = 2578 THEN
            sigmoid_f := 1596;
        ELSIF x = 2579 THEN
            sigmoid_f := 1596;
        ELSIF x = 2580 THEN
            sigmoid_f := 1596;
        ELSIF x = 2581 THEN
            sigmoid_f := 1596;
        ELSIF x = 2582 THEN
            sigmoid_f := 1596;
        ELSIF x = 2583 THEN
            sigmoid_f := 1596;
        ELSIF x = 2584 THEN
            sigmoid_f := 1597;
        ELSIF x = 2585 THEN
            sigmoid_f := 1597;
        ELSIF x = 2586 THEN
            sigmoid_f := 1597;
        ELSIF x = 2587 THEN
            sigmoid_f := 1597;
        ELSIF x = 2588 THEN
            sigmoid_f := 1597;
        ELSIF x = 2589 THEN
            sigmoid_f := 1597;
        ELSIF x = 2590 THEN
            sigmoid_f := 1598;
        ELSIF x = 2591 THEN
            sigmoid_f := 1598;
        ELSIF x = 2592 THEN
            sigmoid_f := 1598;
        ELSIF x = 2593 THEN
            sigmoid_f := 1598;
        ELSIF x = 2594 THEN
            sigmoid_f := 1598;
        ELSIF x = 2595 THEN
            sigmoid_f := 1598;
        ELSIF x = 2596 THEN
            sigmoid_f := 1599;
        ELSIF x = 2597 THEN
            sigmoid_f := 1599;
        ELSIF x = 2598 THEN
            sigmoid_f := 1599;
        ELSIF x = 2599 THEN
            sigmoid_f := 1599;
        ELSIF x = 2600 THEN
            sigmoid_f := 1599;
        ELSIF x = 2601 THEN
            sigmoid_f := 1599;
        ELSIF x = 2602 THEN
            sigmoid_f := 1599;
        ELSIF x = 2603 THEN
            sigmoid_f := 1600;
        ELSIF x = 2604 THEN
            sigmoid_f := 1600;
        ELSIF x = 2605 THEN
            sigmoid_f := 1600;
        ELSIF x = 2606 THEN
            sigmoid_f := 1600;
        ELSIF x = 2607 THEN
            sigmoid_f := 1600;
        ELSIF x = 2608 THEN
            sigmoid_f := 1600;
        ELSIF x = 2609 THEN
            sigmoid_f := 1601;
        ELSIF x = 2610 THEN
            sigmoid_f := 1601;
        ELSIF x = 2611 THEN
            sigmoid_f := 1601;
        ELSIF x = 2612 THEN
            sigmoid_f := 1601;
        ELSIF x = 2613 THEN
            sigmoid_f := 1601;
        ELSIF x = 2614 THEN
            sigmoid_f := 1601;
        ELSIF x = 2615 THEN
            sigmoid_f := 1602;
        ELSIF x = 2616 THEN
            sigmoid_f := 1602;
        ELSIF x = 2617 THEN
            sigmoid_f := 1602;
        ELSIF x = 2618 THEN
            sigmoid_f := 1602;
        ELSIF x = 2619 THEN
            sigmoid_f := 1602;
        ELSIF x = 2620 THEN
            sigmoid_f := 1602;
        ELSIF x = 2621 THEN
            sigmoid_f := 1603;
        ELSIF x = 2622 THEN
            sigmoid_f := 1603;
        ELSIF x = 2623 THEN
            sigmoid_f := 1603;
        ELSIF x = 2624 THEN
            sigmoid_f := 1603;
        ELSIF x = 2625 THEN
            sigmoid_f := 1603;
        ELSIF x = 2626 THEN
            sigmoid_f := 1603;
        ELSIF x = 2627 THEN
            sigmoid_f := 1604;
        ELSIF x = 2628 THEN
            sigmoid_f := 1604;
        ELSIF x = 2629 THEN
            sigmoid_f := 1604;
        ELSIF x = 2630 THEN
            sigmoid_f := 1604;
        ELSIF x = 2631 THEN
            sigmoid_f := 1604;
        ELSIF x = 2632 THEN
            sigmoid_f := 1604;
        ELSIF x = 2633 THEN
            sigmoid_f := 1604;
        ELSIF x = 2634 THEN
            sigmoid_f := 1605;
        ELSIF x = 2635 THEN
            sigmoid_f := 1605;
        ELSIF x = 2636 THEN
            sigmoid_f := 1605;
        ELSIF x = 2637 THEN
            sigmoid_f := 1605;
        ELSIF x = 2638 THEN
            sigmoid_f := 1605;
        ELSIF x = 2639 THEN
            sigmoid_f := 1605;
        ELSIF x = 2640 THEN
            sigmoid_f := 1606;
        ELSIF x = 2641 THEN
            sigmoid_f := 1606;
        ELSIF x = 2642 THEN
            sigmoid_f := 1606;
        ELSIF x = 2643 THEN
            sigmoid_f := 1606;
        ELSIF x = 2644 THEN
            sigmoid_f := 1606;
        ELSIF x = 2645 THEN
            sigmoid_f := 1606;
        ELSIF x = 2646 THEN
            sigmoid_f := 1607;
        ELSIF x = 2647 THEN
            sigmoid_f := 1607;
        ELSIF x = 2648 THEN
            sigmoid_f := 1607;
        ELSIF x = 2649 THEN
            sigmoid_f := 1607;
        ELSIF x = 2650 THEN
            sigmoid_f := 1607;
        ELSIF x = 2651 THEN
            sigmoid_f := 1607;
        ELSIF x = 2652 THEN
            sigmoid_f := 1608;
        ELSIF x = 2653 THEN
            sigmoid_f := 1608;
        ELSIF x = 2654 THEN
            sigmoid_f := 1608;
        ELSIF x = 2655 THEN
            sigmoid_f := 1608;
        ELSIF x = 2656 THEN
            sigmoid_f := 1608;
        ELSIF x = 2657 THEN
            sigmoid_f := 1608;
        ELSIF x = 2658 THEN
            sigmoid_f := 1608;
        ELSIF x = 2659 THEN
            sigmoid_f := 1609;
        ELSIF x = 2660 THEN
            sigmoid_f := 1609;
        ELSIF x = 2661 THEN
            sigmoid_f := 1609;
        ELSIF x = 2662 THEN
            sigmoid_f := 1609;
        ELSIF x = 2663 THEN
            sigmoid_f := 1609;
        ELSIF x = 2664 THEN
            sigmoid_f := 1609;
        ELSIF x = 2665 THEN
            sigmoid_f := 1610;
        ELSIF x = 2666 THEN
            sigmoid_f := 1610;
        ELSIF x = 2667 THEN
            sigmoid_f := 1610;
        ELSIF x = 2668 THEN
            sigmoid_f := 1610;
        ELSIF x = 2669 THEN
            sigmoid_f := 1610;
        ELSIF x = 2670 THEN
            sigmoid_f := 1610;
        ELSIF x = 2671 THEN
            sigmoid_f := 1611;
        ELSIF x = 2672 THEN
            sigmoid_f := 1611;
        ELSIF x = 2673 THEN
            sigmoid_f := 1611;
        ELSIF x = 2674 THEN
            sigmoid_f := 1611;
        ELSIF x = 2675 THEN
            sigmoid_f := 1611;
        ELSIF x = 2676 THEN
            sigmoid_f := 1611;
        ELSIF x = 2677 THEN
            sigmoid_f := 1612;
        ELSIF x = 2678 THEN
            sigmoid_f := 1612;
        ELSIF x = 2679 THEN
            sigmoid_f := 1612;
        ELSIF x = 2680 THEN
            sigmoid_f := 1612;
        ELSIF x = 2681 THEN
            sigmoid_f := 1612;
        ELSIF x = 2682 THEN
            sigmoid_f := 1612;
        ELSIF x = 2683 THEN
            sigmoid_f := 1613;
        ELSIF x = 2684 THEN
            sigmoid_f := 1613;
        ELSIF x = 2685 THEN
            sigmoid_f := 1613;
        ELSIF x = 2686 THEN
            sigmoid_f := 1613;
        ELSIF x = 2687 THEN
            sigmoid_f := 1613;
        ELSIF x = 2688 THEN
            sigmoid_f := 1613;
        ELSIF x = 2689 THEN
            sigmoid_f := 1613;
        ELSIF x = 2690 THEN
            sigmoid_f := 1614;
        ELSIF x = 2691 THEN
            sigmoid_f := 1614;
        ELSIF x = 2692 THEN
            sigmoid_f := 1614;
        ELSIF x = 2693 THEN
            sigmoid_f := 1614;
        ELSIF x = 2694 THEN
            sigmoid_f := 1614;
        ELSIF x = 2695 THEN
            sigmoid_f := 1614;
        ELSIF x = 2696 THEN
            sigmoid_f := 1615;
        ELSIF x = 2697 THEN
            sigmoid_f := 1615;
        ELSIF x = 2698 THEN
            sigmoid_f := 1615;
        ELSIF x = 2699 THEN
            sigmoid_f := 1615;
        ELSIF x = 2700 THEN
            sigmoid_f := 1615;
        ELSIF x = 2701 THEN
            sigmoid_f := 1615;
        ELSIF x = 2702 THEN
            sigmoid_f := 1616;
        ELSIF x = 2703 THEN
            sigmoid_f := 1616;
        ELSIF x = 2704 THEN
            sigmoid_f := 1616;
        ELSIF x = 2705 THEN
            sigmoid_f := 1616;
        ELSIF x = 2706 THEN
            sigmoid_f := 1616;
        ELSIF x = 2707 THEN
            sigmoid_f := 1616;
        ELSIF x = 2708 THEN
            sigmoid_f := 1617;
        ELSIF x = 2709 THEN
            sigmoid_f := 1617;
        ELSIF x = 2710 THEN
            sigmoid_f := 1617;
        ELSIF x = 2711 THEN
            sigmoid_f := 1617;
        ELSIF x = 2712 THEN
            sigmoid_f := 1617;
        ELSIF x = 2713 THEN
            sigmoid_f := 1617;
        ELSIF x = 2714 THEN
            sigmoid_f := 1617;
        ELSIF x = 2715 THEN
            sigmoid_f := 1618;
        ELSIF x = 2716 THEN
            sigmoid_f := 1618;
        ELSIF x = 2717 THEN
            sigmoid_f := 1618;
        ELSIF x = 2718 THEN
            sigmoid_f := 1618;
        ELSIF x = 2719 THEN
            sigmoid_f := 1618;
        ELSIF x = 2720 THEN
            sigmoid_f := 1618;
        ELSIF x = 2721 THEN
            sigmoid_f := 1619;
        ELSIF x = 2722 THEN
            sigmoid_f := 1619;
        ELSIF x = 2723 THEN
            sigmoid_f := 1619;
        ELSIF x = 2724 THEN
            sigmoid_f := 1619;
        ELSIF x = 2725 THEN
            sigmoid_f := 1619;
        ELSIF x = 2726 THEN
            sigmoid_f := 1619;
        ELSIF x = 2727 THEN
            sigmoid_f := 1620;
        ELSIF x = 2728 THEN
            sigmoid_f := 1620;
        ELSIF x = 2729 THEN
            sigmoid_f := 1620;
        ELSIF x = 2730 THEN
            sigmoid_f := 1620;
        ELSIF x = 2731 THEN
            sigmoid_f := 1620;
        ELSIF x = 2732 THEN
            sigmoid_f := 1620;
        ELSIF x = 2733 THEN
            sigmoid_f := 1621;
        ELSIF x = 2734 THEN
            sigmoid_f := 1621;
        ELSIF x = 2735 THEN
            sigmoid_f := 1621;
        ELSIF x = 2736 THEN
            sigmoid_f := 1621;
        ELSIF x = 2737 THEN
            sigmoid_f := 1621;
        ELSIF x = 2738 THEN
            sigmoid_f := 1621;
        ELSIF x = 2739 THEN
            sigmoid_f := 1622;
        ELSIF x = 2740 THEN
            sigmoid_f := 1622;
        ELSIF x = 2741 THEN
            sigmoid_f := 1622;
        ELSIF x = 2742 THEN
            sigmoid_f := 1622;
        ELSIF x = 2743 THEN
            sigmoid_f := 1622;
        ELSIF x = 2744 THEN
            sigmoid_f := 1622;
        ELSIF x = 2745 THEN
            sigmoid_f := 1622;
        ELSIF x = 2746 THEN
            sigmoid_f := 1623;
        ELSIF x = 2747 THEN
            sigmoid_f := 1623;
        ELSIF x = 2748 THEN
            sigmoid_f := 1623;
        ELSIF x = 2749 THEN
            sigmoid_f := 1623;
        ELSIF x = 2750 THEN
            sigmoid_f := 1623;
        ELSIF x = 2751 THEN
            sigmoid_f := 1623;
        ELSIF x = 2752 THEN
            sigmoid_f := 1624;
        ELSIF x = 2753 THEN
            sigmoid_f := 1624;
        ELSIF x = 2754 THEN
            sigmoid_f := 1624;
        ELSIF x = 2755 THEN
            sigmoid_f := 1624;
        ELSIF x = 2756 THEN
            sigmoid_f := 1624;
        ELSIF x = 2757 THEN
            sigmoid_f := 1624;
        ELSIF x = 2758 THEN
            sigmoid_f := 1625;
        ELSIF x = 2759 THEN
            sigmoid_f := 1625;
        ELSIF x = 2760 THEN
            sigmoid_f := 1625;
        ELSIF x = 2761 THEN
            sigmoid_f := 1625;
        ELSIF x = 2762 THEN
            sigmoid_f := 1625;
        ELSIF x = 2763 THEN
            sigmoid_f := 1625;
        ELSIF x = 2764 THEN
            sigmoid_f := 1626;
        ELSIF x = 2765 THEN
            sigmoid_f := 1626;
        ELSIF x = 2766 THEN
            sigmoid_f := 1626;
        ELSIF x = 2767 THEN
            sigmoid_f := 1626;
        ELSIF x = 2768 THEN
            sigmoid_f := 1626;
        ELSIF x = 2769 THEN
            sigmoid_f := 1626;
        ELSIF x = 2770 THEN
            sigmoid_f := 1626;
        ELSIF x = 2771 THEN
            sigmoid_f := 1627;
        ELSIF x = 2772 THEN
            sigmoid_f := 1627;
        ELSIF x = 2773 THEN
            sigmoid_f := 1627;
        ELSIF x = 2774 THEN
            sigmoid_f := 1627;
        ELSIF x = 2775 THEN
            sigmoid_f := 1627;
        ELSIF x = 2776 THEN
            sigmoid_f := 1627;
        ELSIF x = 2777 THEN
            sigmoid_f := 1628;
        ELSIF x = 2778 THEN
            sigmoid_f := 1628;
        ELSIF x = 2779 THEN
            sigmoid_f := 1628;
        ELSIF x = 2780 THEN
            sigmoid_f := 1628;
        ELSIF x = 2781 THEN
            sigmoid_f := 1628;
        ELSIF x = 2782 THEN
            sigmoid_f := 1628;
        ELSIF x = 2783 THEN
            sigmoid_f := 1629;
        ELSIF x = 2784 THEN
            sigmoid_f := 1629;
        ELSIF x = 2785 THEN
            sigmoid_f := 1629;
        ELSIF x = 2786 THEN
            sigmoid_f := 1629;
        ELSIF x = 2787 THEN
            sigmoid_f := 1629;
        ELSIF x = 2788 THEN
            sigmoid_f := 1629;
        ELSIF x = 2789 THEN
            sigmoid_f := 1630;
        ELSIF x = 2790 THEN
            sigmoid_f := 1630;
        ELSIF x = 2791 THEN
            sigmoid_f := 1630;
        ELSIF x = 2792 THEN
            sigmoid_f := 1630;
        ELSIF x = 2793 THEN
            sigmoid_f := 1630;
        ELSIF x = 2794 THEN
            sigmoid_f := 1630;
        ELSIF x = 2795 THEN
            sigmoid_f := 1631;
        ELSIF x = 2796 THEN
            sigmoid_f := 1631;
        ELSIF x = 2797 THEN
            sigmoid_f := 1631;
        ELSIF x = 2798 THEN
            sigmoid_f := 1631;
        ELSIF x = 2799 THEN
            sigmoid_f := 1631;
        ELSIF x = 2800 THEN
            sigmoid_f := 1631;
        ELSIF x = 2801 THEN
            sigmoid_f := 1631;
        ELSIF x = 2802 THEN
            sigmoid_f := 1632;
        ELSIF x = 2803 THEN
            sigmoid_f := 1632;
        ELSIF x = 2804 THEN
            sigmoid_f := 1632;
        ELSIF x = 2805 THEN
            sigmoid_f := 1632;
        ELSIF x = 2806 THEN
            sigmoid_f := 1632;
        ELSIF x = 2807 THEN
            sigmoid_f := 1632;
        ELSIF x = 2808 THEN
            sigmoid_f := 1633;
        ELSIF x = 2809 THEN
            sigmoid_f := 1633;
        ELSIF x = 2810 THEN
            sigmoid_f := 1633;
        ELSIF x = 2811 THEN
            sigmoid_f := 1633;
        ELSIF x = 2812 THEN
            sigmoid_f := 1633;
        ELSIF x = 2813 THEN
            sigmoid_f := 1633;
        ELSIF x = 2814 THEN
            sigmoid_f := 1634;
        ELSIF x = 2815 THEN
            sigmoid_f := 1634;
        ELSIF x = 2816 THEN
            sigmoid_f := 1634;
        ELSIF x = 2817 THEN
            sigmoid_f := 1634;
        ELSIF x = 2818 THEN
            sigmoid_f := 1634;
        ELSIF x = 2819 THEN
            sigmoid_f := 1634;
        ELSIF x = 2820 THEN
            sigmoid_f := 1635;
        ELSIF x = 2821 THEN
            sigmoid_f := 1635;
        ELSIF x = 2822 THEN
            sigmoid_f := 1635;
        ELSIF x = 2823 THEN
            sigmoid_f := 1635;
        ELSIF x = 2824 THEN
            sigmoid_f := 1635;
        ELSIF x = 2825 THEN
            sigmoid_f := 1635;
        ELSIF x = 2826 THEN
            sigmoid_f := 1635;
        ELSIF x = 2827 THEN
            sigmoid_f := 1636;
        ELSIF x = 2828 THEN
            sigmoid_f := 1636;
        ELSIF x = 2829 THEN
            sigmoid_f := 1636;
        ELSIF x = 2830 THEN
            sigmoid_f := 1636;
        ELSIF x = 2831 THEN
            sigmoid_f := 1636;
        ELSIF x = 2832 THEN
            sigmoid_f := 1636;
        ELSIF x = 2833 THEN
            sigmoid_f := 1637;
        ELSIF x = 2834 THEN
            sigmoid_f := 1637;
        ELSIF x = 2835 THEN
            sigmoid_f := 1637;
        ELSIF x = 2836 THEN
            sigmoid_f := 1637;
        ELSIF x = 2837 THEN
            sigmoid_f := 1637;
        ELSIF x = 2838 THEN
            sigmoid_f := 1637;
        ELSIF x = 2839 THEN
            sigmoid_f := 1638;
        ELSIF x = 2840 THEN
            sigmoid_f := 1638;
        ELSIF x = 2841 THEN
            sigmoid_f := 1638;
        ELSIF x = 2842 THEN
            sigmoid_f := 1638;
        ELSIF x = 2843 THEN
            sigmoid_f := 1638;
        ELSIF x = 2844 THEN
            sigmoid_f := 1638;
        ELSIF x = 2845 THEN
            sigmoid_f := 1639;
        ELSIF x = 2846 THEN
            sigmoid_f := 1639;
        ELSIF x = 2847 THEN
            sigmoid_f := 1639;
        ELSIF x = 2848 THEN
            sigmoid_f := 1639;
        ELSIF x = 2849 THEN
            sigmoid_f := 1639;
        ELSIF x = 2850 THEN
            sigmoid_f := 1639;
        ELSIF x = 2851 THEN
            sigmoid_f := 1639;
        ELSIF x = 2852 THEN
            sigmoid_f := 1640;
        ELSIF x = 2853 THEN
            sigmoid_f := 1640;
        ELSIF x = 2854 THEN
            sigmoid_f := 1640;
        ELSIF x = 2855 THEN
            sigmoid_f := 1640;
        ELSIF x = 2856 THEN
            sigmoid_f := 1640;
        ELSIF x = 2857 THEN
            sigmoid_f := 1640;
        ELSIF x = 2858 THEN
            sigmoid_f := 1641;
        ELSIF x = 2859 THEN
            sigmoid_f := 1641;
        ELSIF x = 2860 THEN
            sigmoid_f := 1641;
        ELSIF x = 2861 THEN
            sigmoid_f := 1641;
        ELSIF x = 2862 THEN
            sigmoid_f := 1641;
        ELSIF x = 2863 THEN
            sigmoid_f := 1641;
        ELSIF x = 2864 THEN
            sigmoid_f := 1642;
        ELSIF x = 2865 THEN
            sigmoid_f := 1642;
        ELSIF x = 2866 THEN
            sigmoid_f := 1642;
        ELSIF x = 2867 THEN
            sigmoid_f := 1642;
        ELSIF x = 2868 THEN
            sigmoid_f := 1642;
        ELSIF x = 2869 THEN
            sigmoid_f := 1642;
        ELSIF x = 2870 THEN
            sigmoid_f := 1643;
        ELSIF x = 2871 THEN
            sigmoid_f := 1643;
        ELSIF x = 2872 THEN
            sigmoid_f := 1643;
        ELSIF x = 2873 THEN
            sigmoid_f := 1643;
        ELSIF x = 2874 THEN
            sigmoid_f := 1643;
        ELSIF x = 2875 THEN
            sigmoid_f := 1643;
        ELSIF x = 2876 THEN
            sigmoid_f := 1644;
        ELSIF x = 2877 THEN
            sigmoid_f := 1644;
        ELSIF x = 2878 THEN
            sigmoid_f := 1644;
        ELSIF x = 2879 THEN
            sigmoid_f := 1644;
        ELSIF x = 2880 THEN
            sigmoid_f := 1644;
        ELSIF x = 2881 THEN
            sigmoid_f := 1644;
        ELSIF x = 2882 THEN
            sigmoid_f := 1644;
        ELSIF x = 2883 THEN
            sigmoid_f := 1645;
        ELSIF x = 2884 THEN
            sigmoid_f := 1645;
        ELSIF x = 2885 THEN
            sigmoid_f := 1645;
        ELSIF x = 2886 THEN
            sigmoid_f := 1645;
        ELSIF x = 2887 THEN
            sigmoid_f := 1645;
        ELSIF x = 2888 THEN
            sigmoid_f := 1645;
        ELSIF x = 2889 THEN
            sigmoid_f := 1646;
        ELSIF x = 2890 THEN
            sigmoid_f := 1646;
        ELSIF x = 2891 THEN
            sigmoid_f := 1646;
        ELSIF x = 2892 THEN
            sigmoid_f := 1646;
        ELSIF x = 2893 THEN
            sigmoid_f := 1646;
        ELSIF x = 2894 THEN
            sigmoid_f := 1646;
        ELSIF x = 2895 THEN
            sigmoid_f := 1647;
        ELSIF x = 2896 THEN
            sigmoid_f := 1647;
        ELSIF x = 2897 THEN
            sigmoid_f := 1647;
        ELSIF x = 2898 THEN
            sigmoid_f := 1647;
        ELSIF x = 2899 THEN
            sigmoid_f := 1647;
        ELSIF x = 2900 THEN
            sigmoid_f := 1647;
        ELSIF x = 2901 THEN
            sigmoid_f := 1648;
        ELSIF x = 2902 THEN
            sigmoid_f := 1648;
        ELSIF x = 2903 THEN
            sigmoid_f := 1648;
        ELSIF x = 2904 THEN
            sigmoid_f := 1648;
        ELSIF x = 2905 THEN
            sigmoid_f := 1648;
        ELSIF x = 2906 THEN
            sigmoid_f := 1648;
        ELSIF x = 2907 THEN
            sigmoid_f := 1648;
        ELSIF x = 2908 THEN
            sigmoid_f := 1649;
        ELSIF x = 2909 THEN
            sigmoid_f := 1649;
        ELSIF x = 2910 THEN
            sigmoid_f := 1649;
        ELSIF x = 2911 THEN
            sigmoid_f := 1649;
        ELSIF x = 2912 THEN
            sigmoid_f := 1649;
        ELSIF x = 2913 THEN
            sigmoid_f := 1649;
        ELSIF x = 2914 THEN
            sigmoid_f := 1650;
        ELSIF x = 2915 THEN
            sigmoid_f := 1650;
        ELSIF x = 2916 THEN
            sigmoid_f := 1650;
        ELSIF x = 2917 THEN
            sigmoid_f := 1650;
        ELSIF x = 2918 THEN
            sigmoid_f := 1650;
        ELSIF x = 2919 THEN
            sigmoid_f := 1650;
        ELSIF x = 2920 THEN
            sigmoid_f := 1651;
        ELSIF x = 2921 THEN
            sigmoid_f := 1651;
        ELSIF x = 2922 THEN
            sigmoid_f := 1651;
        ELSIF x = 2923 THEN
            sigmoid_f := 1651;
        ELSIF x = 2924 THEN
            sigmoid_f := 1651;
        ELSIF x = 2925 THEN
            sigmoid_f := 1651;
        ELSIF x = 2926 THEN
            sigmoid_f := 1652;
        ELSIF x = 2927 THEN
            sigmoid_f := 1652;
        ELSIF x = 2928 THEN
            sigmoid_f := 1652;
        ELSIF x = 2929 THEN
            sigmoid_f := 1652;
        ELSIF x = 2930 THEN
            sigmoid_f := 1652;
        ELSIF x = 2931 THEN
            sigmoid_f := 1652;
        ELSIF x = 2932 THEN
            sigmoid_f := 1653;
        ELSIF x = 2933 THEN
            sigmoid_f := 1653;
        ELSIF x = 2934 THEN
            sigmoid_f := 1653;
        ELSIF x = 2935 THEN
            sigmoid_f := 1653;
        ELSIF x = 2936 THEN
            sigmoid_f := 1653;
        ELSIF x = 2937 THEN
            sigmoid_f := 1653;
        ELSIF x = 2938 THEN
            sigmoid_f := 1653;
        ELSIF x = 2939 THEN
            sigmoid_f := 1654;
        ELSIF x = 2940 THEN
            sigmoid_f := 1654;
        ELSIF x = 2941 THEN
            sigmoid_f := 1654;
        ELSIF x = 2942 THEN
            sigmoid_f := 1654;
        ELSIF x = 2943 THEN
            sigmoid_f := 1654;
        ELSIF x = 2944 THEN
            sigmoid_f := 1654;
        ELSIF x = 2945 THEN
            sigmoid_f := 1655;
        ELSIF x = 2946 THEN
            sigmoid_f := 1655;
        ELSIF x = 2947 THEN
            sigmoid_f := 1655;
        ELSIF x = 2948 THEN
            sigmoid_f := 1655;
        ELSIF x = 2949 THEN
            sigmoid_f := 1655;
        ELSIF x = 2950 THEN
            sigmoid_f := 1655;
        ELSIF x = 2951 THEN
            sigmoid_f := 1656;
        ELSIF x = 2952 THEN
            sigmoid_f := 1656;
        ELSIF x = 2953 THEN
            sigmoid_f := 1656;
        ELSIF x = 2954 THEN
            sigmoid_f := 1656;
        ELSIF x = 2955 THEN
            sigmoid_f := 1656;
        ELSIF x = 2956 THEN
            sigmoid_f := 1656;
        ELSIF x = 2957 THEN
            sigmoid_f := 1657;
        ELSIF x = 2958 THEN
            sigmoid_f := 1657;
        ELSIF x = 2959 THEN
            sigmoid_f := 1657;
        ELSIF x = 2960 THEN
            sigmoid_f := 1657;
        ELSIF x = 2961 THEN
            sigmoid_f := 1657;
        ELSIF x = 2962 THEN
            sigmoid_f := 1657;
        ELSIF x = 2963 THEN
            sigmoid_f := 1657;
        ELSIF x = 2964 THEN
            sigmoid_f := 1658;
        ELSIF x = 2965 THEN
            sigmoid_f := 1658;
        ELSIF x = 2966 THEN
            sigmoid_f := 1658;
        ELSIF x = 2967 THEN
            sigmoid_f := 1658;
        ELSIF x = 2968 THEN
            sigmoid_f := 1658;
        ELSIF x = 2969 THEN
            sigmoid_f := 1658;
        ELSIF x = 2970 THEN
            sigmoid_f := 1659;
        ELSIF x = 2971 THEN
            sigmoid_f := 1659;
        ELSIF x = 2972 THEN
            sigmoid_f := 1659;
        ELSIF x = 2973 THEN
            sigmoid_f := 1659;
        ELSIF x = 2974 THEN
            sigmoid_f := 1659;
        ELSIF x = 2975 THEN
            sigmoid_f := 1659;
        ELSIF x = 2976 THEN
            sigmoid_f := 1660;
        ELSIF x = 2977 THEN
            sigmoid_f := 1660;
        ELSIF x = 2978 THEN
            sigmoid_f := 1660;
        ELSIF x = 2979 THEN
            sigmoid_f := 1660;
        ELSIF x = 2980 THEN
            sigmoid_f := 1660;
        ELSIF x = 2981 THEN
            sigmoid_f := 1660;
        ELSIF x = 2982 THEN
            sigmoid_f := 1661;
        ELSIF x = 2983 THEN
            sigmoid_f := 1661;
        ELSIF x = 2984 THEN
            sigmoid_f := 1661;
        ELSIF x = 2985 THEN
            sigmoid_f := 1661;
        ELSIF x = 2986 THEN
            sigmoid_f := 1661;
        ELSIF x = 2987 THEN
            sigmoid_f := 1661;
        ELSIF x = 2988 THEN
            sigmoid_f := 1662;
        ELSIF x = 2989 THEN
            sigmoid_f := 1662;
        ELSIF x = 2990 THEN
            sigmoid_f := 1662;
        ELSIF x = 2991 THEN
            sigmoid_f := 1662;
        ELSIF x = 2992 THEN
            sigmoid_f := 1662;
        ELSIF x = 2993 THEN
            sigmoid_f := 1662;
        ELSIF x = 2994 THEN
            sigmoid_f := 1662;
        ELSIF x = 2995 THEN
            sigmoid_f := 1663;
        ELSIF x = 2996 THEN
            sigmoid_f := 1663;
        ELSIF x = 2997 THEN
            sigmoid_f := 1663;
        ELSIF x = 2998 THEN
            sigmoid_f := 1663;
        ELSIF x = 2999 THEN
            sigmoid_f := 1663;
        ELSIF x = 3000 THEN
            sigmoid_f := 1663;
        ELSIF x = 3001 THEN
            sigmoid_f := 1664;
        ELSIF x = 3002 THEN
            sigmoid_f := 1664;
        ELSIF x = 3003 THEN
            sigmoid_f := 1664;
        ELSIF x = 3004 THEN
            sigmoid_f := 1664;
        ELSIF x = 3005 THEN
            sigmoid_f := 1664;
        ELSIF x = 3006 THEN
            sigmoid_f := 1664;
        ELSIF x = 3007 THEN
            sigmoid_f := 1665;
        ELSIF x = 3008 THEN
            sigmoid_f := 1665;
        ELSIF x = 3009 THEN
            sigmoid_f := 1665;
        ELSIF x = 3010 THEN
            sigmoid_f := 1665;
        ELSIF x = 3011 THEN
            sigmoid_f := 1665;
        ELSIF x = 3012 THEN
            sigmoid_f := 1665;
        ELSIF x = 3013 THEN
            sigmoid_f := 1666;
        ELSIF x = 3014 THEN
            sigmoid_f := 1666;
        ELSIF x = 3015 THEN
            sigmoid_f := 1666;
        ELSIF x = 3016 THEN
            sigmoid_f := 1666;
        ELSIF x = 3017 THEN
            sigmoid_f := 1666;
        ELSIF x = 3018 THEN
            sigmoid_f := 1666;
        ELSIF x = 3019 THEN
            sigmoid_f := 1666;
        ELSIF x = 3020 THEN
            sigmoid_f := 1667;
        ELSIF x = 3021 THEN
            sigmoid_f := 1667;
        ELSIF x = 3022 THEN
            sigmoid_f := 1667;
        ELSIF x = 3023 THEN
            sigmoid_f := 1667;
        ELSIF x = 3024 THEN
            sigmoid_f := 1667;
        ELSIF x = 3025 THEN
            sigmoid_f := 1667;
        ELSIF x = 3026 THEN
            sigmoid_f := 1668;
        ELSIF x = 3027 THEN
            sigmoid_f := 1668;
        ELSIF x = 3028 THEN
            sigmoid_f := 1668;
        ELSIF x = 3029 THEN
            sigmoid_f := 1668;
        ELSIF x = 3030 THEN
            sigmoid_f := 1668;
        ELSIF x = 3031 THEN
            sigmoid_f := 1668;
        ELSIF x = 3032 THEN
            sigmoid_f := 1669;
        ELSIF x = 3033 THEN
            sigmoid_f := 1669;
        ELSIF x = 3034 THEN
            sigmoid_f := 1669;
        ELSIF x = 3035 THEN
            sigmoid_f := 1669;
        ELSIF x = 3036 THEN
            sigmoid_f := 1669;
        ELSIF x = 3037 THEN
            sigmoid_f := 1669;
        ELSIF x = 3038 THEN
            sigmoid_f := 1670;
        ELSIF x = 3039 THEN
            sigmoid_f := 1670;
        ELSIF x = 3040 THEN
            sigmoid_f := 1670;
        ELSIF x = 3041 THEN
            sigmoid_f := 1670;
        ELSIF x = 3042 THEN
            sigmoid_f := 1670;
        ELSIF x = 3043 THEN
            sigmoid_f := 1670;
        ELSIF x = 3044 THEN
            sigmoid_f := 1671;
        ELSIF x = 3045 THEN
            sigmoid_f := 1671;
        ELSIF x = 3046 THEN
            sigmoid_f := 1671;
        ELSIF x = 3047 THEN
            sigmoid_f := 1671;
        ELSIF x = 3048 THEN
            sigmoid_f := 1671;
        ELSIF x = 3049 THEN
            sigmoid_f := 1671;
        ELSIF x = 3050 THEN
            sigmoid_f := 1671;
        ELSIF x = 3051 THEN
            sigmoid_f := 1672;
        ELSIF x = 3052 THEN
            sigmoid_f := 1672;
        ELSIF x = 3053 THEN
            sigmoid_f := 1672;
        ELSIF x = 3054 THEN
            sigmoid_f := 1672;
        ELSIF x = 3055 THEN
            sigmoid_f := 1672;
        ELSIF x = 3056 THEN
            sigmoid_f := 1672;
        ELSIF x = 3057 THEN
            sigmoid_f := 1673;
        ELSIF x = 3058 THEN
            sigmoid_f := 1673;
        ELSIF x = 3059 THEN
            sigmoid_f := 1673;
        ELSIF x = 3060 THEN
            sigmoid_f := 1673;
        ELSIF x = 3061 THEN
            sigmoid_f := 1673;
        ELSIF x = 3062 THEN
            sigmoid_f := 1673;
        ELSIF x = 3063 THEN
            sigmoid_f := 1674;
        ELSIF x = 3064 THEN
            sigmoid_f := 1674;
        ELSIF x = 3065 THEN
            sigmoid_f := 1674;
        ELSIF x = 3066 THEN
            sigmoid_f := 1674;
        ELSIF x = 3067 THEN
            sigmoid_f := 1674;
        ELSIF x = 3068 THEN
            sigmoid_f := 1674;
        ELSIF x = 3069 THEN
            sigmoid_f := 1675;
        ELSIF x = 3070 THEN
            sigmoid_f := 1675;
        ELSIF x = 3071 THEN
            sigmoid_f := 1675;
        ELSIF x = 3072 THEN
            sigmoid_f := 1675;
        ELSIF x = 3073 THEN
            sigmoid_f := 1675;
        ELSIF x = 3074 THEN
            sigmoid_f := 1675;
        ELSIF x = 3075 THEN
            sigmoid_f := 1675;
        ELSIF x = 3076 THEN
            sigmoid_f := 1676;
        ELSIF x = 3077 THEN
            sigmoid_f := 1676;
        ELSIF x = 3078 THEN
            sigmoid_f := 1676;
        ELSIF x = 3079 THEN
            sigmoid_f := 1676;
        ELSIF x = 3080 THEN
            sigmoid_f := 1676;
        ELSIF x = 3081 THEN
            sigmoid_f := 1676;
        ELSIF x = 3082 THEN
            sigmoid_f := 1676;
        ELSIF x = 3083 THEN
            sigmoid_f := 1677;
        ELSIF x = 3084 THEN
            sigmoid_f := 1677;
        ELSIF x = 3085 THEN
            sigmoid_f := 1677;
        ELSIF x = 3086 THEN
            sigmoid_f := 1677;
        ELSIF x = 3087 THEN
            sigmoid_f := 1677;
        ELSIF x = 3088 THEN
            sigmoid_f := 1677;
        ELSIF x = 3089 THEN
            sigmoid_f := 1677;
        ELSIF x = 3090 THEN
            sigmoid_f := 1677;
        ELSIF x = 3091 THEN
            sigmoid_f := 1678;
        ELSIF x = 3092 THEN
            sigmoid_f := 1678;
        ELSIF x = 3093 THEN
            sigmoid_f := 1678;
        ELSIF x = 3094 THEN
            sigmoid_f := 1678;
        ELSIF x = 3095 THEN
            sigmoid_f := 1678;
        ELSIF x = 3096 THEN
            sigmoid_f := 1678;
        ELSIF x = 3097 THEN
            sigmoid_f := 1678;
        ELSIF x = 3098 THEN
            sigmoid_f := 1679;
        ELSIF x = 3099 THEN
            sigmoid_f := 1679;
        ELSIF x = 3100 THEN
            sigmoid_f := 1679;
        ELSIF x = 3101 THEN
            sigmoid_f := 1679;
        ELSIF x = 3102 THEN
            sigmoid_f := 1679;
        ELSIF x = 3103 THEN
            sigmoid_f := 1679;
        ELSIF x = 3104 THEN
            sigmoid_f := 1679;
        ELSIF x = 3105 THEN
            sigmoid_f := 1680;
        ELSIF x = 3106 THEN
            sigmoid_f := 1680;
        ELSIF x = 3107 THEN
            sigmoid_f := 1680;
        ELSIF x = 3108 THEN
            sigmoid_f := 1680;
        ELSIF x = 3109 THEN
            sigmoid_f := 1680;
        ELSIF x = 3110 THEN
            sigmoid_f := 1680;
        ELSIF x = 3111 THEN
            sigmoid_f := 1680;
        ELSIF x = 3112 THEN
            sigmoid_f := 1680;
        ELSIF x = 3113 THEN
            sigmoid_f := 1681;
        ELSIF x = 3114 THEN
            sigmoid_f := 1681;
        ELSIF x = 3115 THEN
            sigmoid_f := 1681;
        ELSIF x = 3116 THEN
            sigmoid_f := 1681;
        ELSIF x = 3117 THEN
            sigmoid_f := 1681;
        ELSIF x = 3118 THEN
            sigmoid_f := 1681;
        ELSIF x = 3119 THEN
            sigmoid_f := 1681;
        ELSIF x = 3120 THEN
            sigmoid_f := 1682;
        ELSIF x = 3121 THEN
            sigmoid_f := 1682;
        ELSIF x = 3122 THEN
            sigmoid_f := 1682;
        ELSIF x = 3123 THEN
            sigmoid_f := 1682;
        ELSIF x = 3124 THEN
            sigmoid_f := 1682;
        ELSIF x = 3125 THEN
            sigmoid_f := 1682;
        ELSIF x = 3126 THEN
            sigmoid_f := 1682;
        ELSIF x = 3127 THEN
            sigmoid_f := 1683;
        ELSIF x = 3128 THEN
            sigmoid_f := 1683;
        ELSIF x = 3129 THEN
            sigmoid_f := 1683;
        ELSIF x = 3130 THEN
            sigmoid_f := 1683;
        ELSIF x = 3131 THEN
            sigmoid_f := 1683;
        ELSIF x = 3132 THEN
            sigmoid_f := 1683;
        ELSIF x = 3133 THEN
            sigmoid_f := 1683;
        ELSIF x = 3134 THEN
            sigmoid_f := 1684;
        ELSIF x = 3135 THEN
            sigmoid_f := 1684;
        ELSIF x = 3136 THEN
            sigmoid_f := 1684;
        ELSIF x = 3137 THEN
            sigmoid_f := 1684;
        ELSIF x = 3138 THEN
            sigmoid_f := 1684;
        ELSIF x = 3139 THEN
            sigmoid_f := 1684;
        ELSIF x = 3140 THEN
            sigmoid_f := 1684;
        ELSIF x = 3141 THEN
            sigmoid_f := 1684;
        ELSIF x = 3142 THEN
            sigmoid_f := 1685;
        ELSIF x = 3143 THEN
            sigmoid_f := 1685;
        ELSIF x = 3144 THEN
            sigmoid_f := 1685;
        ELSIF x = 3145 THEN
            sigmoid_f := 1685;
        ELSIF x = 3146 THEN
            sigmoid_f := 1685;
        ELSIF x = 3147 THEN
            sigmoid_f := 1685;
        ELSIF x = 3148 THEN
            sigmoid_f := 1685;
        ELSIF x = 3149 THEN
            sigmoid_f := 1686;
        ELSIF x = 3150 THEN
            sigmoid_f := 1686;
        ELSIF x = 3151 THEN
            sigmoid_f := 1686;
        ELSIF x = 3152 THEN
            sigmoid_f := 1686;
        ELSIF x = 3153 THEN
            sigmoid_f := 1686;
        ELSIF x = 3154 THEN
            sigmoid_f := 1686;
        ELSIF x = 3155 THEN
            sigmoid_f := 1686;
        ELSIF x = 3156 THEN
            sigmoid_f := 1687;
        ELSIF x = 3157 THEN
            sigmoid_f := 1687;
        ELSIF x = 3158 THEN
            sigmoid_f := 1687;
        ELSIF x = 3159 THEN
            sigmoid_f := 1687;
        ELSIF x = 3160 THEN
            sigmoid_f := 1687;
        ELSIF x = 3161 THEN
            sigmoid_f := 1687;
        ELSIF x = 3162 THEN
            sigmoid_f := 1687;
        ELSIF x = 3163 THEN
            sigmoid_f := 1687;
        ELSIF x = 3164 THEN
            sigmoid_f := 1688;
        ELSIF x = 3165 THEN
            sigmoid_f := 1688;
        ELSIF x = 3166 THEN
            sigmoid_f := 1688;
        ELSIF x = 3167 THEN
            sigmoid_f := 1688;
        ELSIF x = 3168 THEN
            sigmoid_f := 1688;
        ELSIF x = 3169 THEN
            sigmoid_f := 1688;
        ELSIF x = 3170 THEN
            sigmoid_f := 1688;
        ELSIF x = 3171 THEN
            sigmoid_f := 1689;
        ELSIF x = 3172 THEN
            sigmoid_f := 1689;
        ELSIF x = 3173 THEN
            sigmoid_f := 1689;
        ELSIF x = 3174 THEN
            sigmoid_f := 1689;
        ELSIF x = 3175 THEN
            sigmoid_f := 1689;
        ELSIF x = 3176 THEN
            sigmoid_f := 1689;
        ELSIF x = 3177 THEN
            sigmoid_f := 1689;
        ELSIF x = 3178 THEN
            sigmoid_f := 1690;
        ELSIF x = 3179 THEN
            sigmoid_f := 1690;
        ELSIF x = 3180 THEN
            sigmoid_f := 1690;
        ELSIF x = 3181 THEN
            sigmoid_f := 1690;
        ELSIF x = 3182 THEN
            sigmoid_f := 1690;
        ELSIF x = 3183 THEN
            sigmoid_f := 1690;
        ELSIF x = 3184 THEN
            sigmoid_f := 1690;
        ELSIF x = 3185 THEN
            sigmoid_f := 1691;
        ELSIF x = 3186 THEN
            sigmoid_f := 1691;
        ELSIF x = 3187 THEN
            sigmoid_f := 1691;
        ELSIF x = 3188 THEN
            sigmoid_f := 1691;
        ELSIF x = 3189 THEN
            sigmoid_f := 1691;
        ELSIF x = 3190 THEN
            sigmoid_f := 1691;
        ELSIF x = 3191 THEN
            sigmoid_f := 1691;
        ELSIF x = 3192 THEN
            sigmoid_f := 1691;
        ELSIF x = 3193 THEN
            sigmoid_f := 1692;
        ELSIF x = 3194 THEN
            sigmoid_f := 1692;
        ELSIF x = 3195 THEN
            sigmoid_f := 1692;
        ELSIF x = 3196 THEN
            sigmoid_f := 1692;
        ELSIF x = 3197 THEN
            sigmoid_f := 1692;
        ELSIF x = 3198 THEN
            sigmoid_f := 1692;
        ELSIF x = 3199 THEN
            sigmoid_f := 1692;
        ELSIF x = 3200 THEN
            sigmoid_f := 1693;
        ELSIF x = 3201 THEN
            sigmoid_f := 1693;
        ELSIF x = 3202 THEN
            sigmoid_f := 1693;
        ELSIF x = 3203 THEN
            sigmoid_f := 1693;
        ELSIF x = 3204 THEN
            sigmoid_f := 1693;
        ELSIF x = 3205 THEN
            sigmoid_f := 1693;
        ELSIF x = 3206 THEN
            sigmoid_f := 1693;
        ELSIF x = 3207 THEN
            sigmoid_f := 1694;
        ELSIF x = 3208 THEN
            sigmoid_f := 1694;
        ELSIF x = 3209 THEN
            sigmoid_f := 1694;
        ELSIF x = 3210 THEN
            sigmoid_f := 1694;
        ELSIF x = 3211 THEN
            sigmoid_f := 1694;
        ELSIF x = 3212 THEN
            sigmoid_f := 1694;
        ELSIF x = 3213 THEN
            sigmoid_f := 1694;
        ELSIF x = 3214 THEN
            sigmoid_f := 1694;
        ELSIF x = 3215 THEN
            sigmoid_f := 1695;
        ELSIF x = 3216 THEN
            sigmoid_f := 1695;
        ELSIF x = 3217 THEN
            sigmoid_f := 1695;
        ELSIF x = 3218 THEN
            sigmoid_f := 1695;
        ELSIF x = 3219 THEN
            sigmoid_f := 1695;
        ELSIF x = 3220 THEN
            sigmoid_f := 1695;
        ELSIF x = 3221 THEN
            sigmoid_f := 1695;
        ELSIF x = 3222 THEN
            sigmoid_f := 1696;
        ELSIF x = 3223 THEN
            sigmoid_f := 1696;
        ELSIF x = 3224 THEN
            sigmoid_f := 1696;
        ELSIF x = 3225 THEN
            sigmoid_f := 1696;
        ELSIF x = 3226 THEN
            sigmoid_f := 1696;
        ELSIF x = 3227 THEN
            sigmoid_f := 1696;
        ELSIF x = 3228 THEN
            sigmoid_f := 1696;
        ELSIF x = 3229 THEN
            sigmoid_f := 1697;
        ELSIF x = 3230 THEN
            sigmoid_f := 1697;
        ELSIF x = 3231 THEN
            sigmoid_f := 1697;
        ELSIF x = 3232 THEN
            sigmoid_f := 1697;
        ELSIF x = 3233 THEN
            sigmoid_f := 1697;
        ELSIF x = 3234 THEN
            sigmoid_f := 1697;
        ELSIF x = 3235 THEN
            sigmoid_f := 1697;
        ELSIF x = 3236 THEN
            sigmoid_f := 1698;
        ELSIF x = 3237 THEN
            sigmoid_f := 1698;
        ELSIF x = 3238 THEN
            sigmoid_f := 1698;
        ELSIF x = 3239 THEN
            sigmoid_f := 1698;
        ELSIF x = 3240 THEN
            sigmoid_f := 1698;
        ELSIF x = 3241 THEN
            sigmoid_f := 1698;
        ELSIF x = 3242 THEN
            sigmoid_f := 1698;
        ELSIF x = 3243 THEN
            sigmoid_f := 1698;
        ELSIF x = 3244 THEN
            sigmoid_f := 1699;
        ELSIF x = 3245 THEN
            sigmoid_f := 1699;
        ELSIF x = 3246 THEN
            sigmoid_f := 1699;
        ELSIF x = 3247 THEN
            sigmoid_f := 1699;
        ELSIF x = 3248 THEN
            sigmoid_f := 1699;
        ELSIF x = 3249 THEN
            sigmoid_f := 1699;
        ELSIF x = 3250 THEN
            sigmoid_f := 1699;
        ELSIF x = 3251 THEN
            sigmoid_f := 1700;
        ELSIF x = 3252 THEN
            sigmoid_f := 1700;
        ELSIF x = 3253 THEN
            sigmoid_f := 1700;
        ELSIF x = 3254 THEN
            sigmoid_f := 1700;
        ELSIF x = 3255 THEN
            sigmoid_f := 1700;
        ELSIF x = 3256 THEN
            sigmoid_f := 1700;
        ELSIF x = 3257 THEN
            sigmoid_f := 1700;
        ELSIF x = 3258 THEN
            sigmoid_f := 1701;
        ELSIF x = 3259 THEN
            sigmoid_f := 1701;
        ELSIF x = 3260 THEN
            sigmoid_f := 1701;
        ELSIF x = 3261 THEN
            sigmoid_f := 1701;
        ELSIF x = 3262 THEN
            sigmoid_f := 1701;
        ELSIF x = 3263 THEN
            sigmoid_f := 1701;
        ELSIF x = 3264 THEN
            sigmoid_f := 1701;
        ELSIF x = 3265 THEN
            sigmoid_f := 1701;
        ELSIF x = 3266 THEN
            sigmoid_f := 1702;
        ELSIF x = 3267 THEN
            sigmoid_f := 1702;
        ELSIF x = 3268 THEN
            sigmoid_f := 1702;
        ELSIF x = 3269 THEN
            sigmoid_f := 1702;
        ELSIF x = 3270 THEN
            sigmoid_f := 1702;
        ELSIF x = 3271 THEN
            sigmoid_f := 1702;
        ELSIF x = 3272 THEN
            sigmoid_f := 1702;
        ELSIF x = 3273 THEN
            sigmoid_f := 1703;
        ELSIF x = 3274 THEN
            sigmoid_f := 1703;
        ELSIF x = 3275 THEN
            sigmoid_f := 1703;
        ELSIF x = 3276 THEN
            sigmoid_f := 1703;
        ELSIF x = 3277 THEN
            sigmoid_f := 1703;
        ELSIF x = 3278 THEN
            sigmoid_f := 1703;
        ELSIF x = 3279 THEN
            sigmoid_f := 1703;
        ELSIF x = 3280 THEN
            sigmoid_f := 1704;
        ELSIF x = 3281 THEN
            sigmoid_f := 1704;
        ELSIF x = 3282 THEN
            sigmoid_f := 1704;
        ELSIF x = 3283 THEN
            sigmoid_f := 1704;
        ELSIF x = 3284 THEN
            sigmoid_f := 1704;
        ELSIF x = 3285 THEN
            sigmoid_f := 1704;
        ELSIF x = 3286 THEN
            sigmoid_f := 1704;
        ELSIF x = 3287 THEN
            sigmoid_f := 1704;
        ELSIF x = 3288 THEN
            sigmoid_f := 1705;
        ELSIF x = 3289 THEN
            sigmoid_f := 1705;
        ELSIF x = 3290 THEN
            sigmoid_f := 1705;
        ELSIF x = 3291 THEN
            sigmoid_f := 1705;
        ELSIF x = 3292 THEN
            sigmoid_f := 1705;
        ELSIF x = 3293 THEN
            sigmoid_f := 1705;
        ELSIF x = 3294 THEN
            sigmoid_f := 1705;
        ELSIF x = 3295 THEN
            sigmoid_f := 1706;
        ELSIF x = 3296 THEN
            sigmoid_f := 1706;
        ELSIF x = 3297 THEN
            sigmoid_f := 1706;
        ELSIF x = 3298 THEN
            sigmoid_f := 1706;
        ELSIF x = 3299 THEN
            sigmoid_f := 1706;
        ELSIF x = 3300 THEN
            sigmoid_f := 1706;
        ELSIF x = 3301 THEN
            sigmoid_f := 1706;
        ELSIF x = 3302 THEN
            sigmoid_f := 1707;
        ELSIF x = 3303 THEN
            sigmoid_f := 1707;
        ELSIF x = 3304 THEN
            sigmoid_f := 1707;
        ELSIF x = 3305 THEN
            sigmoid_f := 1707;
        ELSIF x = 3306 THEN
            sigmoid_f := 1707;
        ELSIF x = 3307 THEN
            sigmoid_f := 1707;
        ELSIF x = 3308 THEN
            sigmoid_f := 1707;
        ELSIF x = 3309 THEN
            sigmoid_f := 1708;
        ELSIF x = 3310 THEN
            sigmoid_f := 1708;
        ELSIF x = 3311 THEN
            sigmoid_f := 1708;
        ELSIF x = 3312 THEN
            sigmoid_f := 1708;
        ELSIF x = 3313 THEN
            sigmoid_f := 1708;
        ELSIF x = 3314 THEN
            sigmoid_f := 1708;
        ELSIF x = 3315 THEN
            sigmoid_f := 1708;
        ELSIF x = 3316 THEN
            sigmoid_f := 1708;
        ELSIF x = 3317 THEN
            sigmoid_f := 1709;
        ELSIF x = 3318 THEN
            sigmoid_f := 1709;
        ELSIF x = 3319 THEN
            sigmoid_f := 1709;
        ELSIF x = 3320 THEN
            sigmoid_f := 1709;
        ELSIF x = 3321 THEN
            sigmoid_f := 1709;
        ELSIF x = 3322 THEN
            sigmoid_f := 1709;
        ELSIF x = 3323 THEN
            sigmoid_f := 1709;
        ELSIF x = 3324 THEN
            sigmoid_f := 1710;
        ELSIF x = 3325 THEN
            sigmoid_f := 1710;
        ELSIF x = 3326 THEN
            sigmoid_f := 1710;
        ELSIF x = 3327 THEN
            sigmoid_f := 1710;
        ELSIF x = 3328 THEN
            sigmoid_f := 1710;
        ELSIF x = 3329 THEN
            sigmoid_f := 1710;
        ELSIF x = 3330 THEN
            sigmoid_f := 1710;
        ELSIF x = 3331 THEN
            sigmoid_f := 1711;
        ELSIF x = 3332 THEN
            sigmoid_f := 1711;
        ELSIF x = 3333 THEN
            sigmoid_f := 1711;
        ELSIF x = 3334 THEN
            sigmoid_f := 1711;
        ELSIF x = 3335 THEN
            sigmoid_f := 1711;
        ELSIF x = 3336 THEN
            sigmoid_f := 1711;
        ELSIF x = 3337 THEN
            sigmoid_f := 1711;
        ELSIF x = 3338 THEN
            sigmoid_f := 1711;
        ELSIF x = 3339 THEN
            sigmoid_f := 1712;
        ELSIF x = 3340 THEN
            sigmoid_f := 1712;
        ELSIF x = 3341 THEN
            sigmoid_f := 1712;
        ELSIF x = 3342 THEN
            sigmoid_f := 1712;
        ELSIF x = 3343 THEN
            sigmoid_f := 1712;
        ELSIF x = 3344 THEN
            sigmoid_f := 1712;
        ELSIF x = 3345 THEN
            sigmoid_f := 1712;
        ELSIF x = 3346 THEN
            sigmoid_f := 1713;
        ELSIF x = 3347 THEN
            sigmoid_f := 1713;
        ELSIF x = 3348 THEN
            sigmoid_f := 1713;
        ELSIF x = 3349 THEN
            sigmoid_f := 1713;
        ELSIF x = 3350 THEN
            sigmoid_f := 1713;
        ELSIF x = 3351 THEN
            sigmoid_f := 1713;
        ELSIF x = 3352 THEN
            sigmoid_f := 1713;
        ELSIF x = 3353 THEN
            sigmoid_f := 1714;
        ELSIF x = 3354 THEN
            sigmoid_f := 1714;
        ELSIF x = 3355 THEN
            sigmoid_f := 1714;
        ELSIF x = 3356 THEN
            sigmoid_f := 1714;
        ELSIF x = 3357 THEN
            sigmoid_f := 1714;
        ELSIF x = 3358 THEN
            sigmoid_f := 1714;
        ELSIF x = 3359 THEN
            sigmoid_f := 1714;
        ELSIF x = 3360 THEN
            sigmoid_f := 1715;
        ELSIF x = 3361 THEN
            sigmoid_f := 1715;
        ELSIF x = 3362 THEN
            sigmoid_f := 1715;
        ELSIF x = 3363 THEN
            sigmoid_f := 1715;
        ELSIF x = 3364 THEN
            sigmoid_f := 1715;
        ELSIF x = 3365 THEN
            sigmoid_f := 1715;
        ELSIF x = 3366 THEN
            sigmoid_f := 1715;
        ELSIF x = 3367 THEN
            sigmoid_f := 1715;
        ELSIF x = 3368 THEN
            sigmoid_f := 1716;
        ELSIF x = 3369 THEN
            sigmoid_f := 1716;
        ELSIF x = 3370 THEN
            sigmoid_f := 1716;
        ELSIF x = 3371 THEN
            sigmoid_f := 1716;
        ELSIF x = 3372 THEN
            sigmoid_f := 1716;
        ELSIF x = 3373 THEN
            sigmoid_f := 1716;
        ELSIF x = 3374 THEN
            sigmoid_f := 1716;
        ELSIF x = 3375 THEN
            sigmoid_f := 1717;
        ELSIF x = 3376 THEN
            sigmoid_f := 1717;
        ELSIF x = 3377 THEN
            sigmoid_f := 1717;
        ELSIF x = 3378 THEN
            sigmoid_f := 1717;
        ELSIF x = 3379 THEN
            sigmoid_f := 1717;
        ELSIF x = 3380 THEN
            sigmoid_f := 1717;
        ELSIF x = 3381 THEN
            sigmoid_f := 1717;
        ELSIF x = 3382 THEN
            sigmoid_f := 1718;
        ELSIF x = 3383 THEN
            sigmoid_f := 1718;
        ELSIF x = 3384 THEN
            sigmoid_f := 1718;
        ELSIF x = 3385 THEN
            sigmoid_f := 1718;
        ELSIF x = 3386 THEN
            sigmoid_f := 1718;
        ELSIF x = 3387 THEN
            sigmoid_f := 1718;
        ELSIF x = 3388 THEN
            sigmoid_f := 1718;
        ELSIF x = 3389 THEN
            sigmoid_f := 1718;
        ELSIF x = 3390 THEN
            sigmoid_f := 1719;
        ELSIF x = 3391 THEN
            sigmoid_f := 1719;
        ELSIF x = 3392 THEN
            sigmoid_f := 1719;
        ELSIF x = 3393 THEN
            sigmoid_f := 1719;
        ELSIF x = 3394 THEN
            sigmoid_f := 1719;
        ELSIF x = 3395 THEN
            sigmoid_f := 1719;
        ELSIF x = 3396 THEN
            sigmoid_f := 1719;
        ELSIF x = 3397 THEN
            sigmoid_f := 1720;
        ELSIF x = 3398 THEN
            sigmoid_f := 1720;
        ELSIF x = 3399 THEN
            sigmoid_f := 1720;
        ELSIF x = 3400 THEN
            sigmoid_f := 1720;
        ELSIF x = 3401 THEN
            sigmoid_f := 1720;
        ELSIF x = 3402 THEN
            sigmoid_f := 1720;
        ELSIF x = 3403 THEN
            sigmoid_f := 1720;
        ELSIF x = 3404 THEN
            sigmoid_f := 1721;
        ELSIF x = 3405 THEN
            sigmoid_f := 1721;
        ELSIF x = 3406 THEN
            sigmoid_f := 1721;
        ELSIF x = 3407 THEN
            sigmoid_f := 1721;
        ELSIF x = 3408 THEN
            sigmoid_f := 1721;
        ELSIF x = 3409 THEN
            sigmoid_f := 1721;
        ELSIF x = 3410 THEN
            sigmoid_f := 1721;
        ELSIF x = 3411 THEN
            sigmoid_f := 1722;
        ELSIF x = 3412 THEN
            sigmoid_f := 1722;
        ELSIF x = 3413 THEN
            sigmoid_f := 1722;
        ELSIF x = 3414 THEN
            sigmoid_f := 1722;
        ELSIF x = 3415 THEN
            sigmoid_f := 1722;
        ELSIF x = 3416 THEN
            sigmoid_f := 1722;
        ELSIF x = 3417 THEN
            sigmoid_f := 1722;
        ELSIF x = 3418 THEN
            sigmoid_f := 1722;
        ELSIF x = 3419 THEN
            sigmoid_f := 1723;
        ELSIF x = 3420 THEN
            sigmoid_f := 1723;
        ELSIF x = 3421 THEN
            sigmoid_f := 1723;
        ELSIF x = 3422 THEN
            sigmoid_f := 1723;
        ELSIF x = 3423 THEN
            sigmoid_f := 1723;
        ELSIF x = 3424 THEN
            sigmoid_f := 1723;
        ELSIF x = 3425 THEN
            sigmoid_f := 1723;
        ELSIF x = 3426 THEN
            sigmoid_f := 1724;
        ELSIF x = 3427 THEN
            sigmoid_f := 1724;
        ELSIF x = 3428 THEN
            sigmoid_f := 1724;
        ELSIF x = 3429 THEN
            sigmoid_f := 1724;
        ELSIF x = 3430 THEN
            sigmoid_f := 1724;
        ELSIF x = 3431 THEN
            sigmoid_f := 1724;
        ELSIF x = 3432 THEN
            sigmoid_f := 1724;
        ELSIF x = 3433 THEN
            sigmoid_f := 1725;
        ELSIF x = 3434 THEN
            sigmoid_f := 1725;
        ELSIF x = 3435 THEN
            sigmoid_f := 1725;
        ELSIF x = 3436 THEN
            sigmoid_f := 1725;
        ELSIF x = 3437 THEN
            sigmoid_f := 1725;
        ELSIF x = 3438 THEN
            sigmoid_f := 1725;
        ELSIF x = 3439 THEN
            sigmoid_f := 1725;
        ELSIF x = 3440 THEN
            sigmoid_f := 1725;
        ELSIF x = 3441 THEN
            sigmoid_f := 1726;
        ELSIF x = 3442 THEN
            sigmoid_f := 1726;
        ELSIF x = 3443 THEN
            sigmoid_f := 1726;
        ELSIF x = 3444 THEN
            sigmoid_f := 1726;
        ELSIF x = 3445 THEN
            sigmoid_f := 1726;
        ELSIF x = 3446 THEN
            sigmoid_f := 1726;
        ELSIF x = 3447 THEN
            sigmoid_f := 1726;
        ELSIF x = 3448 THEN
            sigmoid_f := 1727;
        ELSIF x = 3449 THEN
            sigmoid_f := 1727;
        ELSIF x = 3450 THEN
            sigmoid_f := 1727;
        ELSIF x = 3451 THEN
            sigmoid_f := 1727;
        ELSIF x = 3452 THEN
            sigmoid_f := 1727;
        ELSIF x = 3453 THEN
            sigmoid_f := 1727;
        ELSIF x = 3454 THEN
            sigmoid_f := 1727;
        ELSIF x = 3455 THEN
            sigmoid_f := 1728;
        ELSIF x = 3456 THEN
            sigmoid_f := 1728;
        ELSIF x = 3457 THEN
            sigmoid_f := 1728;
        ELSIF x = 3458 THEN
            sigmoid_f := 1728;
        ELSIF x = 3459 THEN
            sigmoid_f := 1728;
        ELSIF x = 3460 THEN
            sigmoid_f := 1728;
        ELSIF x = 3461 THEN
            sigmoid_f := 1728;
        ELSIF x = 3462 THEN
            sigmoid_f := 1729;
        ELSIF x = 3463 THEN
            sigmoid_f := 1729;
        ELSIF x = 3464 THEN
            sigmoid_f := 1729;
        ELSIF x = 3465 THEN
            sigmoid_f := 1729;
        ELSIF x = 3466 THEN
            sigmoid_f := 1729;
        ELSIF x = 3467 THEN
            sigmoid_f := 1729;
        ELSIF x = 3468 THEN
            sigmoid_f := 1729;
        ELSIF x = 3469 THEN
            sigmoid_f := 1729;
        ELSIF x = 3470 THEN
            sigmoid_f := 1730;
        ELSIF x = 3471 THEN
            sigmoid_f := 1730;
        ELSIF x = 3472 THEN
            sigmoid_f := 1730;
        ELSIF x = 3473 THEN
            sigmoid_f := 1730;
        ELSIF x = 3474 THEN
            sigmoid_f := 1730;
        ELSIF x = 3475 THEN
            sigmoid_f := 1730;
        ELSIF x = 3476 THEN
            sigmoid_f := 1730;
        ELSIF x = 3477 THEN
            sigmoid_f := 1731;
        ELSIF x = 3478 THEN
            sigmoid_f := 1731;
        ELSIF x = 3479 THEN
            sigmoid_f := 1731;
        ELSIF x = 3480 THEN
            sigmoid_f := 1731;
        ELSIF x = 3481 THEN
            sigmoid_f := 1731;
        ELSIF x = 3482 THEN
            sigmoid_f := 1731;
        ELSIF x = 3483 THEN
            sigmoid_f := 1731;
        ELSIF x = 3484 THEN
            sigmoid_f := 1732;
        ELSIF x = 3485 THEN
            sigmoid_f := 1732;
        ELSIF x = 3486 THEN
            sigmoid_f := 1732;
        ELSIF x = 3487 THEN
            sigmoid_f := 1732;
        ELSIF x = 3488 THEN
            sigmoid_f := 1732;
        ELSIF x = 3489 THEN
            sigmoid_f := 1732;
        ELSIF x = 3490 THEN
            sigmoid_f := 1732;
        ELSIF x = 3491 THEN
            sigmoid_f := 1732;
        ELSIF x = 3492 THEN
            sigmoid_f := 1733;
        ELSIF x = 3493 THEN
            sigmoid_f := 1733;
        ELSIF x = 3494 THEN
            sigmoid_f := 1733;
        ELSIF x = 3495 THEN
            sigmoid_f := 1733;
        ELSIF x = 3496 THEN
            sigmoid_f := 1733;
        ELSIF x = 3497 THEN
            sigmoid_f := 1733;
        ELSIF x = 3498 THEN
            sigmoid_f := 1733;
        ELSIF x = 3499 THEN
            sigmoid_f := 1734;
        ELSIF x = 3500 THEN
            sigmoid_f := 1734;
        ELSIF x = 3501 THEN
            sigmoid_f := 1734;
        ELSIF x = 3502 THEN
            sigmoid_f := 1734;
        ELSIF x = 3503 THEN
            sigmoid_f := 1734;
        ELSIF x = 3504 THEN
            sigmoid_f := 1734;
        ELSIF x = 3505 THEN
            sigmoid_f := 1734;
        ELSIF x = 3506 THEN
            sigmoid_f := 1735;
        ELSIF x = 3507 THEN
            sigmoid_f := 1735;
        ELSIF x = 3508 THEN
            sigmoid_f := 1735;
        ELSIF x = 3509 THEN
            sigmoid_f := 1735;
        ELSIF x = 3510 THEN
            sigmoid_f := 1735;
        ELSIF x = 3511 THEN
            sigmoid_f := 1735;
        ELSIF x = 3512 THEN
            sigmoid_f := 1735;
        ELSIF x = 3513 THEN
            sigmoid_f := 1736;
        ELSIF x = 3514 THEN
            sigmoid_f := 1736;
        ELSIF x = 3515 THEN
            sigmoid_f := 1736;
        ELSIF x = 3516 THEN
            sigmoid_f := 1736;
        ELSIF x = 3517 THEN
            sigmoid_f := 1736;
        ELSIF x = 3518 THEN
            sigmoid_f := 1736;
        ELSIF x = 3519 THEN
            sigmoid_f := 1736;
        ELSIF x = 3520 THEN
            sigmoid_f := 1736;
        ELSIF x = 3521 THEN
            sigmoid_f := 1737;
        ELSIF x = 3522 THEN
            sigmoid_f := 1737;
        ELSIF x = 3523 THEN
            sigmoid_f := 1737;
        ELSIF x = 3524 THEN
            sigmoid_f := 1737;
        ELSIF x = 3525 THEN
            sigmoid_f := 1737;
        ELSIF x = 3526 THEN
            sigmoid_f := 1737;
        ELSIF x = 3527 THEN
            sigmoid_f := 1737;
        ELSIF x = 3528 THEN
            sigmoid_f := 1738;
        ELSIF x = 3529 THEN
            sigmoid_f := 1738;
        ELSIF x = 3530 THEN
            sigmoid_f := 1738;
        ELSIF x = 3531 THEN
            sigmoid_f := 1738;
        ELSIF x = 3532 THEN
            sigmoid_f := 1738;
        ELSIF x = 3533 THEN
            sigmoid_f := 1738;
        ELSIF x = 3534 THEN
            sigmoid_f := 1738;
        ELSIF x = 3535 THEN
            sigmoid_f := 1739;
        ELSIF x = 3536 THEN
            sigmoid_f := 1739;
        ELSIF x = 3537 THEN
            sigmoid_f := 1739;
        ELSIF x = 3538 THEN
            sigmoid_f := 1739;
        ELSIF x = 3539 THEN
            sigmoid_f := 1739;
        ELSIF x = 3540 THEN
            sigmoid_f := 1739;
        ELSIF x = 3541 THEN
            sigmoid_f := 1739;
        ELSIF x = 3542 THEN
            sigmoid_f := 1739;
        ELSIF x = 3543 THEN
            sigmoid_f := 1740;
        ELSIF x = 3544 THEN
            sigmoid_f := 1740;
        ELSIF x = 3545 THEN
            sigmoid_f := 1740;
        ELSIF x = 3546 THEN
            sigmoid_f := 1740;
        ELSIF x = 3547 THEN
            sigmoid_f := 1740;
        ELSIF x = 3548 THEN
            sigmoid_f := 1740;
        ELSIF x = 3549 THEN
            sigmoid_f := 1740;
        ELSIF x = 3550 THEN
            sigmoid_f := 1741;
        ELSIF x = 3551 THEN
            sigmoid_f := 1741;
        ELSIF x = 3552 THEN
            sigmoid_f := 1741;
        ELSIF x = 3553 THEN
            sigmoid_f := 1741;
        ELSIF x = 3554 THEN
            sigmoid_f := 1741;
        ELSIF x = 3555 THEN
            sigmoid_f := 1741;
        ELSIF x = 3556 THEN
            sigmoid_f := 1741;
        ELSIF x = 3557 THEN
            sigmoid_f := 1742;
        ELSIF x = 3558 THEN
            sigmoid_f := 1742;
        ELSIF x = 3559 THEN
            sigmoid_f := 1742;
        ELSIF x = 3560 THEN
            sigmoid_f := 1742;
        ELSIF x = 3561 THEN
            sigmoid_f := 1742;
        ELSIF x = 3562 THEN
            sigmoid_f := 1742;
        ELSIF x = 3563 THEN
            sigmoid_f := 1742;
        ELSIF x = 3564 THEN
            sigmoid_f := 1743;
        ELSIF x = 3565 THEN
            sigmoid_f := 1743;
        ELSIF x = 3566 THEN
            sigmoid_f := 1743;
        ELSIF x = 3567 THEN
            sigmoid_f := 1743;
        ELSIF x = 3568 THEN
            sigmoid_f := 1743;
        ELSIF x = 3569 THEN
            sigmoid_f := 1743;
        ELSIF x = 3570 THEN
            sigmoid_f := 1743;
        ELSIF x = 3571 THEN
            sigmoid_f := 1743;
        ELSIF x = 3572 THEN
            sigmoid_f := 1744;
        ELSIF x = 3573 THEN
            sigmoid_f := 1744;
        ELSIF x = 3574 THEN
            sigmoid_f := 1744;
        ELSIF x = 3575 THEN
            sigmoid_f := 1744;
        ELSIF x = 3576 THEN
            sigmoid_f := 1744;
        ELSIF x = 3577 THEN
            sigmoid_f := 1744;
        ELSIF x = 3578 THEN
            sigmoid_f := 1744;
        ELSIF x = 3579 THEN
            sigmoid_f := 1745;
        ELSIF x = 3580 THEN
            sigmoid_f := 1745;
        ELSIF x = 3581 THEN
            sigmoid_f := 1745;
        ELSIF x = 3582 THEN
            sigmoid_f := 1745;
        ELSIF x = 3583 THEN
            sigmoid_f := 1745;
        ELSIF x = 3584 THEN
            sigmoid_f := 1745;
        ELSIF x = 3585 THEN
            sigmoid_f := 1745;
        ELSIF x = 3586 THEN
            sigmoid_f := 1745;
        ELSIF x = 3587 THEN
            sigmoid_f := 1745;
        ELSIF x = 3588 THEN
            sigmoid_f := 1745;
        ELSIF x = 3589 THEN
            sigmoid_f := 1746;
        ELSIF x = 3590 THEN
            sigmoid_f := 1746;
        ELSIF x = 3591 THEN
            sigmoid_f := 1746;
        ELSIF x = 3592 THEN
            sigmoid_f := 1746;
        ELSIF x = 3593 THEN
            sigmoid_f := 1746;
        ELSIF x = 3594 THEN
            sigmoid_f := 1746;
        ELSIF x = 3595 THEN
            sigmoid_f := 1746;
        ELSIF x = 3596 THEN
            sigmoid_f := 1746;
        ELSIF x = 3597 THEN
            sigmoid_f := 1747;
        ELSIF x = 3598 THEN
            sigmoid_f := 1747;
        ELSIF x = 3599 THEN
            sigmoid_f := 1747;
        ELSIF x = 3600 THEN
            sigmoid_f := 1747;
        ELSIF x = 3601 THEN
            sigmoid_f := 1747;
        ELSIF x = 3602 THEN
            sigmoid_f := 1747;
        ELSIF x = 3603 THEN
            sigmoid_f := 1747;
        ELSIF x = 3604 THEN
            sigmoid_f := 1747;
        ELSIF x = 3605 THEN
            sigmoid_f := 1747;
        ELSIF x = 3606 THEN
            sigmoid_f := 1748;
        ELSIF x = 3607 THEN
            sigmoid_f := 1748;
        ELSIF x = 3608 THEN
            sigmoid_f := 1748;
        ELSIF x = 3609 THEN
            sigmoid_f := 1748;
        ELSIF x = 3610 THEN
            sigmoid_f := 1748;
        ELSIF x = 3611 THEN
            sigmoid_f := 1748;
        ELSIF x = 3612 THEN
            sigmoid_f := 1748;
        ELSIF x = 3613 THEN
            sigmoid_f := 1748;
        ELSIF x = 3614 THEN
            sigmoid_f := 1748;
        ELSIF x = 3615 THEN
            sigmoid_f := 1749;
        ELSIF x = 3616 THEN
            sigmoid_f := 1749;
        ELSIF x = 3617 THEN
            sigmoid_f := 1749;
        ELSIF x = 3618 THEN
            sigmoid_f := 1749;
        ELSIF x = 3619 THEN
            sigmoid_f := 1749;
        ELSIF x = 3620 THEN
            sigmoid_f := 1749;
        ELSIF x = 3621 THEN
            sigmoid_f := 1749;
        ELSIF x = 3622 THEN
            sigmoid_f := 1749;
        ELSIF x = 3623 THEN
            sigmoid_f := 1750;
        ELSIF x = 3624 THEN
            sigmoid_f := 1750;
        ELSIF x = 3625 THEN
            sigmoid_f := 1750;
        ELSIF x = 3626 THEN
            sigmoid_f := 1750;
        ELSIF x = 3627 THEN
            sigmoid_f := 1750;
        ELSIF x = 3628 THEN
            sigmoid_f := 1750;
        ELSIF x = 3629 THEN
            sigmoid_f := 1750;
        ELSIF x = 3630 THEN
            sigmoid_f := 1750;
        ELSIF x = 3631 THEN
            sigmoid_f := 1750;
        ELSIF x = 3632 THEN
            sigmoid_f := 1751;
        ELSIF x = 3633 THEN
            sigmoid_f := 1751;
        ELSIF x = 3634 THEN
            sigmoid_f := 1751;
        ELSIF x = 3635 THEN
            sigmoid_f := 1751;
        ELSIF x = 3636 THEN
            sigmoid_f := 1751;
        ELSIF x = 3637 THEN
            sigmoid_f := 1751;
        ELSIF x = 3638 THEN
            sigmoid_f := 1751;
        ELSIF x = 3639 THEN
            sigmoid_f := 1751;
        ELSIF x = 3640 THEN
            sigmoid_f := 1752;
        ELSIF x = 3641 THEN
            sigmoid_f := 1752;
        ELSIF x = 3642 THEN
            sigmoid_f := 1752;
        ELSIF x = 3643 THEN
            sigmoid_f := 1752;
        ELSIF x = 3644 THEN
            sigmoid_f := 1752;
        ELSIF x = 3645 THEN
            sigmoid_f := 1752;
        ELSIF x = 3646 THEN
            sigmoid_f := 1752;
        ELSIF x = 3647 THEN
            sigmoid_f := 1752;
        ELSIF x = 3648 THEN
            sigmoid_f := 1752;
        ELSIF x = 3649 THEN
            sigmoid_f := 1753;
        ELSIF x = 3650 THEN
            sigmoid_f := 1753;
        ELSIF x = 3651 THEN
            sigmoid_f := 1753;
        ELSIF x = 3652 THEN
            sigmoid_f := 1753;
        ELSIF x = 3653 THEN
            sigmoid_f := 1753;
        ELSIF x = 3654 THEN
            sigmoid_f := 1753;
        ELSIF x = 3655 THEN
            sigmoid_f := 1753;
        ELSIF x = 3656 THEN
            sigmoid_f := 1753;
        ELSIF x = 3657 THEN
            sigmoid_f := 1753;
        ELSIF x = 3658 THEN
            sigmoid_f := 1754;
        ELSIF x = 3659 THEN
            sigmoid_f := 1754;
        ELSIF x = 3660 THEN
            sigmoid_f := 1754;
        ELSIF x = 3661 THEN
            sigmoid_f := 1754;
        ELSIF x = 3662 THEN
            sigmoid_f := 1754;
        ELSIF x = 3663 THEN
            sigmoid_f := 1754;
        ELSIF x = 3664 THEN
            sigmoid_f := 1754;
        ELSIF x = 3665 THEN
            sigmoid_f := 1754;
        ELSIF x = 3666 THEN
            sigmoid_f := 1755;
        ELSIF x = 3667 THEN
            sigmoid_f := 1755;
        ELSIF x = 3668 THEN
            sigmoid_f := 1755;
        ELSIF x = 3669 THEN
            sigmoid_f := 1755;
        ELSIF x = 3670 THEN
            sigmoid_f := 1755;
        ELSIF x = 3671 THEN
            sigmoid_f := 1755;
        ELSIF x = 3672 THEN
            sigmoid_f := 1755;
        ELSIF x = 3673 THEN
            sigmoid_f := 1755;
        ELSIF x = 3674 THEN
            sigmoid_f := 1755;
        ELSIF x = 3675 THEN
            sigmoid_f := 1756;
        ELSIF x = 3676 THEN
            sigmoid_f := 1756;
        ELSIF x = 3677 THEN
            sigmoid_f := 1756;
        ELSIF x = 3678 THEN
            sigmoid_f := 1756;
        ELSIF x = 3679 THEN
            sigmoid_f := 1756;
        ELSIF x = 3680 THEN
            sigmoid_f := 1756;
        ELSIF x = 3681 THEN
            sigmoid_f := 1756;
        ELSIF x = 3682 THEN
            sigmoid_f := 1756;
        ELSIF x = 3683 THEN
            sigmoid_f := 1757;
        ELSIF x = 3684 THEN
            sigmoid_f := 1757;
        ELSIF x = 3685 THEN
            sigmoid_f := 1757;
        ELSIF x = 3686 THEN
            sigmoid_f := 1757;
        ELSIF x = 3687 THEN
            sigmoid_f := 1757;
        ELSIF x = 3688 THEN
            sigmoid_f := 1757;
        ELSIF x = 3689 THEN
            sigmoid_f := 1757;
        ELSIF x = 3690 THEN
            sigmoid_f := 1757;
        ELSIF x = 3691 THEN
            sigmoid_f := 1757;
        ELSIF x = 3692 THEN
            sigmoid_f := 1758;
        ELSIF x = 3693 THEN
            sigmoid_f := 1758;
        ELSIF x = 3694 THEN
            sigmoid_f := 1758;
        ELSIF x = 3695 THEN
            sigmoid_f := 1758;
        ELSIF x = 3696 THEN
            sigmoid_f := 1758;
        ELSIF x = 3697 THEN
            sigmoid_f := 1758;
        ELSIF x = 3698 THEN
            sigmoid_f := 1758;
        ELSIF x = 3699 THEN
            sigmoid_f := 1758;
        ELSIF x = 3700 THEN
            sigmoid_f := 1758;
        ELSIF x = 3701 THEN
            sigmoid_f := 1759;
        ELSIF x = 3702 THEN
            sigmoid_f := 1759;
        ELSIF x = 3703 THEN
            sigmoid_f := 1759;
        ELSIF x = 3704 THEN
            sigmoid_f := 1759;
        ELSIF x = 3705 THEN
            sigmoid_f := 1759;
        ELSIF x = 3706 THEN
            sigmoid_f := 1759;
        ELSIF x = 3707 THEN
            sigmoid_f := 1759;
        ELSIF x = 3708 THEN
            sigmoid_f := 1759;
        ELSIF x = 3709 THEN
            sigmoid_f := 1760;
        ELSIF x = 3710 THEN
            sigmoid_f := 1760;
        ELSIF x = 3711 THEN
            sigmoid_f := 1760;
        ELSIF x = 3712 THEN
            sigmoid_f := 1760;
        ELSIF x = 3713 THEN
            sigmoid_f := 1760;
        ELSIF x = 3714 THEN
            sigmoid_f := 1760;
        ELSIF x = 3715 THEN
            sigmoid_f := 1760;
        ELSIF x = 3716 THEN
            sigmoid_f := 1760;
        ELSIF x = 3717 THEN
            sigmoid_f := 1760;
        ELSIF x = 3718 THEN
            sigmoid_f := 1761;
        ELSIF x = 3719 THEN
            sigmoid_f := 1761;
        ELSIF x = 3720 THEN
            sigmoid_f := 1761;
        ELSIF x = 3721 THEN
            sigmoid_f := 1761;
        ELSIF x = 3722 THEN
            sigmoid_f := 1761;
        ELSIF x = 3723 THEN
            sigmoid_f := 1761;
        ELSIF x = 3724 THEN
            sigmoid_f := 1761;
        ELSIF x = 3725 THEN
            sigmoid_f := 1761;
        ELSIF x = 3726 THEN
            sigmoid_f := 1762;
        ELSIF x = 3727 THEN
            sigmoid_f := 1762;
        ELSIF x = 3728 THEN
            sigmoid_f := 1762;
        ELSIF x = 3729 THEN
            sigmoid_f := 1762;
        ELSIF x = 3730 THEN
            sigmoid_f := 1762;
        ELSIF x = 3731 THEN
            sigmoid_f := 1762;
        ELSIF x = 3732 THEN
            sigmoid_f := 1762;
        ELSIF x = 3733 THEN
            sigmoid_f := 1762;
        ELSIF x = 3734 THEN
            sigmoid_f := 1762;
        ELSIF x = 3735 THEN
            sigmoid_f := 1763;
        ELSIF x = 3736 THEN
            sigmoid_f := 1763;
        ELSIF x = 3737 THEN
            sigmoid_f := 1763;
        ELSIF x = 3738 THEN
            sigmoid_f := 1763;
        ELSIF x = 3739 THEN
            sigmoid_f := 1763;
        ELSIF x = 3740 THEN
            sigmoid_f := 1763;
        ELSIF x = 3741 THEN
            sigmoid_f := 1763;
        ELSIF x = 3742 THEN
            sigmoid_f := 1763;
        ELSIF x = 3743 THEN
            sigmoid_f := 1763;
        ELSIF x = 3744 THEN
            sigmoid_f := 1764;
        ELSIF x = 3745 THEN
            sigmoid_f := 1764;
        ELSIF x = 3746 THEN
            sigmoid_f := 1764;
        ELSIF x = 3747 THEN
            sigmoid_f := 1764;
        ELSIF x = 3748 THEN
            sigmoid_f := 1764;
        ELSIF x = 3749 THEN
            sigmoid_f := 1764;
        ELSIF x = 3750 THEN
            sigmoid_f := 1764;
        ELSIF x = 3751 THEN
            sigmoid_f := 1764;
        ELSIF x = 3752 THEN
            sigmoid_f := 1765;
        ELSIF x = 3753 THEN
            sigmoid_f := 1765;
        ELSIF x = 3754 THEN
            sigmoid_f := 1765;
        ELSIF x = 3755 THEN
            sigmoid_f := 1765;
        ELSIF x = 3756 THEN
            sigmoid_f := 1765;
        ELSIF x = 3757 THEN
            sigmoid_f := 1765;
        ELSIF x = 3758 THEN
            sigmoid_f := 1765;
        ELSIF x = 3759 THEN
            sigmoid_f := 1765;
        ELSIF x = 3760 THEN
            sigmoid_f := 1765;
        ELSIF x = 3761 THEN
            sigmoid_f := 1766;
        ELSIF x = 3762 THEN
            sigmoid_f := 1766;
        ELSIF x = 3763 THEN
            sigmoid_f := 1766;
        ELSIF x = 3764 THEN
            sigmoid_f := 1766;
        ELSIF x = 3765 THEN
            sigmoid_f := 1766;
        ELSIF x = 3766 THEN
            sigmoid_f := 1766;
        ELSIF x = 3767 THEN
            sigmoid_f := 1766;
        ELSIF x = 3768 THEN
            sigmoid_f := 1766;
        ELSIF x = 3769 THEN
            sigmoid_f := 1766;
        ELSIF x = 3770 THEN
            sigmoid_f := 1767;
        ELSIF x = 3771 THEN
            sigmoid_f := 1767;
        ELSIF x = 3772 THEN
            sigmoid_f := 1767;
        ELSIF x = 3773 THEN
            sigmoid_f := 1767;
        ELSIF x = 3774 THEN
            sigmoid_f := 1767;
        ELSIF x = 3775 THEN
            sigmoid_f := 1767;
        ELSIF x = 3776 THEN
            sigmoid_f := 1767;
        ELSIF x = 3777 THEN
            sigmoid_f := 1767;
        ELSIF x = 3778 THEN
            sigmoid_f := 1768;
        ELSIF x = 3779 THEN
            sigmoid_f := 1768;
        ELSIF x = 3780 THEN
            sigmoid_f := 1768;
        ELSIF x = 3781 THEN
            sigmoid_f := 1768;
        ELSIF x = 3782 THEN
            sigmoid_f := 1768;
        ELSIF x = 3783 THEN
            sigmoid_f := 1768;
        ELSIF x = 3784 THEN
            sigmoid_f := 1768;
        ELSIF x = 3785 THEN
            sigmoid_f := 1768;
        ELSIF x = 3786 THEN
            sigmoid_f := 1768;
        ELSIF x = 3787 THEN
            sigmoid_f := 1769;
        ELSIF x = 3788 THEN
            sigmoid_f := 1769;
        ELSIF x = 3789 THEN
            sigmoid_f := 1769;
        ELSIF x = 3790 THEN
            sigmoid_f := 1769;
        ELSIF x = 3791 THEN
            sigmoid_f := 1769;
        ELSIF x = 3792 THEN
            sigmoid_f := 1769;
        ELSIF x = 3793 THEN
            sigmoid_f := 1769;
        ELSIF x = 3794 THEN
            sigmoid_f := 1769;
        ELSIF x = 3795 THEN
            sigmoid_f := 1770;
        ELSIF x = 3796 THEN
            sigmoid_f := 1770;
        ELSIF x = 3797 THEN
            sigmoid_f := 1770;
        ELSIF x = 3798 THEN
            sigmoid_f := 1770;
        ELSIF x = 3799 THEN
            sigmoid_f := 1770;
        ELSIF x = 3800 THEN
            sigmoid_f := 1770;
        ELSIF x = 3801 THEN
            sigmoid_f := 1770;
        ELSIF x = 3802 THEN
            sigmoid_f := 1770;
        ELSIF x = 3803 THEN
            sigmoid_f := 1770;
        ELSIF x = 3804 THEN
            sigmoid_f := 1771;
        ELSIF x = 3805 THEN
            sigmoid_f := 1771;
        ELSIF x = 3806 THEN
            sigmoid_f := 1771;
        ELSIF x = 3807 THEN
            sigmoid_f := 1771;
        ELSIF x = 3808 THEN
            sigmoid_f := 1771;
        ELSIF x = 3809 THEN
            sigmoid_f := 1771;
        ELSIF x = 3810 THEN
            sigmoid_f := 1771;
        ELSIF x = 3811 THEN
            sigmoid_f := 1771;
        ELSIF x = 3812 THEN
            sigmoid_f := 1771;
        ELSIF x = 3813 THEN
            sigmoid_f := 1772;
        ELSIF x = 3814 THEN
            sigmoid_f := 1772;
        ELSIF x = 3815 THEN
            sigmoid_f := 1772;
        ELSIF x = 3816 THEN
            sigmoid_f := 1772;
        ELSIF x = 3817 THEN
            sigmoid_f := 1772;
        ELSIF x = 3818 THEN
            sigmoid_f := 1772;
        ELSIF x = 3819 THEN
            sigmoid_f := 1772;
        ELSIF x = 3820 THEN
            sigmoid_f := 1772;
        ELSIF x = 3821 THEN
            sigmoid_f := 1773;
        ELSIF x = 3822 THEN
            sigmoid_f := 1773;
        ELSIF x = 3823 THEN
            sigmoid_f := 1773;
        ELSIF x = 3824 THEN
            sigmoid_f := 1773;
        ELSIF x = 3825 THEN
            sigmoid_f := 1773;
        ELSIF x = 3826 THEN
            sigmoid_f := 1773;
        ELSIF x = 3827 THEN
            sigmoid_f := 1773;
        ELSIF x = 3828 THEN
            sigmoid_f := 1773;
        ELSIF x = 3829 THEN
            sigmoid_f := 1773;
        ELSIF x = 3830 THEN
            sigmoid_f := 1774;
        ELSIF x = 3831 THEN
            sigmoid_f := 1774;
        ELSIF x = 3832 THEN
            sigmoid_f := 1774;
        ELSIF x = 3833 THEN
            sigmoid_f := 1774;
        ELSIF x = 3834 THEN
            sigmoid_f := 1774;
        ELSIF x = 3835 THEN
            sigmoid_f := 1774;
        ELSIF x = 3836 THEN
            sigmoid_f := 1774;
        ELSIF x = 3837 THEN
            sigmoid_f := 1774;
        ELSIF x = 3838 THEN
            sigmoid_f := 1775;
        ELSIF x = 3839 THEN
            sigmoid_f := 1775;
        ELSIF x = 3840 THEN
            sigmoid_f := 1775;
        ELSIF x = 3841 THEN
            sigmoid_f := 1775;
        ELSIF x = 3842 THEN
            sigmoid_f := 1775;
        ELSIF x = 3843 THEN
            sigmoid_f := 1775;
        ELSIF x = 3844 THEN
            sigmoid_f := 1775;
        ELSIF x = 3845 THEN
            sigmoid_f := 1775;
        ELSIF x = 3846 THEN
            sigmoid_f := 1775;
        ELSIF x = 3847 THEN
            sigmoid_f := 1776;
        ELSIF x = 3848 THEN
            sigmoid_f := 1776;
        ELSIF x = 3849 THEN
            sigmoid_f := 1776;
        ELSIF x = 3850 THEN
            sigmoid_f := 1776;
        ELSIF x = 3851 THEN
            sigmoid_f := 1776;
        ELSIF x = 3852 THEN
            sigmoid_f := 1776;
        ELSIF x = 3853 THEN
            sigmoid_f := 1776;
        ELSIF x = 3854 THEN
            sigmoid_f := 1776;
        ELSIF x = 3855 THEN
            sigmoid_f := 1776;
        ELSIF x = 3856 THEN
            sigmoid_f := 1777;
        ELSIF x = 3857 THEN
            sigmoid_f := 1777;
        ELSIF x = 3858 THEN
            sigmoid_f := 1777;
        ELSIF x = 3859 THEN
            sigmoid_f := 1777;
        ELSIF x = 3860 THEN
            sigmoid_f := 1777;
        ELSIF x = 3861 THEN
            sigmoid_f := 1777;
        ELSIF x = 3862 THEN
            sigmoid_f := 1777;
        ELSIF x = 3863 THEN
            sigmoid_f := 1777;
        ELSIF x = 3864 THEN
            sigmoid_f := 1778;
        ELSIF x = 3865 THEN
            sigmoid_f := 1778;
        ELSIF x = 3866 THEN
            sigmoid_f := 1778;
        ELSIF x = 3867 THEN
            sigmoid_f := 1778;
        ELSIF x = 3868 THEN
            sigmoid_f := 1778;
        ELSIF x = 3869 THEN
            sigmoid_f := 1778;
        ELSIF x = 3870 THEN
            sigmoid_f := 1778;
        ELSIF x = 3871 THEN
            sigmoid_f := 1778;
        ELSIF x = 3872 THEN
            sigmoid_f := 1778;
        ELSIF x = 3873 THEN
            sigmoid_f := 1779;
        ELSIF x = 3874 THEN
            sigmoid_f := 1779;
        ELSIF x = 3875 THEN
            sigmoid_f := 1779;
        ELSIF x = 3876 THEN
            sigmoid_f := 1779;
        ELSIF x = 3877 THEN
            sigmoid_f := 1779;
        ELSIF x = 3878 THEN
            sigmoid_f := 1779;
        ELSIF x = 3879 THEN
            sigmoid_f := 1779;
        ELSIF x = 3880 THEN
            sigmoid_f := 1779;
        ELSIF x = 3881 THEN
            sigmoid_f := 1780;
        ELSIF x = 3882 THEN
            sigmoid_f := 1780;
        ELSIF x = 3883 THEN
            sigmoid_f := 1780;
        ELSIF x = 3884 THEN
            sigmoid_f := 1780;
        ELSIF x = 3885 THEN
            sigmoid_f := 1780;
        ELSIF x = 3886 THEN
            sigmoid_f := 1780;
        ELSIF x = 3887 THEN
            sigmoid_f := 1780;
        ELSIF x = 3888 THEN
            sigmoid_f := 1780;
        ELSIF x = 3889 THEN
            sigmoid_f := 1780;
        ELSIF x = 3890 THEN
            sigmoid_f := 1781;
        ELSIF x = 3891 THEN
            sigmoid_f := 1781;
        ELSIF x = 3892 THEN
            sigmoid_f := 1781;
        ELSIF x = 3893 THEN
            sigmoid_f := 1781;
        ELSIF x = 3894 THEN
            sigmoid_f := 1781;
        ELSIF x = 3895 THEN
            sigmoid_f := 1781;
        ELSIF x = 3896 THEN
            sigmoid_f := 1781;
        ELSIF x = 3897 THEN
            sigmoid_f := 1781;
        ELSIF x = 3898 THEN
            sigmoid_f := 1781;
        ELSIF x = 3899 THEN
            sigmoid_f := 1782;
        ELSIF x = 3900 THEN
            sigmoid_f := 1782;
        ELSIF x = 3901 THEN
            sigmoid_f := 1782;
        ELSIF x = 3902 THEN
            sigmoid_f := 1782;
        ELSIF x = 3903 THEN
            sigmoid_f := 1782;
        ELSIF x = 3904 THEN
            sigmoid_f := 1782;
        ELSIF x = 3905 THEN
            sigmoid_f := 1782;
        ELSIF x = 3906 THEN
            sigmoid_f := 1782;
        ELSIF x = 3907 THEN
            sigmoid_f := 1783;
        ELSIF x = 3908 THEN
            sigmoid_f := 1783;
        ELSIF x = 3909 THEN
            sigmoid_f := 1783;
        ELSIF x = 3910 THEN
            sigmoid_f := 1783;
        ELSIF x = 3911 THEN
            sigmoid_f := 1783;
        ELSIF x = 3912 THEN
            sigmoid_f := 1783;
        ELSIF x = 3913 THEN
            sigmoid_f := 1783;
        ELSIF x = 3914 THEN
            sigmoid_f := 1783;
        ELSIF x = 3915 THEN
            sigmoid_f := 1783;
        ELSIF x = 3916 THEN
            sigmoid_f := 1784;
        ELSIF x = 3917 THEN
            sigmoid_f := 1784;
        ELSIF x = 3918 THEN
            sigmoid_f := 1784;
        ELSIF x = 3919 THEN
            sigmoid_f := 1784;
        ELSIF x = 3920 THEN
            sigmoid_f := 1784;
        ELSIF x = 3921 THEN
            sigmoid_f := 1784;
        ELSIF x = 3922 THEN
            sigmoid_f := 1784;
        ELSIF x = 3923 THEN
            sigmoid_f := 1784;
        ELSIF x = 3924 THEN
            sigmoid_f := 1785;
        ELSIF x = 3925 THEN
            sigmoid_f := 1785;
        ELSIF x = 3926 THEN
            sigmoid_f := 1785;
        ELSIF x = 3927 THEN
            sigmoid_f := 1785;
        ELSIF x = 3928 THEN
            sigmoid_f := 1785;
        ELSIF x = 3929 THEN
            sigmoid_f := 1785;
        ELSIF x = 3930 THEN
            sigmoid_f := 1785;
        ELSIF x = 3931 THEN
            sigmoid_f := 1785;
        ELSIF x = 3932 THEN
            sigmoid_f := 1785;
        ELSIF x = 3933 THEN
            sigmoid_f := 1786;
        ELSIF x = 3934 THEN
            sigmoid_f := 1786;
        ELSIF x = 3935 THEN
            sigmoid_f := 1786;
        ELSIF x = 3936 THEN
            sigmoid_f := 1786;
        ELSIF x = 3937 THEN
            sigmoid_f := 1786;
        ELSIF x = 3938 THEN
            sigmoid_f := 1786;
        ELSIF x = 3939 THEN
            sigmoid_f := 1786;
        ELSIF x = 3940 THEN
            sigmoid_f := 1786;
        ELSIF x = 3941 THEN
            sigmoid_f := 1786;
        ELSIF x = 3942 THEN
            sigmoid_f := 1787;
        ELSIF x = 3943 THEN
            sigmoid_f := 1787;
        ELSIF x = 3944 THEN
            sigmoid_f := 1787;
        ELSIF x = 3945 THEN
            sigmoid_f := 1787;
        ELSIF x = 3946 THEN
            sigmoid_f := 1787;
        ELSIF x = 3947 THEN
            sigmoid_f := 1787;
        ELSIF x = 3948 THEN
            sigmoid_f := 1787;
        ELSIF x = 3949 THEN
            sigmoid_f := 1787;
        ELSIF x = 3950 THEN
            sigmoid_f := 1788;
        ELSIF x = 3951 THEN
            sigmoid_f := 1788;
        ELSIF x = 3952 THEN
            sigmoid_f := 1788;
        ELSIF x = 3953 THEN
            sigmoid_f := 1788;
        ELSIF x = 3954 THEN
            sigmoid_f := 1788;
        ELSIF x = 3955 THEN
            sigmoid_f := 1788;
        ELSIF x = 3956 THEN
            sigmoid_f := 1788;
        ELSIF x = 3957 THEN
            sigmoid_f := 1788;
        ELSIF x = 3958 THEN
            sigmoid_f := 1788;
        ELSIF x = 3959 THEN
            sigmoid_f := 1789;
        ELSIF x = 3960 THEN
            sigmoid_f := 1789;
        ELSIF x = 3961 THEN
            sigmoid_f := 1789;
        ELSIF x = 3962 THEN
            sigmoid_f := 1789;
        ELSIF x = 3963 THEN
            sigmoid_f := 1789;
        ELSIF x = 3964 THEN
            sigmoid_f := 1789;
        ELSIF x = 3965 THEN
            sigmoid_f := 1789;
        ELSIF x = 3966 THEN
            sigmoid_f := 1789;
        ELSIF x = 3967 THEN
            sigmoid_f := 1790;
        ELSIF x = 3968 THEN
            sigmoid_f := 1790;
        ELSIF x = 3969 THEN
            sigmoid_f := 1790;
        ELSIF x = 3970 THEN
            sigmoid_f := 1790;
        ELSIF x = 3971 THEN
            sigmoid_f := 1790;
        ELSIF x = 3972 THEN
            sigmoid_f := 1790;
        ELSIF x = 3973 THEN
            sigmoid_f := 1790;
        ELSIF x = 3974 THEN
            sigmoid_f := 1790;
        ELSIF x = 3975 THEN
            sigmoid_f := 1790;
        ELSIF x = 3976 THEN
            sigmoid_f := 1791;
        ELSIF x = 3977 THEN
            sigmoid_f := 1791;
        ELSIF x = 3978 THEN
            sigmoid_f := 1791;
        ELSIF x = 3979 THEN
            sigmoid_f := 1791;
        ELSIF x = 3980 THEN
            sigmoid_f := 1791;
        ELSIF x = 3981 THEN
            sigmoid_f := 1791;
        ELSIF x = 3982 THEN
            sigmoid_f := 1791;
        ELSIF x = 3983 THEN
            sigmoid_f := 1791;
        ELSIF x = 3984 THEN
            sigmoid_f := 1791;
        ELSIF x = 3985 THEN
            sigmoid_f := 1792;
        ELSIF x = 3986 THEN
            sigmoid_f := 1792;
        ELSIF x = 3987 THEN
            sigmoid_f := 1792;
        ELSIF x = 3988 THEN
            sigmoid_f := 1792;
        ELSIF x = 3989 THEN
            sigmoid_f := 1792;
        ELSIF x = 3990 THEN
            sigmoid_f := 1792;
        ELSIF x = 3991 THEN
            sigmoid_f := 1792;
        ELSIF x = 3992 THEN
            sigmoid_f := 1792;
        ELSIF x = 3993 THEN
            sigmoid_f := 1793;
        ELSIF x = 3994 THEN
            sigmoid_f := 1793;
        ELSIF x = 3995 THEN
            sigmoid_f := 1793;
        ELSIF x = 3996 THEN
            sigmoid_f := 1793;
        ELSIF x = 3997 THEN
            sigmoid_f := 1793;
        ELSIF x = 3998 THEN
            sigmoid_f := 1793;
        ELSIF x = 3999 THEN
            sigmoid_f := 1793;
        ELSIF x = 4000 THEN
            sigmoid_f := 1793;
        ELSIF x = 4001 THEN
            sigmoid_f := 1793;
        ELSIF x = 4002 THEN
            sigmoid_f := 1794;
        ELSIF x = 4003 THEN
            sigmoid_f := 1794;
        ELSIF x = 4004 THEN
            sigmoid_f := 1794;
        ELSIF x = 4005 THEN
            sigmoid_f := 1794;
        ELSIF x = 4006 THEN
            sigmoid_f := 1794;
        ELSIF x = 4007 THEN
            sigmoid_f := 1794;
        ELSIF x = 4008 THEN
            sigmoid_f := 1794;
        ELSIF x = 4009 THEN
            sigmoid_f := 1794;
        ELSIF x = 4010 THEN
            sigmoid_f := 1795;
        ELSIF x = 4011 THEN
            sigmoid_f := 1795;
        ELSIF x = 4012 THEN
            sigmoid_f := 1795;
        ELSIF x = 4013 THEN
            sigmoid_f := 1795;
        ELSIF x = 4014 THEN
            sigmoid_f := 1795;
        ELSIF x = 4015 THEN
            sigmoid_f := 1795;
        ELSIF x = 4016 THEN
            sigmoid_f := 1795;
        ELSIF x = 4017 THEN
            sigmoid_f := 1795;
        ELSIF x = 4018 THEN
            sigmoid_f := 1795;
        ELSIF x = 4019 THEN
            sigmoid_f := 1796;
        ELSIF x = 4020 THEN
            sigmoid_f := 1796;
        ELSIF x = 4021 THEN
            sigmoid_f := 1796;
        ELSIF x = 4022 THEN
            sigmoid_f := 1796;
        ELSIF x = 4023 THEN
            sigmoid_f := 1796;
        ELSIF x = 4024 THEN
            sigmoid_f := 1796;
        ELSIF x = 4025 THEN
            sigmoid_f := 1796;
        ELSIF x = 4026 THEN
            sigmoid_f := 1796;
        ELSIF x = 4027 THEN
            sigmoid_f := 1796;
        ELSIF x = 4028 THEN
            sigmoid_f := 1797;
        ELSIF x = 4029 THEN
            sigmoid_f := 1797;
        ELSIF x = 4030 THEN
            sigmoid_f := 1797;
        ELSIF x = 4031 THEN
            sigmoid_f := 1797;
        ELSIF x = 4032 THEN
            sigmoid_f := 1797;
        ELSIF x = 4033 THEN
            sigmoid_f := 1797;
        ELSIF x = 4034 THEN
            sigmoid_f := 1797;
        ELSIF x = 4035 THEN
            sigmoid_f := 1797;
        ELSIF x = 4036 THEN
            sigmoid_f := 1798;
        ELSIF x = 4037 THEN
            sigmoid_f := 1798;
        ELSIF x = 4038 THEN
            sigmoid_f := 1798;
        ELSIF x = 4039 THEN
            sigmoid_f := 1798;
        ELSIF x = 4040 THEN
            sigmoid_f := 1798;
        ELSIF x = 4041 THEN
            sigmoid_f := 1798;
        ELSIF x = 4042 THEN
            sigmoid_f := 1798;
        ELSIF x = 4043 THEN
            sigmoid_f := 1798;
        ELSIF x = 4044 THEN
            sigmoid_f := 1798;
        ELSIF x = 4045 THEN
            sigmoid_f := 1799;
        ELSIF x = 4046 THEN
            sigmoid_f := 1799;
        ELSIF x = 4047 THEN
            sigmoid_f := 1799;
        ELSIF x = 4048 THEN
            sigmoid_f := 1799;
        ELSIF x = 4049 THEN
            sigmoid_f := 1799;
        ELSIF x = 4050 THEN
            sigmoid_f := 1799;
        ELSIF x = 4051 THEN
            sigmoid_f := 1799;
        ELSIF x = 4052 THEN
            sigmoid_f := 1799;
        ELSIF x = 4053 THEN
            sigmoid_f := 1800;
        ELSIF x = 4054 THEN
            sigmoid_f := 1800;
        ELSIF x = 4055 THEN
            sigmoid_f := 1800;
        ELSIF x = 4056 THEN
            sigmoid_f := 1800;
        ELSIF x = 4057 THEN
            sigmoid_f := 1800;
        ELSIF x = 4058 THEN
            sigmoid_f := 1800;
        ELSIF x = 4059 THEN
            sigmoid_f := 1800;
        ELSIF x = 4060 THEN
            sigmoid_f := 1800;
        ELSIF x = 4061 THEN
            sigmoid_f := 1800;
        ELSIF x = 4062 THEN
            sigmoid_f := 1801;
        ELSIF x = 4063 THEN
            sigmoid_f := 1801;
        ELSIF x = 4064 THEN
            sigmoid_f := 1801;
        ELSIF x = 4065 THEN
            sigmoid_f := 1801;
        ELSIF x = 4066 THEN
            sigmoid_f := 1801;
        ELSIF x = 4067 THEN
            sigmoid_f := 1801;
        ELSIF x = 4068 THEN
            sigmoid_f := 1801;
        ELSIF x = 4069 THEN
            sigmoid_f := 1801;
        ELSIF x = 4070 THEN
            sigmoid_f := 1801;
        ELSIF x = 4071 THEN
            sigmoid_f := 1802;
        ELSIF x = 4072 THEN
            sigmoid_f := 1802;
        ELSIF x = 4073 THEN
            sigmoid_f := 1802;
        ELSIF x = 4074 THEN
            sigmoid_f := 1802;
        ELSIF x = 4075 THEN
            sigmoid_f := 1802;
        ELSIF x = 4076 THEN
            sigmoid_f := 1802;
        ELSIF x = 4077 THEN
            sigmoid_f := 1802;
        ELSIF x = 4078 THEN
            sigmoid_f := 1802;
        ELSIF x = 4079 THEN
            sigmoid_f := 1803;
        ELSIF x = 4080 THEN
            sigmoid_f := 1803;
        ELSIF x = 4081 THEN
            sigmoid_f := 1803;
        ELSIF x = 4082 THEN
            sigmoid_f := 1803;
        ELSIF x = 4083 THEN
            sigmoid_f := 1803;
        ELSIF x = 4084 THEN
            sigmoid_f := 1803;
        ELSIF x = 4085 THEN
            sigmoid_f := 1803;
        ELSIF x = 4086 THEN
            sigmoid_f := 1803;
        ELSIF x = 4087 THEN
            sigmoid_f := 1803;
        ELSIF x = 4088 THEN
            sigmoid_f := 1804;
        ELSIF x = 4089 THEN
            sigmoid_f := 1804;
        ELSIF x = 4090 THEN
            sigmoid_f := 1804;
        ELSIF x = 4091 THEN
            sigmoid_f := 1804;
        ELSIF x = 4092 THEN
            sigmoid_f := 1804;
        ELSIF x = 4093 THEN
            sigmoid_f := 1804;
        ELSIF x = 4094 THEN
            sigmoid_f := 1804;
        ELSIF x = 4095 THEN
            sigmoid_f := 1804;
        ELSIF x = 4096 THEN
            sigmoid_f := 1805;
        ELSIF x = 4097 THEN
            sigmoid_f := 1805;
        ELSIF x = 4098 THEN
            sigmoid_f := 1805;
        ELSIF x = 4099 THEN
            sigmoid_f := 1805;
        ELSIF x = 4100 THEN
            sigmoid_f := 1805;
        ELSIF x = 4101 THEN
            sigmoid_f := 1805;
        ELSIF x = 4102 THEN
            sigmoid_f := 1805;
        ELSIF x = 4103 THEN
            sigmoid_f := 1805;
        ELSIF x = 4104 THEN
            sigmoid_f := 1805;
        ELSIF x = 4105 THEN
            sigmoid_f := 1805;
        ELSIF x = 4106 THEN
            sigmoid_f := 1805;
        ELSIF x = 4107 THEN
            sigmoid_f := 1806;
        ELSIF x = 4108 THEN
            sigmoid_f := 1806;
        ELSIF x = 4109 THEN
            sigmoid_f := 1806;
        ELSIF x = 4110 THEN
            sigmoid_f := 1806;
        ELSIF x = 4111 THEN
            sigmoid_f := 1806;
        ELSIF x = 4112 THEN
            sigmoid_f := 1806;
        ELSIF x = 4113 THEN
            sigmoid_f := 1806;
        ELSIF x = 4114 THEN
            sigmoid_f := 1806;
        ELSIF x = 4115 THEN
            sigmoid_f := 1806;
        ELSIF x = 4116 THEN
            sigmoid_f := 1806;
        ELSIF x = 4117 THEN
            sigmoid_f := 1806;
        ELSIF x = 4118 THEN
            sigmoid_f := 1807;
        ELSIF x = 4119 THEN
            sigmoid_f := 1807;
        ELSIF x = 4120 THEN
            sigmoid_f := 1807;
        ELSIF x = 4121 THEN
            sigmoid_f := 1807;
        ELSIF x = 4122 THEN
            sigmoid_f := 1807;
        ELSIF x = 4123 THEN
            sigmoid_f := 1807;
        ELSIF x = 4124 THEN
            sigmoid_f := 1807;
        ELSIF x = 4125 THEN
            sigmoid_f := 1807;
        ELSIF x = 4126 THEN
            sigmoid_f := 1807;
        ELSIF x = 4127 THEN
            sigmoid_f := 1807;
        ELSIF x = 4128 THEN
            sigmoid_f := 1808;
        ELSIF x = 4129 THEN
            sigmoid_f := 1808;
        ELSIF x = 4130 THEN
            sigmoid_f := 1808;
        ELSIF x = 4131 THEN
            sigmoid_f := 1808;
        ELSIF x = 4132 THEN
            sigmoid_f := 1808;
        ELSIF x = 4133 THEN
            sigmoid_f := 1808;
        ELSIF x = 4134 THEN
            sigmoid_f := 1808;
        ELSIF x = 4135 THEN
            sigmoid_f := 1808;
        ELSIF x = 4136 THEN
            sigmoid_f := 1808;
        ELSIF x = 4137 THEN
            sigmoid_f := 1808;
        ELSIF x = 4138 THEN
            sigmoid_f := 1808;
        ELSIF x = 4139 THEN
            sigmoid_f := 1809;
        ELSIF x = 4140 THEN
            sigmoid_f := 1809;
        ELSIF x = 4141 THEN
            sigmoid_f := 1809;
        ELSIF x = 4142 THEN
            sigmoid_f := 1809;
        ELSIF x = 4143 THEN
            sigmoid_f := 1809;
        ELSIF x = 4144 THEN
            sigmoid_f := 1809;
        ELSIF x = 4145 THEN
            sigmoid_f := 1809;
        ELSIF x = 4146 THEN
            sigmoid_f := 1809;
        ELSIF x = 4147 THEN
            sigmoid_f := 1809;
        ELSIF x = 4148 THEN
            sigmoid_f := 1809;
        ELSIF x = 4149 THEN
            sigmoid_f := 1809;
        ELSIF x = 4150 THEN
            sigmoid_f := 1810;
        ELSIF x = 4151 THEN
            sigmoid_f := 1810;
        ELSIF x = 4152 THEN
            sigmoid_f := 1810;
        ELSIF x = 4153 THEN
            sigmoid_f := 1810;
        ELSIF x = 4154 THEN
            sigmoid_f := 1810;
        ELSIF x = 4155 THEN
            sigmoid_f := 1810;
        ELSIF x = 4156 THEN
            sigmoid_f := 1810;
        ELSIF x = 4157 THEN
            sigmoid_f := 1810;
        ELSIF x = 4158 THEN
            sigmoid_f := 1810;
        ELSIF x = 4159 THEN
            sigmoid_f := 1810;
        ELSIF x = 4160 THEN
            sigmoid_f := 1811;
        ELSIF x = 4161 THEN
            sigmoid_f := 1811;
        ELSIF x = 4162 THEN
            sigmoid_f := 1811;
        ELSIF x = 4163 THEN
            sigmoid_f := 1811;
        ELSIF x = 4164 THEN
            sigmoid_f := 1811;
        ELSIF x = 4165 THEN
            sigmoid_f := 1811;
        ELSIF x = 4166 THEN
            sigmoid_f := 1811;
        ELSIF x = 4167 THEN
            sigmoid_f := 1811;
        ELSIF x = 4168 THEN
            sigmoid_f := 1811;
        ELSIF x = 4169 THEN
            sigmoid_f := 1811;
        ELSIF x = 4170 THEN
            sigmoid_f := 1811;
        ELSIF x = 4171 THEN
            sigmoid_f := 1812;
        ELSIF x = 4172 THEN
            sigmoid_f := 1812;
        ELSIF x = 4173 THEN
            sigmoid_f := 1812;
        ELSIF x = 4174 THEN
            sigmoid_f := 1812;
        ELSIF x = 4175 THEN
            sigmoid_f := 1812;
        ELSIF x = 4176 THEN
            sigmoid_f := 1812;
        ELSIF x = 4177 THEN
            sigmoid_f := 1812;
        ELSIF x = 4178 THEN
            sigmoid_f := 1812;
        ELSIF x = 4179 THEN
            sigmoid_f := 1812;
        ELSIF x = 4180 THEN
            sigmoid_f := 1812;
        ELSIF x = 4181 THEN
            sigmoid_f := 1813;
        ELSIF x = 4182 THEN
            sigmoid_f := 1813;
        ELSIF x = 4183 THEN
            sigmoid_f := 1813;
        ELSIF x = 4184 THEN
            sigmoid_f := 1813;
        ELSIF x = 4185 THEN
            sigmoid_f := 1813;
        ELSIF x = 4186 THEN
            sigmoid_f := 1813;
        ELSIF x = 4187 THEN
            sigmoid_f := 1813;
        ELSIF x = 4188 THEN
            sigmoid_f := 1813;
        ELSIF x = 4189 THEN
            sigmoid_f := 1813;
        ELSIF x = 4190 THEN
            sigmoid_f := 1813;
        ELSIF x = 4191 THEN
            sigmoid_f := 1813;
        ELSIF x = 4192 THEN
            sigmoid_f := 1814;
        ELSIF x = 4193 THEN
            sigmoid_f := 1814;
        ELSIF x = 4194 THEN
            sigmoid_f := 1814;
        ELSIF x = 4195 THEN
            sigmoid_f := 1814;
        ELSIF x = 4196 THEN
            sigmoid_f := 1814;
        ELSIF x = 4197 THEN
            sigmoid_f := 1814;
        ELSIF x = 4198 THEN
            sigmoid_f := 1814;
        ELSIF x = 4199 THEN
            sigmoid_f := 1814;
        ELSIF x = 4200 THEN
            sigmoid_f := 1814;
        ELSIF x = 4201 THEN
            sigmoid_f := 1814;
        ELSIF x = 4202 THEN
            sigmoid_f := 1814;
        ELSIF x = 4203 THEN
            sigmoid_f := 1815;
        ELSIF x = 4204 THEN
            sigmoid_f := 1815;
        ELSIF x = 4205 THEN
            sigmoid_f := 1815;
        ELSIF x = 4206 THEN
            sigmoid_f := 1815;
        ELSIF x = 4207 THEN
            sigmoid_f := 1815;
        ELSIF x = 4208 THEN
            sigmoid_f := 1815;
        ELSIF x = 4209 THEN
            sigmoid_f := 1815;
        ELSIF x = 4210 THEN
            sigmoid_f := 1815;
        ELSIF x = 4211 THEN
            sigmoid_f := 1815;
        ELSIF x = 4212 THEN
            sigmoid_f := 1815;
        ELSIF x = 4213 THEN
            sigmoid_f := 1816;
        ELSIF x = 4214 THEN
            sigmoid_f := 1816;
        ELSIF x = 4215 THEN
            sigmoid_f := 1816;
        ELSIF x = 4216 THEN
            sigmoid_f := 1816;
        ELSIF x = 4217 THEN
            sigmoid_f := 1816;
        ELSIF x = 4218 THEN
            sigmoid_f := 1816;
        ELSIF x = 4219 THEN
            sigmoid_f := 1816;
        ELSIF x = 4220 THEN
            sigmoid_f := 1816;
        ELSIF x = 4221 THEN
            sigmoid_f := 1816;
        ELSIF x = 4222 THEN
            sigmoid_f := 1816;
        ELSIF x = 4223 THEN
            sigmoid_f := 1816;
        ELSIF x = 4224 THEN
            sigmoid_f := 1817;
        ELSIF x = 4225 THEN
            sigmoid_f := 1817;
        ELSIF x = 4226 THEN
            sigmoid_f := 1817;
        ELSIF x = 4227 THEN
            sigmoid_f := 1817;
        ELSIF x = 4228 THEN
            sigmoid_f := 1817;
        ELSIF x = 4229 THEN
            sigmoid_f := 1817;
        ELSIF x = 4230 THEN
            sigmoid_f := 1817;
        ELSIF x = 4231 THEN
            sigmoid_f := 1817;
        ELSIF x = 4232 THEN
            sigmoid_f := 1817;
        ELSIF x = 4233 THEN
            sigmoid_f := 1817;
        ELSIF x = 4234 THEN
            sigmoid_f := 1818;
        ELSIF x = 4235 THEN
            sigmoid_f := 1818;
        ELSIF x = 4236 THEN
            sigmoid_f := 1818;
        ELSIF x = 4237 THEN
            sigmoid_f := 1818;
        ELSIF x = 4238 THEN
            sigmoid_f := 1818;
        ELSIF x = 4239 THEN
            sigmoid_f := 1818;
        ELSIF x = 4240 THEN
            sigmoid_f := 1818;
        ELSIF x = 4241 THEN
            sigmoid_f := 1818;
        ELSIF x = 4242 THEN
            sigmoid_f := 1818;
        ELSIF x = 4243 THEN
            sigmoid_f := 1818;
        ELSIF x = 4244 THEN
            sigmoid_f := 1818;
        ELSIF x = 4245 THEN
            sigmoid_f := 1819;
        ELSIF x = 4246 THEN
            sigmoid_f := 1819;
        ELSIF x = 4247 THEN
            sigmoid_f := 1819;
        ELSIF x = 4248 THEN
            sigmoid_f := 1819;
        ELSIF x = 4249 THEN
            sigmoid_f := 1819;
        ELSIF x = 4250 THEN
            sigmoid_f := 1819;
        ELSIF x = 4251 THEN
            sigmoid_f := 1819;
        ELSIF x = 4252 THEN
            sigmoid_f := 1819;
        ELSIF x = 4253 THEN
            sigmoid_f := 1819;
        ELSIF x = 4254 THEN
            sigmoid_f := 1819;
        ELSIF x = 4255 THEN
            sigmoid_f := 1819;
        ELSIF x = 4256 THEN
            sigmoid_f := 1820;
        ELSIF x = 4257 THEN
            sigmoid_f := 1820;
        ELSIF x = 4258 THEN
            sigmoid_f := 1820;
        ELSIF x = 4259 THEN
            sigmoid_f := 1820;
        ELSIF x = 4260 THEN
            sigmoid_f := 1820;
        ELSIF x = 4261 THEN
            sigmoid_f := 1820;
        ELSIF x = 4262 THEN
            sigmoid_f := 1820;
        ELSIF x = 4263 THEN
            sigmoid_f := 1820;
        ELSIF x = 4264 THEN
            sigmoid_f := 1820;
        ELSIF x = 4265 THEN
            sigmoid_f := 1820;
        ELSIF x = 4266 THEN
            sigmoid_f := 1821;
        ELSIF x = 4267 THEN
            sigmoid_f := 1821;
        ELSIF x = 4268 THEN
            sigmoid_f := 1821;
        ELSIF x = 4269 THEN
            sigmoid_f := 1821;
        ELSIF x = 4270 THEN
            sigmoid_f := 1821;
        ELSIF x = 4271 THEN
            sigmoid_f := 1821;
        ELSIF x = 4272 THEN
            sigmoid_f := 1821;
        ELSIF x = 4273 THEN
            sigmoid_f := 1821;
        ELSIF x = 4274 THEN
            sigmoid_f := 1821;
        ELSIF x = 4275 THEN
            sigmoid_f := 1821;
        ELSIF x = 4276 THEN
            sigmoid_f := 1821;
        ELSIF x = 4277 THEN
            sigmoid_f := 1822;
        ELSIF x = 4278 THEN
            sigmoid_f := 1822;
        ELSIF x = 4279 THEN
            sigmoid_f := 1822;
        ELSIF x = 4280 THEN
            sigmoid_f := 1822;
        ELSIF x = 4281 THEN
            sigmoid_f := 1822;
        ELSIF x = 4282 THEN
            sigmoid_f := 1822;
        ELSIF x = 4283 THEN
            sigmoid_f := 1822;
        ELSIF x = 4284 THEN
            sigmoid_f := 1822;
        ELSIF x = 4285 THEN
            sigmoid_f := 1822;
        ELSIF x = 4286 THEN
            sigmoid_f := 1822;
        ELSIF x = 4287 THEN
            sigmoid_f := 1822;
        ELSIF x = 4288 THEN
            sigmoid_f := 1823;
        ELSIF x = 4289 THEN
            sigmoid_f := 1823;
        ELSIF x = 4290 THEN
            sigmoid_f := 1823;
        ELSIF x = 4291 THEN
            sigmoid_f := 1823;
        ELSIF x = 4292 THEN
            sigmoid_f := 1823;
        ELSIF x = 4293 THEN
            sigmoid_f := 1823;
        ELSIF x = 4294 THEN
            sigmoid_f := 1823;
        ELSIF x = 4295 THEN
            sigmoid_f := 1823;
        ELSIF x = 4296 THEN
            sigmoid_f := 1823;
        ELSIF x = 4297 THEN
            sigmoid_f := 1823;
        ELSIF x = 4298 THEN
            sigmoid_f := 1824;
        ELSIF x = 4299 THEN
            sigmoid_f := 1824;
        ELSIF x = 4300 THEN
            sigmoid_f := 1824;
        ELSIF x = 4301 THEN
            sigmoid_f := 1824;
        ELSIF x = 4302 THEN
            sigmoid_f := 1824;
        ELSIF x = 4303 THEN
            sigmoid_f := 1824;
        ELSIF x = 4304 THEN
            sigmoid_f := 1824;
        ELSIF x = 4305 THEN
            sigmoid_f := 1824;
        ELSIF x = 4306 THEN
            sigmoid_f := 1824;
        ELSIF x = 4307 THEN
            sigmoid_f := 1824;
        ELSIF x = 4308 THEN
            sigmoid_f := 1824;
        ELSIF x = 4309 THEN
            sigmoid_f := 1825;
        ELSIF x = 4310 THEN
            sigmoid_f := 1825;
        ELSIF x = 4311 THEN
            sigmoid_f := 1825;
        ELSIF x = 4312 THEN
            sigmoid_f := 1825;
        ELSIF x = 4313 THEN
            sigmoid_f := 1825;
        ELSIF x = 4314 THEN
            sigmoid_f := 1825;
        ELSIF x = 4315 THEN
            sigmoid_f := 1825;
        ELSIF x = 4316 THEN
            sigmoid_f := 1825;
        ELSIF x = 4317 THEN
            sigmoid_f := 1825;
        ELSIF x = 4318 THEN
            sigmoid_f := 1825;
        ELSIF x = 4319 THEN
            sigmoid_f := 1826;
        ELSIF x = 4320 THEN
            sigmoid_f := 1826;
        ELSIF x = 4321 THEN
            sigmoid_f := 1826;
        ELSIF x = 4322 THEN
            sigmoid_f := 1826;
        ELSIF x = 4323 THEN
            sigmoid_f := 1826;
        ELSIF x = 4324 THEN
            sigmoid_f := 1826;
        ELSIF x = 4325 THEN
            sigmoid_f := 1826;
        ELSIF x = 4326 THEN
            sigmoid_f := 1826;
        ELSIF x = 4327 THEN
            sigmoid_f := 1826;
        ELSIF x = 4328 THEN
            sigmoid_f := 1826;
        ELSIF x = 4329 THEN
            sigmoid_f := 1826;
        ELSIF x = 4330 THEN
            sigmoid_f := 1827;
        ELSIF x = 4331 THEN
            sigmoid_f := 1827;
        ELSIF x = 4332 THEN
            sigmoid_f := 1827;
        ELSIF x = 4333 THEN
            sigmoid_f := 1827;
        ELSIF x = 4334 THEN
            sigmoid_f := 1827;
        ELSIF x = 4335 THEN
            sigmoid_f := 1827;
        ELSIF x = 4336 THEN
            sigmoid_f := 1827;
        ELSIF x = 4337 THEN
            sigmoid_f := 1827;
        ELSIF x = 4338 THEN
            sigmoid_f := 1827;
        ELSIF x = 4339 THEN
            sigmoid_f := 1827;
        ELSIF x = 4340 THEN
            sigmoid_f := 1827;
        ELSIF x = 4341 THEN
            sigmoid_f := 1828;
        ELSIF x = 4342 THEN
            sigmoid_f := 1828;
        ELSIF x = 4343 THEN
            sigmoid_f := 1828;
        ELSIF x = 4344 THEN
            sigmoid_f := 1828;
        ELSIF x = 4345 THEN
            sigmoid_f := 1828;
        ELSIF x = 4346 THEN
            sigmoid_f := 1828;
        ELSIF x = 4347 THEN
            sigmoid_f := 1828;
        ELSIF x = 4348 THEN
            sigmoid_f := 1828;
        ELSIF x = 4349 THEN
            sigmoid_f := 1828;
        ELSIF x = 4350 THEN
            sigmoid_f := 1828;
        ELSIF x = 4351 THEN
            sigmoid_f := 1829;
        ELSIF x = 4352 THEN
            sigmoid_f := 1829;
        ELSIF x = 4353 THEN
            sigmoid_f := 1829;
        ELSIF x = 4354 THEN
            sigmoid_f := 1829;
        ELSIF x = 4355 THEN
            sigmoid_f := 1829;
        ELSIF x = 4356 THEN
            sigmoid_f := 1829;
        ELSIF x = 4357 THEN
            sigmoid_f := 1829;
        ELSIF x = 4358 THEN
            sigmoid_f := 1829;
        ELSIF x = 4359 THEN
            sigmoid_f := 1829;
        ELSIF x = 4360 THEN
            sigmoid_f := 1829;
        ELSIF x = 4361 THEN
            sigmoid_f := 1829;
        ELSIF x = 4362 THEN
            sigmoid_f := 1830;
        ELSIF x = 4363 THEN
            sigmoid_f := 1830;
        ELSIF x = 4364 THEN
            sigmoid_f := 1830;
        ELSIF x = 4365 THEN
            sigmoid_f := 1830;
        ELSIF x = 4366 THEN
            sigmoid_f := 1830;
        ELSIF x = 4367 THEN
            sigmoid_f := 1830;
        ELSIF x = 4368 THEN
            sigmoid_f := 1830;
        ELSIF x = 4369 THEN
            sigmoid_f := 1830;
        ELSIF x = 4370 THEN
            sigmoid_f := 1830;
        ELSIF x = 4371 THEN
            sigmoid_f := 1830;
        ELSIF x = 4372 THEN
            sigmoid_f := 1831;
        ELSIF x = 4373 THEN
            sigmoid_f := 1831;
        ELSIF x = 4374 THEN
            sigmoid_f := 1831;
        ELSIF x = 4375 THEN
            sigmoid_f := 1831;
        ELSIF x = 4376 THEN
            sigmoid_f := 1831;
        ELSIF x = 4377 THEN
            sigmoid_f := 1831;
        ELSIF x = 4378 THEN
            sigmoid_f := 1831;
        ELSIF x = 4379 THEN
            sigmoid_f := 1831;
        ELSIF x = 4380 THEN
            sigmoid_f := 1831;
        ELSIF x = 4381 THEN
            sigmoid_f := 1831;
        ELSIF x = 4382 THEN
            sigmoid_f := 1831;
        ELSIF x = 4383 THEN
            sigmoid_f := 1832;
        ELSIF x = 4384 THEN
            sigmoid_f := 1832;
        ELSIF x = 4385 THEN
            sigmoid_f := 1832;
        ELSIF x = 4386 THEN
            sigmoid_f := 1832;
        ELSIF x = 4387 THEN
            sigmoid_f := 1832;
        ELSIF x = 4388 THEN
            sigmoid_f := 1832;
        ELSIF x = 4389 THEN
            sigmoid_f := 1832;
        ELSIF x = 4390 THEN
            sigmoid_f := 1832;
        ELSIF x = 4391 THEN
            sigmoid_f := 1832;
        ELSIF x = 4392 THEN
            sigmoid_f := 1832;
        ELSIF x = 4393 THEN
            sigmoid_f := 1832;
        ELSIF x = 4394 THEN
            sigmoid_f := 1833;
        ELSIF x = 4395 THEN
            sigmoid_f := 1833;
        ELSIF x = 4396 THEN
            sigmoid_f := 1833;
        ELSIF x = 4397 THEN
            sigmoid_f := 1833;
        ELSIF x = 4398 THEN
            sigmoid_f := 1833;
        ELSIF x = 4399 THEN
            sigmoid_f := 1833;
        ELSIF x = 4400 THEN
            sigmoid_f := 1833;
        ELSIF x = 4401 THEN
            sigmoid_f := 1833;
        ELSIF x = 4402 THEN
            sigmoid_f := 1833;
        ELSIF x = 4403 THEN
            sigmoid_f := 1833;
        ELSIF x = 4404 THEN
            sigmoid_f := 1834;
        ELSIF x = 4405 THEN
            sigmoid_f := 1834;
        ELSIF x = 4406 THEN
            sigmoid_f := 1834;
        ELSIF x = 4407 THEN
            sigmoid_f := 1834;
        ELSIF x = 4408 THEN
            sigmoid_f := 1834;
        ELSIF x = 4409 THEN
            sigmoid_f := 1834;
        ELSIF x = 4410 THEN
            sigmoid_f := 1834;
        ELSIF x = 4411 THEN
            sigmoid_f := 1834;
        ELSIF x = 4412 THEN
            sigmoid_f := 1834;
        ELSIF x = 4413 THEN
            sigmoid_f := 1834;
        ELSIF x = 4414 THEN
            sigmoid_f := 1834;
        ELSIF x = 4415 THEN
            sigmoid_f := 1835;
        ELSIF x = 4416 THEN
            sigmoid_f := 1835;
        ELSIF x = 4417 THEN
            sigmoid_f := 1835;
        ELSIF x = 4418 THEN
            sigmoid_f := 1835;
        ELSIF x = 4419 THEN
            sigmoid_f := 1835;
        ELSIF x = 4420 THEN
            sigmoid_f := 1835;
        ELSIF x = 4421 THEN
            sigmoid_f := 1835;
        ELSIF x = 4422 THEN
            sigmoid_f := 1835;
        ELSIF x = 4423 THEN
            sigmoid_f := 1835;
        ELSIF x = 4424 THEN
            sigmoid_f := 1835;
        ELSIF x = 4425 THEN
            sigmoid_f := 1836;
        ELSIF x = 4426 THEN
            sigmoid_f := 1836;
        ELSIF x = 4427 THEN
            sigmoid_f := 1836;
        ELSIF x = 4428 THEN
            sigmoid_f := 1836;
        ELSIF x = 4429 THEN
            sigmoid_f := 1836;
        ELSIF x = 4430 THEN
            sigmoid_f := 1836;
        ELSIF x = 4431 THEN
            sigmoid_f := 1836;
        ELSIF x = 4432 THEN
            sigmoid_f := 1836;
        ELSIF x = 4433 THEN
            sigmoid_f := 1836;
        ELSIF x = 4434 THEN
            sigmoid_f := 1836;
        ELSIF x = 4435 THEN
            sigmoid_f := 1836;
        ELSIF x = 4436 THEN
            sigmoid_f := 1837;
        ELSIF x = 4437 THEN
            sigmoid_f := 1837;
        ELSIF x = 4438 THEN
            sigmoid_f := 1837;
        ELSIF x = 4439 THEN
            sigmoid_f := 1837;
        ELSIF x = 4440 THEN
            sigmoid_f := 1837;
        ELSIF x = 4441 THEN
            sigmoid_f := 1837;
        ELSIF x = 4442 THEN
            sigmoid_f := 1837;
        ELSIF x = 4443 THEN
            sigmoid_f := 1837;
        ELSIF x = 4444 THEN
            sigmoid_f := 1837;
        ELSIF x = 4445 THEN
            sigmoid_f := 1837;
        ELSIF x = 4446 THEN
            sigmoid_f := 1837;
        ELSIF x = 4447 THEN
            sigmoid_f := 1838;
        ELSIF x = 4448 THEN
            sigmoid_f := 1838;
        ELSIF x = 4449 THEN
            sigmoid_f := 1838;
        ELSIF x = 4450 THEN
            sigmoid_f := 1838;
        ELSIF x = 4451 THEN
            sigmoid_f := 1838;
        ELSIF x = 4452 THEN
            sigmoid_f := 1838;
        ELSIF x = 4453 THEN
            sigmoid_f := 1838;
        ELSIF x = 4454 THEN
            sigmoid_f := 1838;
        ELSIF x = 4455 THEN
            sigmoid_f := 1838;
        ELSIF x = 4456 THEN
            sigmoid_f := 1838;
        ELSIF x = 4457 THEN
            sigmoid_f := 1839;
        ELSIF x = 4458 THEN
            sigmoid_f := 1839;
        ELSIF x = 4459 THEN
            sigmoid_f := 1839;
        ELSIF x = 4460 THEN
            sigmoid_f := 1839;
        ELSIF x = 4461 THEN
            sigmoid_f := 1839;
        ELSIF x = 4462 THEN
            sigmoid_f := 1839;
        ELSIF x = 4463 THEN
            sigmoid_f := 1839;
        ELSIF x = 4464 THEN
            sigmoid_f := 1839;
        ELSIF x = 4465 THEN
            sigmoid_f := 1839;
        ELSIF x = 4466 THEN
            sigmoid_f := 1839;
        ELSIF x = 4467 THEN
            sigmoid_f := 1839;
        ELSIF x = 4468 THEN
            sigmoid_f := 1840;
        ELSIF x = 4469 THEN
            sigmoid_f := 1840;
        ELSIF x = 4470 THEN
            sigmoid_f := 1840;
        ELSIF x = 4471 THEN
            sigmoid_f := 1840;
        ELSIF x = 4472 THEN
            sigmoid_f := 1840;
        ELSIF x = 4473 THEN
            sigmoid_f := 1840;
        ELSIF x = 4474 THEN
            sigmoid_f := 1840;
        ELSIF x = 4475 THEN
            sigmoid_f := 1840;
        ELSIF x = 4476 THEN
            sigmoid_f := 1840;
        ELSIF x = 4477 THEN
            sigmoid_f := 1840;
        ELSIF x = 4478 THEN
            sigmoid_f := 1840;
        ELSIF x = 4479 THEN
            sigmoid_f := 1841;
        ELSIF x = 4480 THEN
            sigmoid_f := 1841;
        ELSIF x = 4481 THEN
            sigmoid_f := 1841;
        ELSIF x = 4482 THEN
            sigmoid_f := 1841;
        ELSIF x = 4483 THEN
            sigmoid_f := 1841;
        ELSIF x = 4484 THEN
            sigmoid_f := 1841;
        ELSIF x = 4485 THEN
            sigmoid_f := 1841;
        ELSIF x = 4486 THEN
            sigmoid_f := 1841;
        ELSIF x = 4487 THEN
            sigmoid_f := 1841;
        ELSIF x = 4488 THEN
            sigmoid_f := 1841;
        ELSIF x = 4489 THEN
            sigmoid_f := 1842;
        ELSIF x = 4490 THEN
            sigmoid_f := 1842;
        ELSIF x = 4491 THEN
            sigmoid_f := 1842;
        ELSIF x = 4492 THEN
            sigmoid_f := 1842;
        ELSIF x = 4493 THEN
            sigmoid_f := 1842;
        ELSIF x = 4494 THEN
            sigmoid_f := 1842;
        ELSIF x = 4495 THEN
            sigmoid_f := 1842;
        ELSIF x = 4496 THEN
            sigmoid_f := 1842;
        ELSIF x = 4497 THEN
            sigmoid_f := 1842;
        ELSIF x = 4498 THEN
            sigmoid_f := 1842;
        ELSIF x = 4499 THEN
            sigmoid_f := 1842;
        ELSIF x = 4500 THEN
            sigmoid_f := 1843;
        ELSIF x = 4501 THEN
            sigmoid_f := 1843;
        ELSIF x = 4502 THEN
            sigmoid_f := 1843;
        ELSIF x = 4503 THEN
            sigmoid_f := 1843;
        ELSIF x = 4504 THEN
            sigmoid_f := 1843;
        ELSIF x = 4505 THEN
            sigmoid_f := 1843;
        ELSIF x = 4506 THEN
            sigmoid_f := 1843;
        ELSIF x = 4507 THEN
            sigmoid_f := 1843;
        ELSIF x = 4508 THEN
            sigmoid_f := 1843;
        ELSIF x = 4509 THEN
            sigmoid_f := 1843;
        ELSIF x = 4510 THEN
            sigmoid_f := 1844;
        ELSIF x = 4511 THEN
            sigmoid_f := 1844;
        ELSIF x = 4512 THEN
            sigmoid_f := 1844;
        ELSIF x = 4513 THEN
            sigmoid_f := 1844;
        ELSIF x = 4514 THEN
            sigmoid_f := 1844;
        ELSIF x = 4515 THEN
            sigmoid_f := 1844;
        ELSIF x = 4516 THEN
            sigmoid_f := 1844;
        ELSIF x = 4517 THEN
            sigmoid_f := 1844;
        ELSIF x = 4518 THEN
            sigmoid_f := 1844;
        ELSIF x = 4519 THEN
            sigmoid_f := 1844;
        ELSIF x = 4520 THEN
            sigmoid_f := 1844;
        ELSIF x = 4521 THEN
            sigmoid_f := 1845;
        ELSIF x = 4522 THEN
            sigmoid_f := 1845;
        ELSIF x = 4523 THEN
            sigmoid_f := 1845;
        ELSIF x = 4524 THEN
            sigmoid_f := 1845;
        ELSIF x = 4525 THEN
            sigmoid_f := 1845;
        ELSIF x = 4526 THEN
            sigmoid_f := 1845;
        ELSIF x = 4527 THEN
            sigmoid_f := 1845;
        ELSIF x = 4528 THEN
            sigmoid_f := 1845;
        ELSIF x = 4529 THEN
            sigmoid_f := 1845;
        ELSIF x = 4530 THEN
            sigmoid_f := 1845;
        ELSIF x = 4531 THEN
            sigmoid_f := 1845;
        ELSIF x = 4532 THEN
            sigmoid_f := 1846;
        ELSIF x = 4533 THEN
            sigmoid_f := 1846;
        ELSIF x = 4534 THEN
            sigmoid_f := 1846;
        ELSIF x = 4535 THEN
            sigmoid_f := 1846;
        ELSIF x = 4536 THEN
            sigmoid_f := 1846;
        ELSIF x = 4537 THEN
            sigmoid_f := 1846;
        ELSIF x = 4538 THEN
            sigmoid_f := 1846;
        ELSIF x = 4539 THEN
            sigmoid_f := 1846;
        ELSIF x = 4540 THEN
            sigmoid_f := 1846;
        ELSIF x = 4541 THEN
            sigmoid_f := 1846;
        ELSIF x = 4542 THEN
            sigmoid_f := 1847;
        ELSIF x = 4543 THEN
            sigmoid_f := 1847;
        ELSIF x = 4544 THEN
            sigmoid_f := 1847;
        ELSIF x = 4545 THEN
            sigmoid_f := 1847;
        ELSIF x = 4546 THEN
            sigmoid_f := 1847;
        ELSIF x = 4547 THEN
            sigmoid_f := 1847;
        ELSIF x = 4548 THEN
            sigmoid_f := 1847;
        ELSIF x = 4549 THEN
            sigmoid_f := 1847;
        ELSIF x = 4550 THEN
            sigmoid_f := 1847;
        ELSIF x = 4551 THEN
            sigmoid_f := 1847;
        ELSIF x = 4552 THEN
            sigmoid_f := 1847;
        ELSIF x = 4553 THEN
            sigmoid_f := 1848;
        ELSIF x = 4554 THEN
            sigmoid_f := 1848;
        ELSIF x = 4555 THEN
            sigmoid_f := 1848;
        ELSIF x = 4556 THEN
            sigmoid_f := 1848;
        ELSIF x = 4557 THEN
            sigmoid_f := 1848;
        ELSIF x = 4558 THEN
            sigmoid_f := 1848;
        ELSIF x = 4559 THEN
            sigmoid_f := 1848;
        ELSIF x = 4560 THEN
            sigmoid_f := 1848;
        ELSIF x = 4561 THEN
            sigmoid_f := 1848;
        ELSIF x = 4562 THEN
            sigmoid_f := 1848;
        ELSIF x = 4563 THEN
            sigmoid_f := 1849;
        ELSIF x = 4564 THEN
            sigmoid_f := 1849;
        ELSIF x = 4565 THEN
            sigmoid_f := 1849;
        ELSIF x = 4566 THEN
            sigmoid_f := 1849;
        ELSIF x = 4567 THEN
            sigmoid_f := 1849;
        ELSIF x = 4568 THEN
            sigmoid_f := 1849;
        ELSIF x = 4569 THEN
            sigmoid_f := 1849;
        ELSIF x = 4570 THEN
            sigmoid_f := 1849;
        ELSIF x = 4571 THEN
            sigmoid_f := 1849;
        ELSIF x = 4572 THEN
            sigmoid_f := 1849;
        ELSIF x = 4573 THEN
            sigmoid_f := 1849;
        ELSIF x = 4574 THEN
            sigmoid_f := 1850;
        ELSIF x = 4575 THEN
            sigmoid_f := 1850;
        ELSIF x = 4576 THEN
            sigmoid_f := 1850;
        ELSIF x = 4577 THEN
            sigmoid_f := 1850;
        ELSIF x = 4578 THEN
            sigmoid_f := 1850;
        ELSIF x = 4579 THEN
            sigmoid_f := 1850;
        ELSIF x = 4580 THEN
            sigmoid_f := 1850;
        ELSIF x = 4581 THEN
            sigmoid_f := 1850;
        ELSIF x = 4582 THEN
            sigmoid_f := 1850;
        ELSIF x = 4583 THEN
            sigmoid_f := 1850;
        ELSIF x = 4584 THEN
            sigmoid_f := 1850;
        ELSIF x = 4585 THEN
            sigmoid_f := 1851;
        ELSIF x = 4586 THEN
            sigmoid_f := 1851;
        ELSIF x = 4587 THEN
            sigmoid_f := 1851;
        ELSIF x = 4588 THEN
            sigmoid_f := 1851;
        ELSIF x = 4589 THEN
            sigmoid_f := 1851;
        ELSIF x = 4590 THEN
            sigmoid_f := 1851;
        ELSIF x = 4591 THEN
            sigmoid_f := 1851;
        ELSIF x = 4592 THEN
            sigmoid_f := 1851;
        ELSIF x = 4593 THEN
            sigmoid_f := 1851;
        ELSIF x = 4594 THEN
            sigmoid_f := 1851;
        ELSIF x = 4595 THEN
            sigmoid_f := 1852;
        ELSIF x = 4596 THEN
            sigmoid_f := 1852;
        ELSIF x = 4597 THEN
            sigmoid_f := 1852;
        ELSIF x = 4598 THEN
            sigmoid_f := 1852;
        ELSIF x = 4599 THEN
            sigmoid_f := 1852;
        ELSIF x = 4600 THEN
            sigmoid_f := 1852;
        ELSIF x = 4601 THEN
            sigmoid_f := 1852;
        ELSIF x = 4602 THEN
            sigmoid_f := 1852;
        ELSIF x = 4603 THEN
            sigmoid_f := 1852;
        ELSIF x = 4604 THEN
            sigmoid_f := 1852;
        ELSIF x = 4605 THEN
            sigmoid_f := 1852;
        ELSIF x = 4606 THEN
            sigmoid_f := 1853;
        ELSIF x = 4607 THEN
            sigmoid_f := 1853;
        ELSIF x = 4608 THEN
            sigmoid_f := 1853;
        ELSIF x = 4609 THEN
            sigmoid_f := 1853;
        ELSIF x = 4610 THEN
            sigmoid_f := 1853;
        ELSIF x = 4611 THEN
            sigmoid_f := 1853;
        ELSIF x = 4612 THEN
            sigmoid_f := 1853;
        ELSIF x = 4613 THEN
            sigmoid_f := 1853;
        ELSIF x = 4614 THEN
            sigmoid_f := 1853;
        ELSIF x = 4615 THEN
            sigmoid_f := 1853;
        ELSIF x = 4616 THEN
            sigmoid_f := 1853;
        ELSIF x = 4617 THEN
            sigmoid_f := 1853;
        ELSIF x = 4618 THEN
            sigmoid_f := 1854;
        ELSIF x = 4619 THEN
            sigmoid_f := 1854;
        ELSIF x = 4620 THEN
            sigmoid_f := 1854;
        ELSIF x = 4621 THEN
            sigmoid_f := 1854;
        ELSIF x = 4622 THEN
            sigmoid_f := 1854;
        ELSIF x = 4623 THEN
            sigmoid_f := 1854;
        ELSIF x = 4624 THEN
            sigmoid_f := 1854;
        ELSIF x = 4625 THEN
            sigmoid_f := 1854;
        ELSIF x = 4626 THEN
            sigmoid_f := 1854;
        ELSIF x = 4627 THEN
            sigmoid_f := 1854;
        ELSIF x = 4628 THEN
            sigmoid_f := 1854;
        ELSIF x = 4629 THEN
            sigmoid_f := 1854;
        ELSIF x = 4630 THEN
            sigmoid_f := 1854;
        ELSIF x = 4631 THEN
            sigmoid_f := 1855;
        ELSIF x = 4632 THEN
            sigmoid_f := 1855;
        ELSIF x = 4633 THEN
            sigmoid_f := 1855;
        ELSIF x = 4634 THEN
            sigmoid_f := 1855;
        ELSIF x = 4635 THEN
            sigmoid_f := 1855;
        ELSIF x = 4636 THEN
            sigmoid_f := 1855;
        ELSIF x = 4637 THEN
            sigmoid_f := 1855;
        ELSIF x = 4638 THEN
            sigmoid_f := 1855;
        ELSIF x = 4639 THEN
            sigmoid_f := 1855;
        ELSIF x = 4640 THEN
            sigmoid_f := 1855;
        ELSIF x = 4641 THEN
            sigmoid_f := 1855;
        ELSIF x = 4642 THEN
            sigmoid_f := 1855;
        ELSIF x = 4643 THEN
            sigmoid_f := 1856;
        ELSIF x = 4644 THEN
            sigmoid_f := 1856;
        ELSIF x = 4645 THEN
            sigmoid_f := 1856;
        ELSIF x = 4646 THEN
            sigmoid_f := 1856;
        ELSIF x = 4647 THEN
            sigmoid_f := 1856;
        ELSIF x = 4648 THEN
            sigmoid_f := 1856;
        ELSIF x = 4649 THEN
            sigmoid_f := 1856;
        ELSIF x = 4650 THEN
            sigmoid_f := 1856;
        ELSIF x = 4651 THEN
            sigmoid_f := 1856;
        ELSIF x = 4652 THEN
            sigmoid_f := 1856;
        ELSIF x = 4653 THEN
            sigmoid_f := 1856;
        ELSIF x = 4654 THEN
            sigmoid_f := 1856;
        ELSIF x = 4655 THEN
            sigmoid_f := 1856;
        ELSIF x = 4656 THEN
            sigmoid_f := 1857;
        ELSIF x = 4657 THEN
            sigmoid_f := 1857;
        ELSIF x = 4658 THEN
            sigmoid_f := 1857;
        ELSIF x = 4659 THEN
            sigmoid_f := 1857;
        ELSIF x = 4660 THEN
            sigmoid_f := 1857;
        ELSIF x = 4661 THEN
            sigmoid_f := 1857;
        ELSIF x = 4662 THEN
            sigmoid_f := 1857;
        ELSIF x = 4663 THEN
            sigmoid_f := 1857;
        ELSIF x = 4664 THEN
            sigmoid_f := 1857;
        ELSIF x = 4665 THEN
            sigmoid_f := 1857;
        ELSIF x = 4666 THEN
            sigmoid_f := 1857;
        ELSIF x = 4667 THEN
            sigmoid_f := 1857;
        ELSIF x = 4668 THEN
            sigmoid_f := 1857;
        ELSIF x = 4669 THEN
            sigmoid_f := 1858;
        ELSIF x = 4670 THEN
            sigmoid_f := 1858;
        ELSIF x = 4671 THEN
            sigmoid_f := 1858;
        ELSIF x = 4672 THEN
            sigmoid_f := 1858;
        ELSIF x = 4673 THEN
            sigmoid_f := 1858;
        ELSIF x = 4674 THEN
            sigmoid_f := 1858;
        ELSIF x = 4675 THEN
            sigmoid_f := 1858;
        ELSIF x = 4676 THEN
            sigmoid_f := 1858;
        ELSIF x = 4677 THEN
            sigmoid_f := 1858;
        ELSIF x = 4678 THEN
            sigmoid_f := 1858;
        ELSIF x = 4679 THEN
            sigmoid_f := 1858;
        ELSIF x = 4680 THEN
            sigmoid_f := 1858;
        ELSIF x = 4681 THEN
            sigmoid_f := 1858;
        ELSIF x = 4682 THEN
            sigmoid_f := 1859;
        ELSIF x = 4683 THEN
            sigmoid_f := 1859;
        ELSIF x = 4684 THEN
            sigmoid_f := 1859;
        ELSIF x = 4685 THEN
            sigmoid_f := 1859;
        ELSIF x = 4686 THEN
            sigmoid_f := 1859;
        ELSIF x = 4687 THEN
            sigmoid_f := 1859;
        ELSIF x = 4688 THEN
            sigmoid_f := 1859;
        ELSIF x = 4689 THEN
            sigmoid_f := 1859;
        ELSIF x = 4690 THEN
            sigmoid_f := 1859;
        ELSIF x = 4691 THEN
            sigmoid_f := 1859;
        ELSIF x = 4692 THEN
            sigmoid_f := 1859;
        ELSIF x = 4693 THEN
            sigmoid_f := 1859;
        ELSIF x = 4694 THEN
            sigmoid_f := 1860;
        ELSIF x = 4695 THEN
            sigmoid_f := 1860;
        ELSIF x = 4696 THEN
            sigmoid_f := 1860;
        ELSIF x = 4697 THEN
            sigmoid_f := 1860;
        ELSIF x = 4698 THEN
            sigmoid_f := 1860;
        ELSIF x = 4699 THEN
            sigmoid_f := 1860;
        ELSIF x = 4700 THEN
            sigmoid_f := 1860;
        ELSIF x = 4701 THEN
            sigmoid_f := 1860;
        ELSIF x = 4702 THEN
            sigmoid_f := 1860;
        ELSIF x = 4703 THEN
            sigmoid_f := 1860;
        ELSIF x = 4704 THEN
            sigmoid_f := 1860;
        ELSIF x = 4705 THEN
            sigmoid_f := 1860;
        ELSIF x = 4706 THEN
            sigmoid_f := 1860;
        ELSIF x = 4707 THEN
            sigmoid_f := 1861;
        ELSIF x = 4708 THEN
            sigmoid_f := 1861;
        ELSIF x = 4709 THEN
            sigmoid_f := 1861;
        ELSIF x = 4710 THEN
            sigmoid_f := 1861;
        ELSIF x = 4711 THEN
            sigmoid_f := 1861;
        ELSIF x = 4712 THEN
            sigmoid_f := 1861;
        ELSIF x = 4713 THEN
            sigmoid_f := 1861;
        ELSIF x = 4714 THEN
            sigmoid_f := 1861;
        ELSIF x = 4715 THEN
            sigmoid_f := 1861;
        ELSIF x = 4716 THEN
            sigmoid_f := 1861;
        ELSIF x = 4717 THEN
            sigmoid_f := 1861;
        ELSIF x = 4718 THEN
            sigmoid_f := 1861;
        ELSIF x = 4719 THEN
            sigmoid_f := 1861;
        ELSIF x = 4720 THEN
            sigmoid_f := 1862;
        ELSIF x = 4721 THEN
            sigmoid_f := 1862;
        ELSIF x = 4722 THEN
            sigmoid_f := 1862;
        ELSIF x = 4723 THEN
            sigmoid_f := 1862;
        ELSIF x = 4724 THEN
            sigmoid_f := 1862;
        ELSIF x = 4725 THEN
            sigmoid_f := 1862;
        ELSIF x = 4726 THEN
            sigmoid_f := 1862;
        ELSIF x = 4727 THEN
            sigmoid_f := 1862;
        ELSIF x = 4728 THEN
            sigmoid_f := 1862;
        ELSIF x = 4729 THEN
            sigmoid_f := 1862;
        ELSIF x = 4730 THEN
            sigmoid_f := 1862;
        ELSIF x = 4731 THEN
            sigmoid_f := 1862;
        ELSIF x = 4732 THEN
            sigmoid_f := 1862;
        ELSIF x = 4733 THEN
            sigmoid_f := 1863;
        ELSIF x = 4734 THEN
            sigmoid_f := 1863;
        ELSIF x = 4735 THEN
            sigmoid_f := 1863;
        ELSIF x = 4736 THEN
            sigmoid_f := 1863;
        ELSIF x = 4737 THEN
            sigmoid_f := 1863;
        ELSIF x = 4738 THEN
            sigmoid_f := 1863;
        ELSIF x = 4739 THEN
            sigmoid_f := 1863;
        ELSIF x = 4740 THEN
            sigmoid_f := 1863;
        ELSIF x = 4741 THEN
            sigmoid_f := 1863;
        ELSIF x = 4742 THEN
            sigmoid_f := 1863;
        ELSIF x = 4743 THEN
            sigmoid_f := 1863;
        ELSIF x = 4744 THEN
            sigmoid_f := 1863;
        ELSIF x = 4745 THEN
            sigmoid_f := 1864;
        ELSIF x = 4746 THEN
            sigmoid_f := 1864;
        ELSIF x = 4747 THEN
            sigmoid_f := 1864;
        ELSIF x = 4748 THEN
            sigmoid_f := 1864;
        ELSIF x = 4749 THEN
            sigmoid_f := 1864;
        ELSIF x = 4750 THEN
            sigmoid_f := 1864;
        ELSIF x = 4751 THEN
            sigmoid_f := 1864;
        ELSIF x = 4752 THEN
            sigmoid_f := 1864;
        ELSIF x = 4753 THEN
            sigmoid_f := 1864;
        ELSIF x = 4754 THEN
            sigmoid_f := 1864;
        ELSIF x = 4755 THEN
            sigmoid_f := 1864;
        ELSIF x = 4756 THEN
            sigmoid_f := 1864;
        ELSIF x = 4757 THEN
            sigmoid_f := 1864;
        ELSIF x = 4758 THEN
            sigmoid_f := 1865;
        ELSIF x = 4759 THEN
            sigmoid_f := 1865;
        ELSIF x = 4760 THEN
            sigmoid_f := 1865;
        ELSIF x = 4761 THEN
            sigmoid_f := 1865;
        ELSIF x = 4762 THEN
            sigmoid_f := 1865;
        ELSIF x = 4763 THEN
            sigmoid_f := 1865;
        ELSIF x = 4764 THEN
            sigmoid_f := 1865;
        ELSIF x = 4765 THEN
            sigmoid_f := 1865;
        ELSIF x = 4766 THEN
            sigmoid_f := 1865;
        ELSIF x = 4767 THEN
            sigmoid_f := 1865;
        ELSIF x = 4768 THEN
            sigmoid_f := 1865;
        ELSIF x = 4769 THEN
            sigmoid_f := 1865;
        ELSIF x = 4770 THEN
            sigmoid_f := 1865;
        ELSIF x = 4771 THEN
            sigmoid_f := 1866;
        ELSIF x = 4772 THEN
            sigmoid_f := 1866;
        ELSIF x = 4773 THEN
            sigmoid_f := 1866;
        ELSIF x = 4774 THEN
            sigmoid_f := 1866;
        ELSIF x = 4775 THEN
            sigmoid_f := 1866;
        ELSIF x = 4776 THEN
            sigmoid_f := 1866;
        ELSIF x = 4777 THEN
            sigmoid_f := 1866;
        ELSIF x = 4778 THEN
            sigmoid_f := 1866;
        ELSIF x = 4779 THEN
            sigmoid_f := 1866;
        ELSIF x = 4780 THEN
            sigmoid_f := 1866;
        ELSIF x = 4781 THEN
            sigmoid_f := 1866;
        ELSIF x = 4782 THEN
            sigmoid_f := 1866;
        ELSIF x = 4783 THEN
            sigmoid_f := 1867;
        ELSIF x = 4784 THEN
            sigmoid_f := 1867;
        ELSIF x = 4785 THEN
            sigmoid_f := 1867;
        ELSIF x = 4786 THEN
            sigmoid_f := 1867;
        ELSIF x = 4787 THEN
            sigmoid_f := 1867;
        ELSIF x = 4788 THEN
            sigmoid_f := 1867;
        ELSIF x = 4789 THEN
            sigmoid_f := 1867;
        ELSIF x = 4790 THEN
            sigmoid_f := 1867;
        ELSIF x = 4791 THEN
            sigmoid_f := 1867;
        ELSIF x = 4792 THEN
            sigmoid_f := 1867;
        ELSIF x = 4793 THEN
            sigmoid_f := 1867;
        ELSIF x = 4794 THEN
            sigmoid_f := 1867;
        ELSIF x = 4795 THEN
            sigmoid_f := 1867;
        ELSIF x = 4796 THEN
            sigmoid_f := 1868;
        ELSIF x = 4797 THEN
            sigmoid_f := 1868;
        ELSIF x = 4798 THEN
            sigmoid_f := 1868;
        ELSIF x = 4799 THEN
            sigmoid_f := 1868;
        ELSIF x = 4800 THEN
            sigmoid_f := 1868;
        ELSIF x = 4801 THEN
            sigmoid_f := 1868;
        ELSIF x = 4802 THEN
            sigmoid_f := 1868;
        ELSIF x = 4803 THEN
            sigmoid_f := 1868;
        ELSIF x = 4804 THEN
            sigmoid_f := 1868;
        ELSIF x = 4805 THEN
            sigmoid_f := 1868;
        ELSIF x = 4806 THEN
            sigmoid_f := 1868;
        ELSIF x = 4807 THEN
            sigmoid_f := 1868;
        ELSIF x = 4808 THEN
            sigmoid_f := 1868;
        ELSIF x = 4809 THEN
            sigmoid_f := 1869;
        ELSIF x = 4810 THEN
            sigmoid_f := 1869;
        ELSIF x = 4811 THEN
            sigmoid_f := 1869;
        ELSIF x = 4812 THEN
            sigmoid_f := 1869;
        ELSIF x = 4813 THEN
            sigmoid_f := 1869;
        ELSIF x = 4814 THEN
            sigmoid_f := 1869;
        ELSIF x = 4815 THEN
            sigmoid_f := 1869;
        ELSIF x = 4816 THEN
            sigmoid_f := 1869;
        ELSIF x = 4817 THEN
            sigmoid_f := 1869;
        ELSIF x = 4818 THEN
            sigmoid_f := 1869;
        ELSIF x = 4819 THEN
            sigmoid_f := 1869;
        ELSIF x = 4820 THEN
            sigmoid_f := 1869;
        ELSIF x = 4821 THEN
            sigmoid_f := 1869;
        ELSIF x = 4822 THEN
            sigmoid_f := 1870;
        ELSIF x = 4823 THEN
            sigmoid_f := 1870;
        ELSIF x = 4824 THEN
            sigmoid_f := 1870;
        ELSIF x = 4825 THEN
            sigmoid_f := 1870;
        ELSIF x = 4826 THEN
            sigmoid_f := 1870;
        ELSIF x = 4827 THEN
            sigmoid_f := 1870;
        ELSIF x = 4828 THEN
            sigmoid_f := 1870;
        ELSIF x = 4829 THEN
            sigmoid_f := 1870;
        ELSIF x = 4830 THEN
            sigmoid_f := 1870;
        ELSIF x = 4831 THEN
            sigmoid_f := 1870;
        ELSIF x = 4832 THEN
            sigmoid_f := 1870;
        ELSIF x = 4833 THEN
            sigmoid_f := 1870;
        ELSIF x = 4834 THEN
            sigmoid_f := 1871;
        ELSIF x = 4835 THEN
            sigmoid_f := 1871;
        ELSIF x = 4836 THEN
            sigmoid_f := 1871;
        ELSIF x = 4837 THEN
            sigmoid_f := 1871;
        ELSIF x = 4838 THEN
            sigmoid_f := 1871;
        ELSIF x = 4839 THEN
            sigmoid_f := 1871;
        ELSIF x = 4840 THEN
            sigmoid_f := 1871;
        ELSIF x = 4841 THEN
            sigmoid_f := 1871;
        ELSIF x = 4842 THEN
            sigmoid_f := 1871;
        ELSIF x = 4843 THEN
            sigmoid_f := 1871;
        ELSIF x = 4844 THEN
            sigmoid_f := 1871;
        ELSIF x = 4845 THEN
            sigmoid_f := 1871;
        ELSIF x = 4846 THEN
            sigmoid_f := 1871;
        ELSIF x = 4847 THEN
            sigmoid_f := 1872;
        ELSIF x = 4848 THEN
            sigmoid_f := 1872;
        ELSIF x = 4849 THEN
            sigmoid_f := 1872;
        ELSIF x = 4850 THEN
            sigmoid_f := 1872;
        ELSIF x = 4851 THEN
            sigmoid_f := 1872;
        ELSIF x = 4852 THEN
            sigmoid_f := 1872;
        ELSIF x = 4853 THEN
            sigmoid_f := 1872;
        ELSIF x = 4854 THEN
            sigmoid_f := 1872;
        ELSIF x = 4855 THEN
            sigmoid_f := 1872;
        ELSIF x = 4856 THEN
            sigmoid_f := 1872;
        ELSIF x = 4857 THEN
            sigmoid_f := 1872;
        ELSIF x = 4858 THEN
            sigmoid_f := 1872;
        ELSIF x = 4859 THEN
            sigmoid_f := 1872;
        ELSIF x = 4860 THEN
            sigmoid_f := 1873;
        ELSIF x = 4861 THEN
            sigmoid_f := 1873;
        ELSIF x = 4862 THEN
            sigmoid_f := 1873;
        ELSIF x = 4863 THEN
            sigmoid_f := 1873;
        ELSIF x = 4864 THEN
            sigmoid_f := 1873;
        ELSIF x = 4865 THEN
            sigmoid_f := 1873;
        ELSIF x = 4866 THEN
            sigmoid_f := 1873;
        ELSIF x = 4867 THEN
            sigmoid_f := 1873;
        ELSIF x = 4868 THEN
            sigmoid_f := 1873;
        ELSIF x = 4869 THEN
            sigmoid_f := 1873;
        ELSIF x = 4870 THEN
            sigmoid_f := 1873;
        ELSIF x = 4871 THEN
            sigmoid_f := 1873;
        ELSIF x = 4872 THEN
            sigmoid_f := 1874;
        ELSIF x = 4873 THEN
            sigmoid_f := 1874;
        ELSIF x = 4874 THEN
            sigmoid_f := 1874;
        ELSIF x = 4875 THEN
            sigmoid_f := 1874;
        ELSIF x = 4876 THEN
            sigmoid_f := 1874;
        ELSIF x = 4877 THEN
            sigmoid_f := 1874;
        ELSIF x = 4878 THEN
            sigmoid_f := 1874;
        ELSIF x = 4879 THEN
            sigmoid_f := 1874;
        ELSIF x = 4880 THEN
            sigmoid_f := 1874;
        ELSIF x = 4881 THEN
            sigmoid_f := 1874;
        ELSIF x = 4882 THEN
            sigmoid_f := 1874;
        ELSIF x = 4883 THEN
            sigmoid_f := 1874;
        ELSIF x = 4884 THEN
            sigmoid_f := 1874;
        ELSIF x = 4885 THEN
            sigmoid_f := 1875;
        ELSIF x = 4886 THEN
            sigmoid_f := 1875;
        ELSIF x = 4887 THEN
            sigmoid_f := 1875;
        ELSIF x = 4888 THEN
            sigmoid_f := 1875;
        ELSIF x = 4889 THEN
            sigmoid_f := 1875;
        ELSIF x = 4890 THEN
            sigmoid_f := 1875;
        ELSIF x = 4891 THEN
            sigmoid_f := 1875;
        ELSIF x = 4892 THEN
            sigmoid_f := 1875;
        ELSIF x = 4893 THEN
            sigmoid_f := 1875;
        ELSIF x = 4894 THEN
            sigmoid_f := 1875;
        ELSIF x = 4895 THEN
            sigmoid_f := 1875;
        ELSIF x = 4896 THEN
            sigmoid_f := 1875;
        ELSIF x = 4897 THEN
            sigmoid_f := 1875;
        ELSIF x = 4898 THEN
            sigmoid_f := 1876;
        ELSIF x = 4899 THEN
            sigmoid_f := 1876;
        ELSIF x = 4900 THEN
            sigmoid_f := 1876;
        ELSIF x = 4901 THEN
            sigmoid_f := 1876;
        ELSIF x = 4902 THEN
            sigmoid_f := 1876;
        ELSIF x = 4903 THEN
            sigmoid_f := 1876;
        ELSIF x = 4904 THEN
            sigmoid_f := 1876;
        ELSIF x = 4905 THEN
            sigmoid_f := 1876;
        ELSIF x = 4906 THEN
            sigmoid_f := 1876;
        ELSIF x = 4907 THEN
            sigmoid_f := 1876;
        ELSIF x = 4908 THEN
            sigmoid_f := 1876;
        ELSIF x = 4909 THEN
            sigmoid_f := 1876;
        ELSIF x = 4910 THEN
            sigmoid_f := 1876;
        ELSIF x = 4911 THEN
            sigmoid_f := 1877;
        ELSIF x = 4912 THEN
            sigmoid_f := 1877;
        ELSIF x = 4913 THEN
            sigmoid_f := 1877;
        ELSIF x = 4914 THEN
            sigmoid_f := 1877;
        ELSIF x = 4915 THEN
            sigmoid_f := 1877;
        ELSIF x = 4916 THEN
            sigmoid_f := 1877;
        ELSIF x = 4917 THEN
            sigmoid_f := 1877;
        ELSIF x = 4918 THEN
            sigmoid_f := 1877;
        ELSIF x = 4919 THEN
            sigmoid_f := 1877;
        ELSIF x = 4920 THEN
            sigmoid_f := 1877;
        ELSIF x = 4921 THEN
            sigmoid_f := 1877;
        ELSIF x = 4922 THEN
            sigmoid_f := 1877;
        ELSIF x = 4923 THEN
            sigmoid_f := 1878;
        ELSIF x = 4924 THEN
            sigmoid_f := 1878;
        ELSIF x = 4925 THEN
            sigmoid_f := 1878;
        ELSIF x = 4926 THEN
            sigmoid_f := 1878;
        ELSIF x = 4927 THEN
            sigmoid_f := 1878;
        ELSIF x = 4928 THEN
            sigmoid_f := 1878;
        ELSIF x = 4929 THEN
            sigmoid_f := 1878;
        ELSIF x = 4930 THEN
            sigmoid_f := 1878;
        ELSIF x = 4931 THEN
            sigmoid_f := 1878;
        ELSIF x = 4932 THEN
            sigmoid_f := 1878;
        ELSIF x = 4933 THEN
            sigmoid_f := 1878;
        ELSIF x = 4934 THEN
            sigmoid_f := 1878;
        ELSIF x = 4935 THEN
            sigmoid_f := 1878;
        ELSIF x = 4936 THEN
            sigmoid_f := 1879;
        ELSIF x = 4937 THEN
            sigmoid_f := 1879;
        ELSIF x = 4938 THEN
            sigmoid_f := 1879;
        ELSIF x = 4939 THEN
            sigmoid_f := 1879;
        ELSIF x = 4940 THEN
            sigmoid_f := 1879;
        ELSIF x = 4941 THEN
            sigmoid_f := 1879;
        ELSIF x = 4942 THEN
            sigmoid_f := 1879;
        ELSIF x = 4943 THEN
            sigmoid_f := 1879;
        ELSIF x = 4944 THEN
            sigmoid_f := 1879;
        ELSIF x = 4945 THEN
            sigmoid_f := 1879;
        ELSIF x = 4946 THEN
            sigmoid_f := 1879;
        ELSIF x = 4947 THEN
            sigmoid_f := 1879;
        ELSIF x = 4948 THEN
            sigmoid_f := 1879;
        ELSIF x = 4949 THEN
            sigmoid_f := 1880;
        ELSIF x = 4950 THEN
            sigmoid_f := 1880;
        ELSIF x = 4951 THEN
            sigmoid_f := 1880;
        ELSIF x = 4952 THEN
            sigmoid_f := 1880;
        ELSIF x = 4953 THEN
            sigmoid_f := 1880;
        ELSIF x = 4954 THEN
            sigmoid_f := 1880;
        ELSIF x = 4955 THEN
            sigmoid_f := 1880;
        ELSIF x = 4956 THEN
            sigmoid_f := 1880;
        ELSIF x = 4957 THEN
            sigmoid_f := 1880;
        ELSIF x = 4958 THEN
            sigmoid_f := 1880;
        ELSIF x = 4959 THEN
            sigmoid_f := 1880;
        ELSIF x = 4960 THEN
            sigmoid_f := 1880;
        ELSIF x = 4961 THEN
            sigmoid_f := 1881;
        ELSIF x = 4962 THEN
            sigmoid_f := 1881;
        ELSIF x = 4963 THEN
            sigmoid_f := 1881;
        ELSIF x = 4964 THEN
            sigmoid_f := 1881;
        ELSIF x = 4965 THEN
            sigmoid_f := 1881;
        ELSIF x = 4966 THEN
            sigmoid_f := 1881;
        ELSIF x = 4967 THEN
            sigmoid_f := 1881;
        ELSIF x = 4968 THEN
            sigmoid_f := 1881;
        ELSIF x = 4969 THEN
            sigmoid_f := 1881;
        ELSIF x = 4970 THEN
            sigmoid_f := 1881;
        ELSIF x = 4971 THEN
            sigmoid_f := 1881;
        ELSIF x = 4972 THEN
            sigmoid_f := 1881;
        ELSIF x = 4973 THEN
            sigmoid_f := 1881;
        ELSIF x = 4974 THEN
            sigmoid_f := 1882;
        ELSIF x = 4975 THEN
            sigmoid_f := 1882;
        ELSIF x = 4976 THEN
            sigmoid_f := 1882;
        ELSIF x = 4977 THEN
            sigmoid_f := 1882;
        ELSIF x = 4978 THEN
            sigmoid_f := 1882;
        ELSIF x = 4979 THEN
            sigmoid_f := 1882;
        ELSIF x = 4980 THEN
            sigmoid_f := 1882;
        ELSIF x = 4981 THEN
            sigmoid_f := 1882;
        ELSIF x = 4982 THEN
            sigmoid_f := 1882;
        ELSIF x = 4983 THEN
            sigmoid_f := 1882;
        ELSIF x = 4984 THEN
            sigmoid_f := 1882;
        ELSIF x = 4985 THEN
            sigmoid_f := 1882;
        ELSIF x = 4986 THEN
            sigmoid_f := 1882;
        ELSIF x = 4987 THEN
            sigmoid_f := 1883;
        ELSIF x = 4988 THEN
            sigmoid_f := 1883;
        ELSIF x = 4989 THEN
            sigmoid_f := 1883;
        ELSIF x = 4990 THEN
            sigmoid_f := 1883;
        ELSIF x = 4991 THEN
            sigmoid_f := 1883;
        ELSIF x = 4992 THEN
            sigmoid_f := 1883;
        ELSIF x = 4993 THEN
            sigmoid_f := 1883;
        ELSIF x = 4994 THEN
            sigmoid_f := 1883;
        ELSIF x = 4995 THEN
            sigmoid_f := 1883;
        ELSIF x = 4996 THEN
            sigmoid_f := 1883;
        ELSIF x = 4997 THEN
            sigmoid_f := 1883;
        ELSIF x = 4998 THEN
            sigmoid_f := 1883;
        ELSIF x = 4999 THEN
            sigmoid_f := 1883;
        ELSIF x = 5000 THEN
            sigmoid_f := 1884;
        ELSIF x = 5001 THEN
            sigmoid_f := 1884;
        ELSIF x = 5002 THEN
            sigmoid_f := 1884;
        ELSIF x = 5003 THEN
            sigmoid_f := 1884;
        ELSIF x = 5004 THEN
            sigmoid_f := 1884;
        ELSIF x = 5005 THEN
            sigmoid_f := 1884;
        ELSIF x = 5006 THEN
            sigmoid_f := 1884;
        ELSIF x = 5007 THEN
            sigmoid_f := 1884;
        ELSIF x = 5008 THEN
            sigmoid_f := 1884;
        ELSIF x = 5009 THEN
            sigmoid_f := 1884;
        ELSIF x = 5010 THEN
            sigmoid_f := 1884;
        ELSIF x = 5011 THEN
            sigmoid_f := 1884;
        ELSIF x = 5012 THEN
            sigmoid_f := 1885;
        ELSIF x = 5013 THEN
            sigmoid_f := 1885;
        ELSIF x = 5014 THEN
            sigmoid_f := 1885;
        ELSIF x = 5015 THEN
            sigmoid_f := 1885;
        ELSIF x = 5016 THEN
            sigmoid_f := 1885;
        ELSIF x = 5017 THEN
            sigmoid_f := 1885;
        ELSIF x = 5018 THEN
            sigmoid_f := 1885;
        ELSIF x = 5019 THEN
            sigmoid_f := 1885;
        ELSIF x = 5020 THEN
            sigmoid_f := 1885;
        ELSIF x = 5021 THEN
            sigmoid_f := 1885;
        ELSIF x = 5022 THEN
            sigmoid_f := 1885;
        ELSIF x = 5023 THEN
            sigmoid_f := 1885;
        ELSIF x = 5024 THEN
            sigmoid_f := 1885;
        ELSIF x = 5025 THEN
            sigmoid_f := 1886;
        ELSIF x = 5026 THEN
            sigmoid_f := 1886;
        ELSIF x = 5027 THEN
            sigmoid_f := 1886;
        ELSIF x = 5028 THEN
            sigmoid_f := 1886;
        ELSIF x = 5029 THEN
            sigmoid_f := 1886;
        ELSIF x = 5030 THEN
            sigmoid_f := 1886;
        ELSIF x = 5031 THEN
            sigmoid_f := 1886;
        ELSIF x = 5032 THEN
            sigmoid_f := 1886;
        ELSIF x = 5033 THEN
            sigmoid_f := 1886;
        ELSIF x = 5034 THEN
            sigmoid_f := 1886;
        ELSIF x = 5035 THEN
            sigmoid_f := 1886;
        ELSIF x = 5036 THEN
            sigmoid_f := 1886;
        ELSIF x = 5037 THEN
            sigmoid_f := 1886;
        ELSIF x = 5038 THEN
            sigmoid_f := 1887;
        ELSIF x = 5039 THEN
            sigmoid_f := 1887;
        ELSIF x = 5040 THEN
            sigmoid_f := 1887;
        ELSIF x = 5041 THEN
            sigmoid_f := 1887;
        ELSIF x = 5042 THEN
            sigmoid_f := 1887;
        ELSIF x = 5043 THEN
            sigmoid_f := 1887;
        ELSIF x = 5044 THEN
            sigmoid_f := 1887;
        ELSIF x = 5045 THEN
            sigmoid_f := 1887;
        ELSIF x = 5046 THEN
            sigmoid_f := 1887;
        ELSIF x = 5047 THEN
            sigmoid_f := 1887;
        ELSIF x = 5048 THEN
            sigmoid_f := 1887;
        ELSIF x = 5049 THEN
            sigmoid_f := 1887;
        ELSIF x = 5050 THEN
            sigmoid_f := 1887;
        ELSIF x = 5051 THEN
            sigmoid_f := 1888;
        ELSIF x = 5052 THEN
            sigmoid_f := 1888;
        ELSIF x = 5053 THEN
            sigmoid_f := 1888;
        ELSIF x = 5054 THEN
            sigmoid_f := 1888;
        ELSIF x = 5055 THEN
            sigmoid_f := 1888;
        ELSIF x = 5056 THEN
            sigmoid_f := 1888;
        ELSIF x = 5057 THEN
            sigmoid_f := 1888;
        ELSIF x = 5058 THEN
            sigmoid_f := 1888;
        ELSIF x = 5059 THEN
            sigmoid_f := 1888;
        ELSIF x = 5060 THEN
            sigmoid_f := 1888;
        ELSIF x = 5061 THEN
            sigmoid_f := 1888;
        ELSIF x = 5062 THEN
            sigmoid_f := 1888;
        ELSIF x = 5063 THEN
            sigmoid_f := 1889;
        ELSIF x = 5064 THEN
            sigmoid_f := 1889;
        ELSIF x = 5065 THEN
            sigmoid_f := 1889;
        ELSIF x = 5066 THEN
            sigmoid_f := 1889;
        ELSIF x = 5067 THEN
            sigmoid_f := 1889;
        ELSIF x = 5068 THEN
            sigmoid_f := 1889;
        ELSIF x = 5069 THEN
            sigmoid_f := 1889;
        ELSIF x = 5070 THEN
            sigmoid_f := 1889;
        ELSIF x = 5071 THEN
            sigmoid_f := 1889;
        ELSIF x = 5072 THEN
            sigmoid_f := 1889;
        ELSIF x = 5073 THEN
            sigmoid_f := 1889;
        ELSIF x = 5074 THEN
            sigmoid_f := 1889;
        ELSIF x = 5075 THEN
            sigmoid_f := 1889;
        ELSIF x = 5076 THEN
            sigmoid_f := 1890;
        ELSIF x = 5077 THEN
            sigmoid_f := 1890;
        ELSIF x = 5078 THEN
            sigmoid_f := 1890;
        ELSIF x = 5079 THEN
            sigmoid_f := 1890;
        ELSIF x = 5080 THEN
            sigmoid_f := 1890;
        ELSIF x = 5081 THEN
            sigmoid_f := 1890;
        ELSIF x = 5082 THEN
            sigmoid_f := 1890;
        ELSIF x = 5083 THEN
            sigmoid_f := 1890;
        ELSIF x = 5084 THEN
            sigmoid_f := 1890;
        ELSIF x = 5085 THEN
            sigmoid_f := 1890;
        ELSIF x = 5086 THEN
            sigmoid_f := 1890;
        ELSIF x = 5087 THEN
            sigmoid_f := 1890;
        ELSIF x = 5088 THEN
            sigmoid_f := 1890;
        ELSIF x = 5089 THEN
            sigmoid_f := 1891;
        ELSIF x = 5090 THEN
            sigmoid_f := 1891;
        ELSIF x = 5091 THEN
            sigmoid_f := 1891;
        ELSIF x = 5092 THEN
            sigmoid_f := 1891;
        ELSIF x = 5093 THEN
            sigmoid_f := 1891;
        ELSIF x = 5094 THEN
            sigmoid_f := 1891;
        ELSIF x = 5095 THEN
            sigmoid_f := 1891;
        ELSIF x = 5096 THEN
            sigmoid_f := 1891;
        ELSIF x = 5097 THEN
            sigmoid_f := 1891;
        ELSIF x = 5098 THEN
            sigmoid_f := 1891;
        ELSIF x = 5099 THEN
            sigmoid_f := 1891;
        ELSIF x = 5100 THEN
            sigmoid_f := 1891;
        ELSIF x = 5101 THEN
            sigmoid_f := 1892;
        ELSIF x = 5102 THEN
            sigmoid_f := 1892;
        ELSIF x = 5103 THEN
            sigmoid_f := 1892;
        ELSIF x = 5104 THEN
            sigmoid_f := 1892;
        ELSIF x = 5105 THEN
            sigmoid_f := 1892;
        ELSIF x = 5106 THEN
            sigmoid_f := 1892;
        ELSIF x = 5107 THEN
            sigmoid_f := 1892;
        ELSIF x = 5108 THEN
            sigmoid_f := 1892;
        ELSIF x = 5109 THEN
            sigmoid_f := 1892;
        ELSIF x = 5110 THEN
            sigmoid_f := 1892;
        ELSIF x = 5111 THEN
            sigmoid_f := 1892;
        ELSIF x = 5112 THEN
            sigmoid_f := 1892;
        ELSIF x = 5113 THEN
            sigmoid_f := 1892;
        ELSIF x = 5114 THEN
            sigmoid_f := 1893;
        ELSIF x = 5115 THEN
            sigmoid_f := 1893;
        ELSIF x = 5116 THEN
            sigmoid_f := 1893;
        ELSIF x = 5117 THEN
            sigmoid_f := 1893;
        ELSIF x = 5118 THEN
            sigmoid_f := 1893;
        ELSIF x = 5119 THEN
            sigmoid_f := 1893;
        ELSIF x = 5120 THEN
            sigmoid_f := 1893;
        ELSIF x = 5121 THEN
            sigmoid_f := 1893;
        ELSIF x = 5122 THEN
            sigmoid_f := 1893;
        ELSIF x = 5123 THEN
            sigmoid_f := 1893;
        ELSIF x = 5124 THEN
            sigmoid_f := 1893;
        ELSIF x = 5125 THEN
            sigmoid_f := 1893;
        ELSIF x = 5126 THEN
            sigmoid_f := 1893;
        ELSIF x = 5127 THEN
            sigmoid_f := 1893;
        ELSIF x = 5128 THEN
            sigmoid_f := 1893;
        ELSIF x = 5129 THEN
            sigmoid_f := 1894;
        ELSIF x = 5130 THEN
            sigmoid_f := 1894;
        ELSIF x = 5131 THEN
            sigmoid_f := 1894;
        ELSIF x = 5132 THEN
            sigmoid_f := 1894;
        ELSIF x = 5133 THEN
            sigmoid_f := 1894;
        ELSIF x = 5134 THEN
            sigmoid_f := 1894;
        ELSIF x = 5135 THEN
            sigmoid_f := 1894;
        ELSIF x = 5136 THEN
            sigmoid_f := 1894;
        ELSIF x = 5137 THEN
            sigmoid_f := 1894;
        ELSIF x = 5138 THEN
            sigmoid_f := 1894;
        ELSIF x = 5139 THEN
            sigmoid_f := 1894;
        ELSIF x = 5140 THEN
            sigmoid_f := 1894;
        ELSIF x = 5141 THEN
            sigmoid_f := 1894;
        ELSIF x = 5142 THEN
            sigmoid_f := 1894;
        ELSIF x = 5143 THEN
            sigmoid_f := 1894;
        ELSIF x = 5144 THEN
            sigmoid_f := 1894;
        ELSIF x = 5145 THEN
            sigmoid_f := 1895;
        ELSIF x = 5146 THEN
            sigmoid_f := 1895;
        ELSIF x = 5147 THEN
            sigmoid_f := 1895;
        ELSIF x = 5148 THEN
            sigmoid_f := 1895;
        ELSIF x = 5149 THEN
            sigmoid_f := 1895;
        ELSIF x = 5150 THEN
            sigmoid_f := 1895;
        ELSIF x = 5151 THEN
            sigmoid_f := 1895;
        ELSIF x = 5152 THEN
            sigmoid_f := 1895;
        ELSIF x = 5153 THEN
            sigmoid_f := 1895;
        ELSIF x = 5154 THEN
            sigmoid_f := 1895;
        ELSIF x = 5155 THEN
            sigmoid_f := 1895;
        ELSIF x = 5156 THEN
            sigmoid_f := 1895;
        ELSIF x = 5157 THEN
            sigmoid_f := 1895;
        ELSIF x = 5158 THEN
            sigmoid_f := 1895;
        ELSIF x = 5159 THEN
            sigmoid_f := 1895;
        ELSIF x = 5160 THEN
            sigmoid_f := 1895;
        ELSIF x = 5161 THEN
            sigmoid_f := 1896;
        ELSIF x = 5162 THEN
            sigmoid_f := 1896;
        ELSIF x = 5163 THEN
            sigmoid_f := 1896;
        ELSIF x = 5164 THEN
            sigmoid_f := 1896;
        ELSIF x = 5165 THEN
            sigmoid_f := 1896;
        ELSIF x = 5166 THEN
            sigmoid_f := 1896;
        ELSIF x = 5167 THEN
            sigmoid_f := 1896;
        ELSIF x = 5168 THEN
            sigmoid_f := 1896;
        ELSIF x = 5169 THEN
            sigmoid_f := 1896;
        ELSIF x = 5170 THEN
            sigmoid_f := 1896;
        ELSIF x = 5171 THEN
            sigmoid_f := 1896;
        ELSIF x = 5172 THEN
            sigmoid_f := 1896;
        ELSIF x = 5173 THEN
            sigmoid_f := 1896;
        ELSIF x = 5174 THEN
            sigmoid_f := 1896;
        ELSIF x = 5175 THEN
            sigmoid_f := 1896;
        ELSIF x = 5176 THEN
            sigmoid_f := 1896;
        ELSIF x = 5177 THEN
            sigmoid_f := 1897;
        ELSIF x = 5178 THEN
            sigmoid_f := 1897;
        ELSIF x = 5179 THEN
            sigmoid_f := 1897;
        ELSIF x = 5180 THEN
            sigmoid_f := 1897;
        ELSIF x = 5181 THEN
            sigmoid_f := 1897;
        ELSIF x = 5182 THEN
            sigmoid_f := 1897;
        ELSIF x = 5183 THEN
            sigmoid_f := 1897;
        ELSIF x = 5184 THEN
            sigmoid_f := 1897;
        ELSIF x = 5185 THEN
            sigmoid_f := 1897;
        ELSIF x = 5186 THEN
            sigmoid_f := 1897;
        ELSIF x = 5187 THEN
            sigmoid_f := 1897;
        ELSIF x = 5188 THEN
            sigmoid_f := 1897;
        ELSIF x = 5189 THEN
            sigmoid_f := 1897;
        ELSIF x = 5190 THEN
            sigmoid_f := 1897;
        ELSIF x = 5191 THEN
            sigmoid_f := 1897;
        ELSIF x = 5192 THEN
            sigmoid_f := 1897;
        ELSIF x = 5193 THEN
            sigmoid_f := 1898;
        ELSIF x = 5194 THEN
            sigmoid_f := 1898;
        ELSIF x = 5195 THEN
            sigmoid_f := 1898;
        ELSIF x = 5196 THEN
            sigmoid_f := 1898;
        ELSIF x = 5197 THEN
            sigmoid_f := 1898;
        ELSIF x = 5198 THEN
            sigmoid_f := 1898;
        ELSIF x = 5199 THEN
            sigmoid_f := 1898;
        ELSIF x = 5200 THEN
            sigmoid_f := 1898;
        ELSIF x = 5201 THEN
            sigmoid_f := 1898;
        ELSIF x = 5202 THEN
            sigmoid_f := 1898;
        ELSIF x = 5203 THEN
            sigmoid_f := 1898;
        ELSIF x = 5204 THEN
            sigmoid_f := 1898;
        ELSIF x = 5205 THEN
            sigmoid_f := 1898;
        ELSIF x = 5206 THEN
            sigmoid_f := 1898;
        ELSIF x = 5207 THEN
            sigmoid_f := 1898;
        ELSIF x = 5208 THEN
            sigmoid_f := 1898;
        ELSIF x = 5209 THEN
            sigmoid_f := 1899;
        ELSIF x = 5210 THEN
            sigmoid_f := 1899;
        ELSIF x = 5211 THEN
            sigmoid_f := 1899;
        ELSIF x = 5212 THEN
            sigmoid_f := 1899;
        ELSIF x = 5213 THEN
            sigmoid_f := 1899;
        ELSIF x = 5214 THEN
            sigmoid_f := 1899;
        ELSIF x = 5215 THEN
            sigmoid_f := 1899;
        ELSIF x = 5216 THEN
            sigmoid_f := 1899;
        ELSIF x = 5217 THEN
            sigmoid_f := 1899;
        ELSIF x = 5218 THEN
            sigmoid_f := 1899;
        ELSIF x = 5219 THEN
            sigmoid_f := 1899;
        ELSIF x = 5220 THEN
            sigmoid_f := 1899;
        ELSIF x = 5221 THEN
            sigmoid_f := 1899;
        ELSIF x = 5222 THEN
            sigmoid_f := 1899;
        ELSIF x = 5223 THEN
            sigmoid_f := 1899;
        ELSIF x = 5224 THEN
            sigmoid_f := 1899;
        ELSIF x = 5225 THEN
            sigmoid_f := 1900;
        ELSIF x = 5226 THEN
            sigmoid_f := 1900;
        ELSIF x = 5227 THEN
            sigmoid_f := 1900;
        ELSIF x = 5228 THEN
            sigmoid_f := 1900;
        ELSIF x = 5229 THEN
            sigmoid_f := 1900;
        ELSIF x = 5230 THEN
            sigmoid_f := 1900;
        ELSIF x = 5231 THEN
            sigmoid_f := 1900;
        ELSIF x = 5232 THEN
            sigmoid_f := 1900;
        ELSIF x = 5233 THEN
            sigmoid_f := 1900;
        ELSIF x = 5234 THEN
            sigmoid_f := 1900;
        ELSIF x = 5235 THEN
            sigmoid_f := 1900;
        ELSIF x = 5236 THEN
            sigmoid_f := 1900;
        ELSIF x = 5237 THEN
            sigmoid_f := 1900;
        ELSIF x = 5238 THEN
            sigmoid_f := 1900;
        ELSIF x = 5239 THEN
            sigmoid_f := 1900;
        ELSIF x = 5240 THEN
            sigmoid_f := 1900;
        ELSIF x = 5241 THEN
            sigmoid_f := 1901;
        ELSIF x = 5242 THEN
            sigmoid_f := 1901;
        ELSIF x = 5243 THEN
            sigmoid_f := 1901;
        ELSIF x = 5244 THEN
            sigmoid_f := 1901;
        ELSIF x = 5245 THEN
            sigmoid_f := 1901;
        ELSIF x = 5246 THEN
            sigmoid_f := 1901;
        ELSIF x = 5247 THEN
            sigmoid_f := 1901;
        ELSIF x = 5248 THEN
            sigmoid_f := 1901;
        ELSIF x = 5249 THEN
            sigmoid_f := 1901;
        ELSIF x = 5250 THEN
            sigmoid_f := 1901;
        ELSIF x = 5251 THEN
            sigmoid_f := 1901;
        ELSIF x = 5252 THEN
            sigmoid_f := 1901;
        ELSIF x = 5253 THEN
            sigmoid_f := 1901;
        ELSIF x = 5254 THEN
            sigmoid_f := 1901;
        ELSIF x = 5255 THEN
            sigmoid_f := 1901;
        ELSIF x = 5256 THEN
            sigmoid_f := 1901;
        ELSIF x = 5257 THEN
            sigmoid_f := 1901;
        ELSIF x = 5258 THEN
            sigmoid_f := 1902;
        ELSIF x = 5259 THEN
            sigmoid_f := 1902;
        ELSIF x = 5260 THEN
            sigmoid_f := 1902;
        ELSIF x = 5261 THEN
            sigmoid_f := 1902;
        ELSIF x = 5262 THEN
            sigmoid_f := 1902;
        ELSIF x = 5263 THEN
            sigmoid_f := 1902;
        ELSIF x = 5264 THEN
            sigmoid_f := 1902;
        ELSIF x = 5265 THEN
            sigmoid_f := 1902;
        ELSIF x = 5266 THEN
            sigmoid_f := 1902;
        ELSIF x = 5267 THEN
            sigmoid_f := 1902;
        ELSIF x = 5268 THEN
            sigmoid_f := 1902;
        ELSIF x = 5269 THEN
            sigmoid_f := 1902;
        ELSIF x = 5270 THEN
            sigmoid_f := 1902;
        ELSIF x = 5271 THEN
            sigmoid_f := 1902;
        ELSIF x = 5272 THEN
            sigmoid_f := 1902;
        ELSIF x = 5273 THEN
            sigmoid_f := 1902;
        ELSIF x = 5274 THEN
            sigmoid_f := 1903;
        ELSIF x = 5275 THEN
            sigmoid_f := 1903;
        ELSIF x = 5276 THEN
            sigmoid_f := 1903;
        ELSIF x = 5277 THEN
            sigmoid_f := 1903;
        ELSIF x = 5278 THEN
            sigmoid_f := 1903;
        ELSIF x = 5279 THEN
            sigmoid_f := 1903;
        ELSIF x = 5280 THEN
            sigmoid_f := 1903;
        ELSIF x = 5281 THEN
            sigmoid_f := 1903;
        ELSIF x = 5282 THEN
            sigmoid_f := 1903;
        ELSIF x = 5283 THEN
            sigmoid_f := 1903;
        ELSIF x = 5284 THEN
            sigmoid_f := 1903;
        ELSIF x = 5285 THEN
            sigmoid_f := 1903;
        ELSIF x = 5286 THEN
            sigmoid_f := 1903;
        ELSIF x = 5287 THEN
            sigmoid_f := 1903;
        ELSIF x = 5288 THEN
            sigmoid_f := 1903;
        ELSIF x = 5289 THEN
            sigmoid_f := 1903;
        ELSIF x = 5290 THEN
            sigmoid_f := 1904;
        ELSIF x = 5291 THEN
            sigmoid_f := 1904;
        ELSIF x = 5292 THEN
            sigmoid_f := 1904;
        ELSIF x = 5293 THEN
            sigmoid_f := 1904;
        ELSIF x = 5294 THEN
            sigmoid_f := 1904;
        ELSIF x = 5295 THEN
            sigmoid_f := 1904;
        ELSIF x = 5296 THEN
            sigmoid_f := 1904;
        ELSIF x = 5297 THEN
            sigmoid_f := 1904;
        ELSIF x = 5298 THEN
            sigmoid_f := 1904;
        ELSIF x = 5299 THEN
            sigmoid_f := 1904;
        ELSIF x = 5300 THEN
            sigmoid_f := 1904;
        ELSIF x = 5301 THEN
            sigmoid_f := 1904;
        ELSIF x = 5302 THEN
            sigmoid_f := 1904;
        ELSIF x = 5303 THEN
            sigmoid_f := 1904;
        ELSIF x = 5304 THEN
            sigmoid_f := 1904;
        ELSIF x = 5305 THEN
            sigmoid_f := 1904;
        ELSIF x = 5306 THEN
            sigmoid_f := 1905;
        ELSIF x = 5307 THEN
            sigmoid_f := 1905;
        ELSIF x = 5308 THEN
            sigmoid_f := 1905;
        ELSIF x = 5309 THEN
            sigmoid_f := 1905;
        ELSIF x = 5310 THEN
            sigmoid_f := 1905;
        ELSIF x = 5311 THEN
            sigmoid_f := 1905;
        ELSIF x = 5312 THEN
            sigmoid_f := 1905;
        ELSIF x = 5313 THEN
            sigmoid_f := 1905;
        ELSIF x = 5314 THEN
            sigmoid_f := 1905;
        ELSIF x = 5315 THEN
            sigmoid_f := 1905;
        ELSIF x = 5316 THEN
            sigmoid_f := 1905;
        ELSIF x = 5317 THEN
            sigmoid_f := 1905;
        ELSIF x = 5318 THEN
            sigmoid_f := 1905;
        ELSIF x = 5319 THEN
            sigmoid_f := 1905;
        ELSIF x = 5320 THEN
            sigmoid_f := 1905;
        ELSIF x = 5321 THEN
            sigmoid_f := 1905;
        ELSIF x = 5322 THEN
            sigmoid_f := 1906;
        ELSIF x = 5323 THEN
            sigmoid_f := 1906;
        ELSIF x = 5324 THEN
            sigmoid_f := 1906;
        ELSIF x = 5325 THEN
            sigmoid_f := 1906;
        ELSIF x = 5326 THEN
            sigmoid_f := 1906;
        ELSIF x = 5327 THEN
            sigmoid_f := 1906;
        ELSIF x = 5328 THEN
            sigmoid_f := 1906;
        ELSIF x = 5329 THEN
            sigmoid_f := 1906;
        ELSIF x = 5330 THEN
            sigmoid_f := 1906;
        ELSIF x = 5331 THEN
            sigmoid_f := 1906;
        ELSIF x = 5332 THEN
            sigmoid_f := 1906;
        ELSIF x = 5333 THEN
            sigmoid_f := 1906;
        ELSIF x = 5334 THEN
            sigmoid_f := 1906;
        ELSIF x = 5335 THEN
            sigmoid_f := 1906;
        ELSIF x = 5336 THEN
            sigmoid_f := 1906;
        ELSIF x = 5337 THEN
            sigmoid_f := 1906;
        ELSIF x = 5338 THEN
            sigmoid_f := 1907;
        ELSIF x = 5339 THEN
            sigmoid_f := 1907;
        ELSIF x = 5340 THEN
            sigmoid_f := 1907;
        ELSIF x = 5341 THEN
            sigmoid_f := 1907;
        ELSIF x = 5342 THEN
            sigmoid_f := 1907;
        ELSIF x = 5343 THEN
            sigmoid_f := 1907;
        ELSIF x = 5344 THEN
            sigmoid_f := 1907;
        ELSIF x = 5345 THEN
            sigmoid_f := 1907;
        ELSIF x = 5346 THEN
            sigmoid_f := 1907;
        ELSIF x = 5347 THEN
            sigmoid_f := 1907;
        ELSIF x = 5348 THEN
            sigmoid_f := 1907;
        ELSIF x = 5349 THEN
            sigmoid_f := 1907;
        ELSIF x = 5350 THEN
            sigmoid_f := 1907;
        ELSIF x = 5351 THEN
            sigmoid_f := 1907;
        ELSIF x = 5352 THEN
            sigmoid_f := 1907;
        ELSIF x = 5353 THEN
            sigmoid_f := 1907;
        ELSIF x = 5354 THEN
            sigmoid_f := 1908;
        ELSIF x = 5355 THEN
            sigmoid_f := 1908;
        ELSIF x = 5356 THEN
            sigmoid_f := 1908;
        ELSIF x = 5357 THEN
            sigmoid_f := 1908;
        ELSIF x = 5358 THEN
            sigmoid_f := 1908;
        ELSIF x = 5359 THEN
            sigmoid_f := 1908;
        ELSIF x = 5360 THEN
            sigmoid_f := 1908;
        ELSIF x = 5361 THEN
            sigmoid_f := 1908;
        ELSIF x = 5362 THEN
            sigmoid_f := 1908;
        ELSIF x = 5363 THEN
            sigmoid_f := 1908;
        ELSIF x = 5364 THEN
            sigmoid_f := 1908;
        ELSIF x = 5365 THEN
            sigmoid_f := 1908;
        ELSIF x = 5366 THEN
            sigmoid_f := 1908;
        ELSIF x = 5367 THEN
            sigmoid_f := 1908;
        ELSIF x = 5368 THEN
            sigmoid_f := 1908;
        ELSIF x = 5369 THEN
            sigmoid_f := 1908;
        ELSIF x = 5370 THEN
            sigmoid_f := 1909;
        ELSIF x = 5371 THEN
            sigmoid_f := 1909;
        ELSIF x = 5372 THEN
            sigmoid_f := 1909;
        ELSIF x = 5373 THEN
            sigmoid_f := 1909;
        ELSIF x = 5374 THEN
            sigmoid_f := 1909;
        ELSIF x = 5375 THEN
            sigmoid_f := 1909;
        ELSIF x = 5376 THEN
            sigmoid_f := 1909;
        ELSIF x = 5377 THEN
            sigmoid_f := 1909;
        ELSIF x = 5378 THEN
            sigmoid_f := 1909;
        ELSIF x = 5379 THEN
            sigmoid_f := 1909;
        ELSIF x = 5380 THEN
            sigmoid_f := 1909;
        ELSIF x = 5381 THEN
            sigmoid_f := 1909;
        ELSIF x = 5382 THEN
            sigmoid_f := 1909;
        ELSIF x = 5383 THEN
            sigmoid_f := 1909;
        ELSIF x = 5384 THEN
            sigmoid_f := 1909;
        ELSIF x = 5385 THEN
            sigmoid_f := 1909;
        ELSIF x = 5386 THEN
            sigmoid_f := 1909;
        ELSIF x = 5387 THEN
            sigmoid_f := 1910;
        ELSIF x = 5388 THEN
            sigmoid_f := 1910;
        ELSIF x = 5389 THEN
            sigmoid_f := 1910;
        ELSIF x = 5390 THEN
            sigmoid_f := 1910;
        ELSIF x = 5391 THEN
            sigmoid_f := 1910;
        ELSIF x = 5392 THEN
            sigmoid_f := 1910;
        ELSIF x = 5393 THEN
            sigmoid_f := 1910;
        ELSIF x = 5394 THEN
            sigmoid_f := 1910;
        ELSIF x = 5395 THEN
            sigmoid_f := 1910;
        ELSIF x = 5396 THEN
            sigmoid_f := 1910;
        ELSIF x = 5397 THEN
            sigmoid_f := 1910;
        ELSIF x = 5398 THEN
            sigmoid_f := 1910;
        ELSIF x = 5399 THEN
            sigmoid_f := 1910;
        ELSIF x = 5400 THEN
            sigmoid_f := 1910;
        ELSIF x = 5401 THEN
            sigmoid_f := 1910;
        ELSIF x = 5402 THEN
            sigmoid_f := 1910;
        ELSIF x = 5403 THEN
            sigmoid_f := 1911;
        ELSIF x = 5404 THEN
            sigmoid_f := 1911;
        ELSIF x = 5405 THEN
            sigmoid_f := 1911;
        ELSIF x = 5406 THEN
            sigmoid_f := 1911;
        ELSIF x = 5407 THEN
            sigmoid_f := 1911;
        ELSIF x = 5408 THEN
            sigmoid_f := 1911;
        ELSIF x = 5409 THEN
            sigmoid_f := 1911;
        ELSIF x = 5410 THEN
            sigmoid_f := 1911;
        ELSIF x = 5411 THEN
            sigmoid_f := 1911;
        ELSIF x = 5412 THEN
            sigmoid_f := 1911;
        ELSIF x = 5413 THEN
            sigmoid_f := 1911;
        ELSIF x = 5414 THEN
            sigmoid_f := 1911;
        ELSIF x = 5415 THEN
            sigmoid_f := 1911;
        ELSIF x = 5416 THEN
            sigmoid_f := 1911;
        ELSIF x = 5417 THEN
            sigmoid_f := 1911;
        ELSIF x = 5418 THEN
            sigmoid_f := 1911;
        ELSIF x = 5419 THEN
            sigmoid_f := 1912;
        ELSIF x = 5420 THEN
            sigmoid_f := 1912;
        ELSIF x = 5421 THEN
            sigmoid_f := 1912;
        ELSIF x = 5422 THEN
            sigmoid_f := 1912;
        ELSIF x = 5423 THEN
            sigmoid_f := 1912;
        ELSIF x = 5424 THEN
            sigmoid_f := 1912;
        ELSIF x = 5425 THEN
            sigmoid_f := 1912;
        ELSIF x = 5426 THEN
            sigmoid_f := 1912;
        ELSIF x = 5427 THEN
            sigmoid_f := 1912;
        ELSIF x = 5428 THEN
            sigmoid_f := 1912;
        ELSIF x = 5429 THEN
            sigmoid_f := 1912;
        ELSIF x = 5430 THEN
            sigmoid_f := 1912;
        ELSIF x = 5431 THEN
            sigmoid_f := 1912;
        ELSIF x = 5432 THEN
            sigmoid_f := 1912;
        ELSIF x = 5433 THEN
            sigmoid_f := 1912;
        ELSIF x = 5434 THEN
            sigmoid_f := 1912;
        ELSIF x = 5435 THEN
            sigmoid_f := 1913;
        ELSIF x = 5436 THEN
            sigmoid_f := 1913;
        ELSIF x = 5437 THEN
            sigmoid_f := 1913;
        ELSIF x = 5438 THEN
            sigmoid_f := 1913;
        ELSIF x = 5439 THEN
            sigmoid_f := 1913;
        ELSIF x = 5440 THEN
            sigmoid_f := 1913;
        ELSIF x = 5441 THEN
            sigmoid_f := 1913;
        ELSIF x = 5442 THEN
            sigmoid_f := 1913;
        ELSIF x = 5443 THEN
            sigmoid_f := 1913;
        ELSIF x = 5444 THEN
            sigmoid_f := 1913;
        ELSIF x = 5445 THEN
            sigmoid_f := 1913;
        ELSIF x = 5446 THEN
            sigmoid_f := 1913;
        ELSIF x = 5447 THEN
            sigmoid_f := 1913;
        ELSIF x = 5448 THEN
            sigmoid_f := 1913;
        ELSIF x = 5449 THEN
            sigmoid_f := 1913;
        ELSIF x = 5450 THEN
            sigmoid_f := 1913;
        ELSIF x = 5451 THEN
            sigmoid_f := 1914;
        ELSIF x = 5452 THEN
            sigmoid_f := 1914;
        ELSIF x = 5453 THEN
            sigmoid_f := 1914;
        ELSIF x = 5454 THEN
            sigmoid_f := 1914;
        ELSIF x = 5455 THEN
            sigmoid_f := 1914;
        ELSIF x = 5456 THEN
            sigmoid_f := 1914;
        ELSIF x = 5457 THEN
            sigmoid_f := 1914;
        ELSIF x = 5458 THEN
            sigmoid_f := 1914;
        ELSIF x = 5459 THEN
            sigmoid_f := 1914;
        ELSIF x = 5460 THEN
            sigmoid_f := 1914;
        ELSIF x = 5461 THEN
            sigmoid_f := 1914;
        ELSIF x = 5462 THEN
            sigmoid_f := 1914;
        ELSIF x = 5463 THEN
            sigmoid_f := 1914;
        ELSIF x = 5464 THEN
            sigmoid_f := 1914;
        ELSIF x = 5465 THEN
            sigmoid_f := 1914;
        ELSIF x = 5466 THEN
            sigmoid_f := 1914;
        ELSIF x = 5467 THEN
            sigmoid_f := 1915;
        ELSIF x = 5468 THEN
            sigmoid_f := 1915;
        ELSIF x = 5469 THEN
            sigmoid_f := 1915;
        ELSIF x = 5470 THEN
            sigmoid_f := 1915;
        ELSIF x = 5471 THEN
            sigmoid_f := 1915;
        ELSIF x = 5472 THEN
            sigmoid_f := 1915;
        ELSIF x = 5473 THEN
            sigmoid_f := 1915;
        ELSIF x = 5474 THEN
            sigmoid_f := 1915;
        ELSIF x = 5475 THEN
            sigmoid_f := 1915;
        ELSIF x = 5476 THEN
            sigmoid_f := 1915;
        ELSIF x = 5477 THEN
            sigmoid_f := 1915;
        ELSIF x = 5478 THEN
            sigmoid_f := 1915;
        ELSIF x = 5479 THEN
            sigmoid_f := 1915;
        ELSIF x = 5480 THEN
            sigmoid_f := 1915;
        ELSIF x = 5481 THEN
            sigmoid_f := 1915;
        ELSIF x = 5482 THEN
            sigmoid_f := 1915;
        ELSIF x = 5483 THEN
            sigmoid_f := 1916;
        ELSIF x = 5484 THEN
            sigmoid_f := 1916;
        ELSIF x = 5485 THEN
            sigmoid_f := 1916;
        ELSIF x = 5486 THEN
            sigmoid_f := 1916;
        ELSIF x = 5487 THEN
            sigmoid_f := 1916;
        ELSIF x = 5488 THEN
            sigmoid_f := 1916;
        ELSIF x = 5489 THEN
            sigmoid_f := 1916;
        ELSIF x = 5490 THEN
            sigmoid_f := 1916;
        ELSIF x = 5491 THEN
            sigmoid_f := 1916;
        ELSIF x = 5492 THEN
            sigmoid_f := 1916;
        ELSIF x = 5493 THEN
            sigmoid_f := 1916;
        ELSIF x = 5494 THEN
            sigmoid_f := 1916;
        ELSIF x = 5495 THEN
            sigmoid_f := 1916;
        ELSIF x = 5496 THEN
            sigmoid_f := 1916;
        ELSIF x = 5497 THEN
            sigmoid_f := 1916;
        ELSIF x = 5498 THEN
            sigmoid_f := 1916;
        ELSIF x = 5499 THEN
            sigmoid_f := 1917;
        ELSIF x = 5500 THEN
            sigmoid_f := 1917;
        ELSIF x = 5501 THEN
            sigmoid_f := 1917;
        ELSIF x = 5502 THEN
            sigmoid_f := 1917;
        ELSIF x = 5503 THEN
            sigmoid_f := 1917;
        ELSIF x = 5504 THEN
            sigmoid_f := 1917;
        ELSIF x = 5505 THEN
            sigmoid_f := 1917;
        ELSIF x = 5506 THEN
            sigmoid_f := 1917;
        ELSIF x = 5507 THEN
            sigmoid_f := 1917;
        ELSIF x = 5508 THEN
            sigmoid_f := 1917;
        ELSIF x = 5509 THEN
            sigmoid_f := 1917;
        ELSIF x = 5510 THEN
            sigmoid_f := 1917;
        ELSIF x = 5511 THEN
            sigmoid_f := 1917;
        ELSIF x = 5512 THEN
            sigmoid_f := 1917;
        ELSIF x = 5513 THEN
            sigmoid_f := 1917;
        ELSIF x = 5514 THEN
            sigmoid_f := 1917;
        ELSIF x = 5515 THEN
            sigmoid_f := 1917;
        ELSIF x = 5516 THEN
            sigmoid_f := 1918;
        ELSIF x = 5517 THEN
            sigmoid_f := 1918;
        ELSIF x = 5518 THEN
            sigmoid_f := 1918;
        ELSIF x = 5519 THEN
            sigmoid_f := 1918;
        ELSIF x = 5520 THEN
            sigmoid_f := 1918;
        ELSIF x = 5521 THEN
            sigmoid_f := 1918;
        ELSIF x = 5522 THEN
            sigmoid_f := 1918;
        ELSIF x = 5523 THEN
            sigmoid_f := 1918;
        ELSIF x = 5524 THEN
            sigmoid_f := 1918;
        ELSIF x = 5525 THEN
            sigmoid_f := 1918;
        ELSIF x = 5526 THEN
            sigmoid_f := 1918;
        ELSIF x = 5527 THEN
            sigmoid_f := 1918;
        ELSIF x = 5528 THEN
            sigmoid_f := 1918;
        ELSIF x = 5529 THEN
            sigmoid_f := 1918;
        ELSIF x = 5530 THEN
            sigmoid_f := 1918;
        ELSIF x = 5531 THEN
            sigmoid_f := 1918;
        ELSIF x = 5532 THEN
            sigmoid_f := 1919;
        ELSIF x = 5533 THEN
            sigmoid_f := 1919;
        ELSIF x = 5534 THEN
            sigmoid_f := 1919;
        ELSIF x = 5535 THEN
            sigmoid_f := 1919;
        ELSIF x = 5536 THEN
            sigmoid_f := 1919;
        ELSIF x = 5537 THEN
            sigmoid_f := 1919;
        ELSIF x = 5538 THEN
            sigmoid_f := 1919;
        ELSIF x = 5539 THEN
            sigmoid_f := 1919;
        ELSIF x = 5540 THEN
            sigmoid_f := 1919;
        ELSIF x = 5541 THEN
            sigmoid_f := 1919;
        ELSIF x = 5542 THEN
            sigmoid_f := 1919;
        ELSIF x = 5543 THEN
            sigmoid_f := 1919;
        ELSIF x = 5544 THEN
            sigmoid_f := 1919;
        ELSIF x = 5545 THEN
            sigmoid_f := 1919;
        ELSIF x = 5546 THEN
            sigmoid_f := 1919;
        ELSIF x = 5547 THEN
            sigmoid_f := 1919;
        ELSIF x = 5548 THEN
            sigmoid_f := 1920;
        ELSIF x = 5549 THEN
            sigmoid_f := 1920;
        ELSIF x = 5550 THEN
            sigmoid_f := 1920;
        ELSIF x = 5551 THEN
            sigmoid_f := 1920;
        ELSIF x = 5552 THEN
            sigmoid_f := 1920;
        ELSIF x = 5553 THEN
            sigmoid_f := 1920;
        ELSIF x = 5554 THEN
            sigmoid_f := 1920;
        ELSIF x = 5555 THEN
            sigmoid_f := 1920;
        ELSIF x = 5556 THEN
            sigmoid_f := 1920;
        ELSIF x = 5557 THEN
            sigmoid_f := 1920;
        ELSIF x = 5558 THEN
            sigmoid_f := 1920;
        ELSIF x = 5559 THEN
            sigmoid_f := 1920;
        ELSIF x = 5560 THEN
            sigmoid_f := 1920;
        ELSIF x = 5561 THEN
            sigmoid_f := 1920;
        ELSIF x = 5562 THEN
            sigmoid_f := 1920;
        ELSIF x = 5563 THEN
            sigmoid_f := 1920;
        ELSIF x = 5564 THEN
            sigmoid_f := 1921;
        ELSIF x = 5565 THEN
            sigmoid_f := 1921;
        ELSIF x = 5566 THEN
            sigmoid_f := 1921;
        ELSIF x = 5567 THEN
            sigmoid_f := 1921;
        ELSIF x = 5568 THEN
            sigmoid_f := 1921;
        ELSIF x = 5569 THEN
            sigmoid_f := 1921;
        ELSIF x = 5570 THEN
            sigmoid_f := 1921;
        ELSIF x = 5571 THEN
            sigmoid_f := 1921;
        ELSIF x = 5572 THEN
            sigmoid_f := 1921;
        ELSIF x = 5573 THEN
            sigmoid_f := 1921;
        ELSIF x = 5574 THEN
            sigmoid_f := 1921;
        ELSIF x = 5575 THEN
            sigmoid_f := 1921;
        ELSIF x = 5576 THEN
            sigmoid_f := 1921;
        ELSIF x = 5577 THEN
            sigmoid_f := 1921;
        ELSIF x = 5578 THEN
            sigmoid_f := 1921;
        ELSIF x = 5579 THEN
            sigmoid_f := 1921;
        ELSIF x = 5580 THEN
            sigmoid_f := 1922;
        ELSIF x = 5581 THEN
            sigmoid_f := 1922;
        ELSIF x = 5582 THEN
            sigmoid_f := 1922;
        ELSIF x = 5583 THEN
            sigmoid_f := 1922;
        ELSIF x = 5584 THEN
            sigmoid_f := 1922;
        ELSIF x = 5585 THEN
            sigmoid_f := 1922;
        ELSIF x = 5586 THEN
            sigmoid_f := 1922;
        ELSIF x = 5587 THEN
            sigmoid_f := 1922;
        ELSIF x = 5588 THEN
            sigmoid_f := 1922;
        ELSIF x = 5589 THEN
            sigmoid_f := 1922;
        ELSIF x = 5590 THEN
            sigmoid_f := 1922;
        ELSIF x = 5591 THEN
            sigmoid_f := 1922;
        ELSIF x = 5592 THEN
            sigmoid_f := 1922;
        ELSIF x = 5593 THEN
            sigmoid_f := 1922;
        ELSIF x = 5594 THEN
            sigmoid_f := 1922;
        ELSIF x = 5595 THEN
            sigmoid_f := 1922;
        ELSIF x = 5596 THEN
            sigmoid_f := 1923;
        ELSIF x = 5597 THEN
            sigmoid_f := 1923;
        ELSIF x = 5598 THEN
            sigmoid_f := 1923;
        ELSIF x = 5599 THEN
            sigmoid_f := 1923;
        ELSIF x = 5600 THEN
            sigmoid_f := 1923;
        ELSIF x = 5601 THEN
            sigmoid_f := 1923;
        ELSIF x = 5602 THEN
            sigmoid_f := 1923;
        ELSIF x = 5603 THEN
            sigmoid_f := 1923;
        ELSIF x = 5604 THEN
            sigmoid_f := 1923;
        ELSIF x = 5605 THEN
            sigmoid_f := 1923;
        ELSIF x = 5606 THEN
            sigmoid_f := 1923;
        ELSIF x = 5607 THEN
            sigmoid_f := 1923;
        ELSIF x = 5608 THEN
            sigmoid_f := 1923;
        ELSIF x = 5609 THEN
            sigmoid_f := 1923;
        ELSIF x = 5610 THEN
            sigmoid_f := 1923;
        ELSIF x = 5611 THEN
            sigmoid_f := 1923;
        ELSIF x = 5612 THEN
            sigmoid_f := 1924;
        ELSIF x = 5613 THEN
            sigmoid_f := 1924;
        ELSIF x = 5614 THEN
            sigmoid_f := 1924;
        ELSIF x = 5615 THEN
            sigmoid_f := 1924;
        ELSIF x = 5616 THEN
            sigmoid_f := 1924;
        ELSIF x = 5617 THEN
            sigmoid_f := 1924;
        ELSIF x = 5618 THEN
            sigmoid_f := 1924;
        ELSIF x = 5619 THEN
            sigmoid_f := 1924;
        ELSIF x = 5620 THEN
            sigmoid_f := 1924;
        ELSIF x = 5621 THEN
            sigmoid_f := 1924;
        ELSIF x = 5622 THEN
            sigmoid_f := 1924;
        ELSIF x = 5623 THEN
            sigmoid_f := 1924;
        ELSIF x = 5624 THEN
            sigmoid_f := 1924;
        ELSIF x = 5625 THEN
            sigmoid_f := 1924;
        ELSIF x = 5626 THEN
            sigmoid_f := 1924;
        ELSIF x = 5627 THEN
            sigmoid_f := 1924;
        ELSIF x = 5628 THEN
            sigmoid_f := 1925;
        ELSIF x = 5629 THEN
            sigmoid_f := 1925;
        ELSIF x = 5630 THEN
            sigmoid_f := 1925;
        ELSIF x = 5631 THEN
            sigmoid_f := 1925;
        ELSIF x = 5632 THEN
            sigmoid_f := 1925;
        ELSIF x = 5633 THEN
            sigmoid_f := 1925;
        ELSIF x = 5634 THEN
            sigmoid_f := 1925;
        ELSIF x = 5635 THEN
            sigmoid_f := 1925;
        ELSIF x = 5636 THEN
            sigmoid_f := 1925;
        ELSIF x = 5637 THEN
            sigmoid_f := 1925;
        ELSIF x = 5638 THEN
            sigmoid_f := 1925;
        ELSIF x = 5639 THEN
            sigmoid_f := 1925;
        ELSIF x = 5640 THEN
            sigmoid_f := 1925;
        ELSIF x = 5641 THEN
            sigmoid_f := 1925;
        ELSIF x = 5642 THEN
            sigmoid_f := 1925;
        ELSIF x = 5643 THEN
            sigmoid_f := 1926;
        ELSIF x = 5644 THEN
            sigmoid_f := 1926;
        ELSIF x = 5645 THEN
            sigmoid_f := 1926;
        ELSIF x = 5646 THEN
            sigmoid_f := 1926;
        ELSIF x = 5647 THEN
            sigmoid_f := 1926;
        ELSIF x = 5648 THEN
            sigmoid_f := 1926;
        ELSIF x = 5649 THEN
            sigmoid_f := 1926;
        ELSIF x = 5650 THEN
            sigmoid_f := 1926;
        ELSIF x = 5651 THEN
            sigmoid_f := 1926;
        ELSIF x = 5652 THEN
            sigmoid_f := 1926;
        ELSIF x = 5653 THEN
            sigmoid_f := 1926;
        ELSIF x = 5654 THEN
            sigmoid_f := 1926;
        ELSIF x = 5655 THEN
            sigmoid_f := 1926;
        ELSIF x = 5656 THEN
            sigmoid_f := 1926;
        ELSIF x = 5657 THEN
            sigmoid_f := 1926;
        ELSIF x = 5658 THEN
            sigmoid_f := 1926;
        ELSIF x = 5659 THEN
            sigmoid_f := 1926;
        ELSIF x = 5660 THEN
            sigmoid_f := 1926;
        ELSIF x = 5661 THEN
            sigmoid_f := 1926;
        ELSIF x = 5662 THEN
            sigmoid_f := 1926;
        ELSIF x = 5663 THEN
            sigmoid_f := 1927;
        ELSIF x = 5664 THEN
            sigmoid_f := 1927;
        ELSIF x = 5665 THEN
            sigmoid_f := 1927;
        ELSIF x = 5666 THEN
            sigmoid_f := 1927;
        ELSIF x = 5667 THEN
            sigmoid_f := 1927;
        ELSIF x = 5668 THEN
            sigmoid_f := 1927;
        ELSIF x = 5669 THEN
            sigmoid_f := 1927;
        ELSIF x = 5670 THEN
            sigmoid_f := 1927;
        ELSIF x = 5671 THEN
            sigmoid_f := 1927;
        ELSIF x = 5672 THEN
            sigmoid_f := 1927;
        ELSIF x = 5673 THEN
            sigmoid_f := 1927;
        ELSIF x = 5674 THEN
            sigmoid_f := 1927;
        ELSIF x = 5675 THEN
            sigmoid_f := 1927;
        ELSIF x = 5676 THEN
            sigmoid_f := 1927;
        ELSIF x = 5677 THEN
            sigmoid_f := 1927;
        ELSIF x = 5678 THEN
            sigmoid_f := 1927;
        ELSIF x = 5679 THEN
            sigmoid_f := 1927;
        ELSIF x = 5680 THEN
            sigmoid_f := 1927;
        ELSIF x = 5681 THEN
            sigmoid_f := 1927;
        ELSIF x = 5682 THEN
            sigmoid_f := 1927;
        ELSIF x = 5683 THEN
            sigmoid_f := 1928;
        ELSIF x = 5684 THEN
            sigmoid_f := 1928;
        ELSIF x = 5685 THEN
            sigmoid_f := 1928;
        ELSIF x = 5686 THEN
            sigmoid_f := 1928;
        ELSIF x = 5687 THEN
            sigmoid_f := 1928;
        ELSIF x = 5688 THEN
            sigmoid_f := 1928;
        ELSIF x = 5689 THEN
            sigmoid_f := 1928;
        ELSIF x = 5690 THEN
            sigmoid_f := 1928;
        ELSIF x = 5691 THEN
            sigmoid_f := 1928;
        ELSIF x = 5692 THEN
            sigmoid_f := 1928;
        ELSIF x = 5693 THEN
            sigmoid_f := 1928;
        ELSIF x = 5694 THEN
            sigmoid_f := 1928;
        ELSIF x = 5695 THEN
            sigmoid_f := 1928;
        ELSIF x = 5696 THEN
            sigmoid_f := 1928;
        ELSIF x = 5697 THEN
            sigmoid_f := 1928;
        ELSIF x = 5698 THEN
            sigmoid_f := 1928;
        ELSIF x = 5699 THEN
            sigmoid_f := 1928;
        ELSIF x = 5700 THEN
            sigmoid_f := 1928;
        ELSIF x = 5701 THEN
            sigmoid_f := 1928;
        ELSIF x = 5702 THEN
            sigmoid_f := 1928;
        ELSIF x = 5703 THEN
            sigmoid_f := 1929;
        ELSIF x = 5704 THEN
            sigmoid_f := 1929;
        ELSIF x = 5705 THEN
            sigmoid_f := 1929;
        ELSIF x = 5706 THEN
            sigmoid_f := 1929;
        ELSIF x = 5707 THEN
            sigmoid_f := 1929;
        ELSIF x = 5708 THEN
            sigmoid_f := 1929;
        ELSIF x = 5709 THEN
            sigmoid_f := 1929;
        ELSIF x = 5710 THEN
            sigmoid_f := 1929;
        ELSIF x = 5711 THEN
            sigmoid_f := 1929;
        ELSIF x = 5712 THEN
            sigmoid_f := 1929;
        ELSIF x = 5713 THEN
            sigmoid_f := 1929;
        ELSIF x = 5714 THEN
            sigmoid_f := 1929;
        ELSIF x = 5715 THEN
            sigmoid_f := 1929;
        ELSIF x = 5716 THEN
            sigmoid_f := 1929;
        ELSIF x = 5717 THEN
            sigmoid_f := 1929;
        ELSIF x = 5718 THEN
            sigmoid_f := 1929;
        ELSIF x = 5719 THEN
            sigmoid_f := 1929;
        ELSIF x = 5720 THEN
            sigmoid_f := 1929;
        ELSIF x = 5721 THEN
            sigmoid_f := 1929;
        ELSIF x = 5722 THEN
            sigmoid_f := 1929;
        ELSIF x = 5723 THEN
            sigmoid_f := 1930;
        ELSIF x = 5724 THEN
            sigmoid_f := 1930;
        ELSIF x = 5725 THEN
            sigmoid_f := 1930;
        ELSIF x = 5726 THEN
            sigmoid_f := 1930;
        ELSIF x = 5727 THEN
            sigmoid_f := 1930;
        ELSIF x = 5728 THEN
            sigmoid_f := 1930;
        ELSIF x = 5729 THEN
            sigmoid_f := 1930;
        ELSIF x = 5730 THEN
            sigmoid_f := 1930;
        ELSIF x = 5731 THEN
            sigmoid_f := 1930;
        ELSIF x = 5732 THEN
            sigmoid_f := 1930;
        ELSIF x = 5733 THEN
            sigmoid_f := 1930;
        ELSIF x = 5734 THEN
            sigmoid_f := 1930;
        ELSIF x = 5735 THEN
            sigmoid_f := 1930;
        ELSIF x = 5736 THEN
            sigmoid_f := 1930;
        ELSIF x = 5737 THEN
            sigmoid_f := 1930;
        ELSIF x = 5738 THEN
            sigmoid_f := 1930;
        ELSIF x = 5739 THEN
            sigmoid_f := 1930;
        ELSIF x = 5740 THEN
            sigmoid_f := 1930;
        ELSIF x = 5741 THEN
            sigmoid_f := 1930;
        ELSIF x = 5742 THEN
            sigmoid_f := 1930;
        ELSIF x = 5743 THEN
            sigmoid_f := 1931;
        ELSIF x = 5744 THEN
            sigmoid_f := 1931;
        ELSIF x = 5745 THEN
            sigmoid_f := 1931;
        ELSIF x = 5746 THEN
            sigmoid_f := 1931;
        ELSIF x = 5747 THEN
            sigmoid_f := 1931;
        ELSIF x = 5748 THEN
            sigmoid_f := 1931;
        ELSIF x = 5749 THEN
            sigmoid_f := 1931;
        ELSIF x = 5750 THEN
            sigmoid_f := 1931;
        ELSIF x = 5751 THEN
            sigmoid_f := 1931;
        ELSIF x = 5752 THEN
            sigmoid_f := 1931;
        ELSIF x = 5753 THEN
            sigmoid_f := 1931;
        ELSIF x = 5754 THEN
            sigmoid_f := 1931;
        ELSIF x = 5755 THEN
            sigmoid_f := 1931;
        ELSIF x = 5756 THEN
            sigmoid_f := 1931;
        ELSIF x = 5757 THEN
            sigmoid_f := 1931;
        ELSIF x = 5758 THEN
            sigmoid_f := 1931;
        ELSIF x = 5759 THEN
            sigmoid_f := 1931;
        ELSIF x = 5760 THEN
            sigmoid_f := 1931;
        ELSIF x = 5761 THEN
            sigmoid_f := 1931;
        ELSIF x = 5762 THEN
            sigmoid_f := 1931;
        ELSIF x = 5763 THEN
            sigmoid_f := 1932;
        ELSIF x = 5764 THEN
            sigmoid_f := 1932;
        ELSIF x = 5765 THEN
            sigmoid_f := 1932;
        ELSIF x = 5766 THEN
            sigmoid_f := 1932;
        ELSIF x = 5767 THEN
            sigmoid_f := 1932;
        ELSIF x = 5768 THEN
            sigmoid_f := 1932;
        ELSIF x = 5769 THEN
            sigmoid_f := 1932;
        ELSIF x = 5770 THEN
            sigmoid_f := 1932;
        ELSIF x = 5771 THEN
            sigmoid_f := 1932;
        ELSIF x = 5772 THEN
            sigmoid_f := 1932;
        ELSIF x = 5773 THEN
            sigmoid_f := 1932;
        ELSIF x = 5774 THEN
            sigmoid_f := 1932;
        ELSIF x = 5775 THEN
            sigmoid_f := 1932;
        ELSIF x = 5776 THEN
            sigmoid_f := 1932;
        ELSIF x = 5777 THEN
            sigmoid_f := 1932;
        ELSIF x = 5778 THEN
            sigmoid_f := 1932;
        ELSIF x = 5779 THEN
            sigmoid_f := 1932;
        ELSIF x = 5780 THEN
            sigmoid_f := 1932;
        ELSIF x = 5781 THEN
            sigmoid_f := 1932;
        ELSIF x = 5782 THEN
            sigmoid_f := 1932;
        ELSIF x = 5783 THEN
            sigmoid_f := 1933;
        ELSIF x = 5784 THEN
            sigmoid_f := 1933;
        ELSIF x = 5785 THEN
            sigmoid_f := 1933;
        ELSIF x = 5786 THEN
            sigmoid_f := 1933;
        ELSIF x = 5787 THEN
            sigmoid_f := 1933;
        ELSIF x = 5788 THEN
            sigmoid_f := 1933;
        ELSIF x = 5789 THEN
            sigmoid_f := 1933;
        ELSIF x = 5790 THEN
            sigmoid_f := 1933;
        ELSIF x = 5791 THEN
            sigmoid_f := 1933;
        ELSIF x = 5792 THEN
            sigmoid_f := 1933;
        ELSIF x = 5793 THEN
            sigmoid_f := 1933;
        ELSIF x = 5794 THEN
            sigmoid_f := 1933;
        ELSIF x = 5795 THEN
            sigmoid_f := 1933;
        ELSIF x = 5796 THEN
            sigmoid_f := 1933;
        ELSIF x = 5797 THEN
            sigmoid_f := 1933;
        ELSIF x = 5798 THEN
            sigmoid_f := 1933;
        ELSIF x = 5799 THEN
            sigmoid_f := 1933;
        ELSIF x = 5800 THEN
            sigmoid_f := 1933;
        ELSIF x = 5801 THEN
            sigmoid_f := 1933;
        ELSIF x = 5802 THEN
            sigmoid_f := 1933;
        ELSIF x = 5803 THEN
            sigmoid_f := 1934;
        ELSIF x = 5804 THEN
            sigmoid_f := 1934;
        ELSIF x = 5805 THEN
            sigmoid_f := 1934;
        ELSIF x = 5806 THEN
            sigmoid_f := 1934;
        ELSIF x = 5807 THEN
            sigmoid_f := 1934;
        ELSIF x = 5808 THEN
            sigmoid_f := 1934;
        ELSIF x = 5809 THEN
            sigmoid_f := 1934;
        ELSIF x = 5810 THEN
            sigmoid_f := 1934;
        ELSIF x = 5811 THEN
            sigmoid_f := 1934;
        ELSIF x = 5812 THEN
            sigmoid_f := 1934;
        ELSIF x = 5813 THEN
            sigmoid_f := 1934;
        ELSIF x = 5814 THEN
            sigmoid_f := 1934;
        ELSIF x = 5815 THEN
            sigmoid_f := 1934;
        ELSIF x = 5816 THEN
            sigmoid_f := 1934;
        ELSIF x = 5817 THEN
            sigmoid_f := 1934;
        ELSIF x = 5818 THEN
            sigmoid_f := 1934;
        ELSIF x = 5819 THEN
            sigmoid_f := 1934;
        ELSIF x = 5820 THEN
            sigmoid_f := 1934;
        ELSIF x = 5821 THEN
            sigmoid_f := 1934;
        ELSIF x = 5822 THEN
            sigmoid_f := 1934;
        ELSIF x = 5823 THEN
            sigmoid_f := 1935;
        ELSIF x = 5824 THEN
            sigmoid_f := 1935;
        ELSIF x = 5825 THEN
            sigmoid_f := 1935;
        ELSIF x = 5826 THEN
            sigmoid_f := 1935;
        ELSIF x = 5827 THEN
            sigmoid_f := 1935;
        ELSIF x = 5828 THEN
            sigmoid_f := 1935;
        ELSIF x = 5829 THEN
            sigmoid_f := 1935;
        ELSIF x = 5830 THEN
            sigmoid_f := 1935;
        ELSIF x = 5831 THEN
            sigmoid_f := 1935;
        ELSIF x = 5832 THEN
            sigmoid_f := 1935;
        ELSIF x = 5833 THEN
            sigmoid_f := 1935;
        ELSIF x = 5834 THEN
            sigmoid_f := 1935;
        ELSIF x = 5835 THEN
            sigmoid_f := 1935;
        ELSIF x = 5836 THEN
            sigmoid_f := 1935;
        ELSIF x = 5837 THEN
            sigmoid_f := 1935;
        ELSIF x = 5838 THEN
            sigmoid_f := 1935;
        ELSIF x = 5839 THEN
            sigmoid_f := 1935;
        ELSIF x = 5840 THEN
            sigmoid_f := 1935;
        ELSIF x = 5841 THEN
            sigmoid_f := 1935;
        ELSIF x = 5842 THEN
            sigmoid_f := 1935;
        ELSIF x = 5843 THEN
            sigmoid_f := 1936;
        ELSIF x = 5844 THEN
            sigmoid_f := 1936;
        ELSIF x = 5845 THEN
            sigmoid_f := 1936;
        ELSIF x = 5846 THEN
            sigmoid_f := 1936;
        ELSIF x = 5847 THEN
            sigmoid_f := 1936;
        ELSIF x = 5848 THEN
            sigmoid_f := 1936;
        ELSIF x = 5849 THEN
            sigmoid_f := 1936;
        ELSIF x = 5850 THEN
            sigmoid_f := 1936;
        ELSIF x = 5851 THEN
            sigmoid_f := 1936;
        ELSIF x = 5852 THEN
            sigmoid_f := 1936;
        ELSIF x = 5853 THEN
            sigmoid_f := 1936;
        ELSIF x = 5854 THEN
            sigmoid_f := 1936;
        ELSIF x = 5855 THEN
            sigmoid_f := 1936;
        ELSIF x = 5856 THEN
            sigmoid_f := 1936;
        ELSIF x = 5857 THEN
            sigmoid_f := 1936;
        ELSIF x = 5858 THEN
            sigmoid_f := 1936;
        ELSIF x = 5859 THEN
            sigmoid_f := 1936;
        ELSIF x = 5860 THEN
            sigmoid_f := 1936;
        ELSIF x = 5861 THEN
            sigmoid_f := 1936;
        ELSIF x = 5862 THEN
            sigmoid_f := 1936;
        ELSIF x = 5863 THEN
            sigmoid_f := 1937;
        ELSIF x = 5864 THEN
            sigmoid_f := 1937;
        ELSIF x = 5865 THEN
            sigmoid_f := 1937;
        ELSIF x = 5866 THEN
            sigmoid_f := 1937;
        ELSIF x = 5867 THEN
            sigmoid_f := 1937;
        ELSIF x = 5868 THEN
            sigmoid_f := 1937;
        ELSIF x = 5869 THEN
            sigmoid_f := 1937;
        ELSIF x = 5870 THEN
            sigmoid_f := 1937;
        ELSIF x = 5871 THEN
            sigmoid_f := 1937;
        ELSIF x = 5872 THEN
            sigmoid_f := 1937;
        ELSIF x = 5873 THEN
            sigmoid_f := 1937;
        ELSIF x = 5874 THEN
            sigmoid_f := 1937;
        ELSIF x = 5875 THEN
            sigmoid_f := 1937;
        ELSIF x = 5876 THEN
            sigmoid_f := 1937;
        ELSIF x = 5877 THEN
            sigmoid_f := 1937;
        ELSIF x = 5878 THEN
            sigmoid_f := 1937;
        ELSIF x = 5879 THEN
            sigmoid_f := 1937;
        ELSIF x = 5880 THEN
            sigmoid_f := 1937;
        ELSIF x = 5881 THEN
            sigmoid_f := 1937;
        ELSIF x = 5882 THEN
            sigmoid_f := 1937;
        ELSIF x = 5883 THEN
            sigmoid_f := 1938;
        ELSIF x = 5884 THEN
            sigmoid_f := 1938;
        ELSIF x = 5885 THEN
            sigmoid_f := 1938;
        ELSIF x = 5886 THEN
            sigmoid_f := 1938;
        ELSIF x = 5887 THEN
            sigmoid_f := 1938;
        ELSIF x = 5888 THEN
            sigmoid_f := 1938;
        ELSIF x = 5889 THEN
            sigmoid_f := 1938;
        ELSIF x = 5890 THEN
            sigmoid_f := 1938;
        ELSIF x = 5891 THEN
            sigmoid_f := 1938;
        ELSIF x = 5892 THEN
            sigmoid_f := 1938;
        ELSIF x = 5893 THEN
            sigmoid_f := 1938;
        ELSIF x = 5894 THEN
            sigmoid_f := 1938;
        ELSIF x = 5895 THEN
            sigmoid_f := 1938;
        ELSIF x = 5896 THEN
            sigmoid_f := 1938;
        ELSIF x = 5897 THEN
            sigmoid_f := 1938;
        ELSIF x = 5898 THEN
            sigmoid_f := 1938;
        ELSIF x = 5899 THEN
            sigmoid_f := 1938;
        ELSIF x = 5900 THEN
            sigmoid_f := 1938;
        ELSIF x = 5901 THEN
            sigmoid_f := 1938;
        ELSIF x = 5902 THEN
            sigmoid_f := 1938;
        ELSIF x = 5903 THEN
            sigmoid_f := 1938;
        ELSIF x = 5904 THEN
            sigmoid_f := 1939;
        ELSIF x = 5905 THEN
            sigmoid_f := 1939;
        ELSIF x = 5906 THEN
            sigmoid_f := 1939;
        ELSIF x = 5907 THEN
            sigmoid_f := 1939;
        ELSIF x = 5908 THEN
            sigmoid_f := 1939;
        ELSIF x = 5909 THEN
            sigmoid_f := 1939;
        ELSIF x = 5910 THEN
            sigmoid_f := 1939;
        ELSIF x = 5911 THEN
            sigmoid_f := 1939;
        ELSIF x = 5912 THEN
            sigmoid_f := 1939;
        ELSIF x = 5913 THEN
            sigmoid_f := 1939;
        ELSIF x = 5914 THEN
            sigmoid_f := 1939;
        ELSIF x = 5915 THEN
            sigmoid_f := 1939;
        ELSIF x = 5916 THEN
            sigmoid_f := 1939;
        ELSIF x = 5917 THEN
            sigmoid_f := 1939;
        ELSIF x = 5918 THEN
            sigmoid_f := 1939;
        ELSIF x = 5919 THEN
            sigmoid_f := 1939;
        ELSIF x = 5920 THEN
            sigmoid_f := 1939;
        ELSIF x = 5921 THEN
            sigmoid_f := 1939;
        ELSIF x = 5922 THEN
            sigmoid_f := 1939;
        ELSIF x = 5923 THEN
            sigmoid_f := 1939;
        ELSIF x = 5924 THEN
            sigmoid_f := 1940;
        ELSIF x = 5925 THEN
            sigmoid_f := 1940;
        ELSIF x = 5926 THEN
            sigmoid_f := 1940;
        ELSIF x = 5927 THEN
            sigmoid_f := 1940;
        ELSIF x = 5928 THEN
            sigmoid_f := 1940;
        ELSIF x = 5929 THEN
            sigmoid_f := 1940;
        ELSIF x = 5930 THEN
            sigmoid_f := 1940;
        ELSIF x = 5931 THEN
            sigmoid_f := 1940;
        ELSIF x = 5932 THEN
            sigmoid_f := 1940;
        ELSIF x = 5933 THEN
            sigmoid_f := 1940;
        ELSIF x = 5934 THEN
            sigmoid_f := 1940;
        ELSIF x = 5935 THEN
            sigmoid_f := 1940;
        ELSIF x = 5936 THEN
            sigmoid_f := 1940;
        ELSIF x = 5937 THEN
            sigmoid_f := 1940;
        ELSIF x = 5938 THEN
            sigmoid_f := 1940;
        ELSIF x = 5939 THEN
            sigmoid_f := 1940;
        ELSIF x = 5940 THEN
            sigmoid_f := 1940;
        ELSIF x = 5941 THEN
            sigmoid_f := 1940;
        ELSIF x = 5942 THEN
            sigmoid_f := 1940;
        ELSIF x = 5943 THEN
            sigmoid_f := 1940;
        ELSIF x = 5944 THEN
            sigmoid_f := 1941;
        ELSIF x = 5945 THEN
            sigmoid_f := 1941;
        ELSIF x = 5946 THEN
            sigmoid_f := 1941;
        ELSIF x = 5947 THEN
            sigmoid_f := 1941;
        ELSIF x = 5948 THEN
            sigmoid_f := 1941;
        ELSIF x = 5949 THEN
            sigmoid_f := 1941;
        ELSIF x = 5950 THEN
            sigmoid_f := 1941;
        ELSIF x = 5951 THEN
            sigmoid_f := 1941;
        ELSIF x = 5952 THEN
            sigmoid_f := 1941;
        ELSIF x = 5953 THEN
            sigmoid_f := 1941;
        ELSIF x = 5954 THEN
            sigmoid_f := 1941;
        ELSIF x = 5955 THEN
            sigmoid_f := 1941;
        ELSIF x = 5956 THEN
            sigmoid_f := 1941;
        ELSIF x = 5957 THEN
            sigmoid_f := 1941;
        ELSIF x = 5958 THEN
            sigmoid_f := 1941;
        ELSIF x = 5959 THEN
            sigmoid_f := 1941;
        ELSIF x = 5960 THEN
            sigmoid_f := 1941;
        ELSIF x = 5961 THEN
            sigmoid_f := 1941;
        ELSIF x = 5962 THEN
            sigmoid_f := 1941;
        ELSIF x = 5963 THEN
            sigmoid_f := 1941;
        ELSIF x = 5964 THEN
            sigmoid_f := 1942;
        ELSIF x = 5965 THEN
            sigmoid_f := 1942;
        ELSIF x = 5966 THEN
            sigmoid_f := 1942;
        ELSIF x = 5967 THEN
            sigmoid_f := 1942;
        ELSIF x = 5968 THEN
            sigmoid_f := 1942;
        ELSIF x = 5969 THEN
            sigmoid_f := 1942;
        ELSIF x = 5970 THEN
            sigmoid_f := 1942;
        ELSIF x = 5971 THEN
            sigmoid_f := 1942;
        ELSIF x = 5972 THEN
            sigmoid_f := 1942;
        ELSIF x = 5973 THEN
            sigmoid_f := 1942;
        ELSIF x = 5974 THEN
            sigmoid_f := 1942;
        ELSIF x = 5975 THEN
            sigmoid_f := 1942;
        ELSIF x = 5976 THEN
            sigmoid_f := 1942;
        ELSIF x = 5977 THEN
            sigmoid_f := 1942;
        ELSIF x = 5978 THEN
            sigmoid_f := 1942;
        ELSIF x = 5979 THEN
            sigmoid_f := 1942;
        ELSIF x = 5980 THEN
            sigmoid_f := 1942;
        ELSIF x = 5981 THEN
            sigmoid_f := 1942;
        ELSIF x = 5982 THEN
            sigmoid_f := 1942;
        ELSIF x = 5983 THEN
            sigmoid_f := 1942;
        ELSIF x = 5984 THEN
            sigmoid_f := 1943;
        ELSIF x = 5985 THEN
            sigmoid_f := 1943;
        ELSIF x = 5986 THEN
            sigmoid_f := 1943;
        ELSIF x = 5987 THEN
            sigmoid_f := 1943;
        ELSIF x = 5988 THEN
            sigmoid_f := 1943;
        ELSIF x = 5989 THEN
            sigmoid_f := 1943;
        ELSIF x = 5990 THEN
            sigmoid_f := 1943;
        ELSIF x = 5991 THEN
            sigmoid_f := 1943;
        ELSIF x = 5992 THEN
            sigmoid_f := 1943;
        ELSIF x = 5993 THEN
            sigmoid_f := 1943;
        ELSIF x = 5994 THEN
            sigmoid_f := 1943;
        ELSIF x = 5995 THEN
            sigmoid_f := 1943;
        ELSIF x = 5996 THEN
            sigmoid_f := 1943;
        ELSIF x = 5997 THEN
            sigmoid_f := 1943;
        ELSIF x = 5998 THEN
            sigmoid_f := 1943;
        ELSIF x = 5999 THEN
            sigmoid_f := 1943;
        ELSIF x = 6000 THEN
            sigmoid_f := 1943;
        ELSIF x = 6001 THEN
            sigmoid_f := 1943;
        ELSIF x = 6002 THEN
            sigmoid_f := 1943;
        ELSIF x = 6003 THEN
            sigmoid_f := 1943;
        ELSIF x = 6004 THEN
            sigmoid_f := 1944;
        ELSIF x = 6005 THEN
            sigmoid_f := 1944;
        ELSIF x = 6006 THEN
            sigmoid_f := 1944;
        ELSIF x = 6007 THEN
            sigmoid_f := 1944;
        ELSIF x = 6008 THEN
            sigmoid_f := 1944;
        ELSIF x = 6009 THEN
            sigmoid_f := 1944;
        ELSIF x = 6010 THEN
            sigmoid_f := 1944;
        ELSIF x = 6011 THEN
            sigmoid_f := 1944;
        ELSIF x = 6012 THEN
            sigmoid_f := 1944;
        ELSIF x = 6013 THEN
            sigmoid_f := 1944;
        ELSIF x = 6014 THEN
            sigmoid_f := 1944;
        ELSIF x = 6015 THEN
            sigmoid_f := 1944;
        ELSIF x = 6016 THEN
            sigmoid_f := 1944;
        ELSIF x = 6017 THEN
            sigmoid_f := 1944;
        ELSIF x = 6018 THEN
            sigmoid_f := 1944;
        ELSIF x = 6019 THEN
            sigmoid_f := 1944;
        ELSIF x = 6020 THEN
            sigmoid_f := 1944;
        ELSIF x = 6021 THEN
            sigmoid_f := 1944;
        ELSIF x = 6022 THEN
            sigmoid_f := 1944;
        ELSIF x = 6023 THEN
            sigmoid_f := 1944;
        ELSIF x = 6024 THEN
            sigmoid_f := 1945;
        ELSIF x = 6025 THEN
            sigmoid_f := 1945;
        ELSIF x = 6026 THEN
            sigmoid_f := 1945;
        ELSIF x = 6027 THEN
            sigmoid_f := 1945;
        ELSIF x = 6028 THEN
            sigmoid_f := 1945;
        ELSIF x = 6029 THEN
            sigmoid_f := 1945;
        ELSIF x = 6030 THEN
            sigmoid_f := 1945;
        ELSIF x = 6031 THEN
            sigmoid_f := 1945;
        ELSIF x = 6032 THEN
            sigmoid_f := 1945;
        ELSIF x = 6033 THEN
            sigmoid_f := 1945;
        ELSIF x = 6034 THEN
            sigmoid_f := 1945;
        ELSIF x = 6035 THEN
            sigmoid_f := 1945;
        ELSIF x = 6036 THEN
            sigmoid_f := 1945;
        ELSIF x = 6037 THEN
            sigmoid_f := 1945;
        ELSIF x = 6038 THEN
            sigmoid_f := 1945;
        ELSIF x = 6039 THEN
            sigmoid_f := 1945;
        ELSIF x = 6040 THEN
            sigmoid_f := 1945;
        ELSIF x = 6041 THEN
            sigmoid_f := 1945;
        ELSIF x = 6042 THEN
            sigmoid_f := 1945;
        ELSIF x = 6043 THEN
            sigmoid_f := 1945;
        ELSIF x = 6044 THEN
            sigmoid_f := 1946;
        ELSIF x = 6045 THEN
            sigmoid_f := 1946;
        ELSIF x = 6046 THEN
            sigmoid_f := 1946;
        ELSIF x = 6047 THEN
            sigmoid_f := 1946;
        ELSIF x = 6048 THEN
            sigmoid_f := 1946;
        ELSIF x = 6049 THEN
            sigmoid_f := 1946;
        ELSIF x = 6050 THEN
            sigmoid_f := 1946;
        ELSIF x = 6051 THEN
            sigmoid_f := 1946;
        ELSIF x = 6052 THEN
            sigmoid_f := 1946;
        ELSIF x = 6053 THEN
            sigmoid_f := 1946;
        ELSIF x = 6054 THEN
            sigmoid_f := 1946;
        ELSIF x = 6055 THEN
            sigmoid_f := 1946;
        ELSIF x = 6056 THEN
            sigmoid_f := 1946;
        ELSIF x = 6057 THEN
            sigmoid_f := 1946;
        ELSIF x = 6058 THEN
            sigmoid_f := 1946;
        ELSIF x = 6059 THEN
            sigmoid_f := 1946;
        ELSIF x = 6060 THEN
            sigmoid_f := 1946;
        ELSIF x = 6061 THEN
            sigmoid_f := 1946;
        ELSIF x = 6062 THEN
            sigmoid_f := 1946;
        ELSIF x = 6063 THEN
            sigmoid_f := 1946;
        ELSIF x = 6064 THEN
            sigmoid_f := 1947;
        ELSIF x = 6065 THEN
            sigmoid_f := 1947;
        ELSIF x = 6066 THEN
            sigmoid_f := 1947;
        ELSIF x = 6067 THEN
            sigmoid_f := 1947;
        ELSIF x = 6068 THEN
            sigmoid_f := 1947;
        ELSIF x = 6069 THEN
            sigmoid_f := 1947;
        ELSIF x = 6070 THEN
            sigmoid_f := 1947;
        ELSIF x = 6071 THEN
            sigmoid_f := 1947;
        ELSIF x = 6072 THEN
            sigmoid_f := 1947;
        ELSIF x = 6073 THEN
            sigmoid_f := 1947;
        ELSIF x = 6074 THEN
            sigmoid_f := 1947;
        ELSIF x = 6075 THEN
            sigmoid_f := 1947;
        ELSIF x = 6076 THEN
            sigmoid_f := 1947;
        ELSIF x = 6077 THEN
            sigmoid_f := 1947;
        ELSIF x = 6078 THEN
            sigmoid_f := 1947;
        ELSIF x = 6079 THEN
            sigmoid_f := 1947;
        ELSIF x = 6080 THEN
            sigmoid_f := 1947;
        ELSIF x = 6081 THEN
            sigmoid_f := 1947;
        ELSIF x = 6082 THEN
            sigmoid_f := 1947;
        ELSIF x = 6083 THEN
            sigmoid_f := 1947;
        ELSIF x = 6084 THEN
            sigmoid_f := 1948;
        ELSIF x = 6085 THEN
            sigmoid_f := 1948;
        ELSIF x = 6086 THEN
            sigmoid_f := 1948;
        ELSIF x = 6087 THEN
            sigmoid_f := 1948;
        ELSIF x = 6088 THEN
            sigmoid_f := 1948;
        ELSIF x = 6089 THEN
            sigmoid_f := 1948;
        ELSIF x = 6090 THEN
            sigmoid_f := 1948;
        ELSIF x = 6091 THEN
            sigmoid_f := 1948;
        ELSIF x = 6092 THEN
            sigmoid_f := 1948;
        ELSIF x = 6093 THEN
            sigmoid_f := 1948;
        ELSIF x = 6094 THEN
            sigmoid_f := 1948;
        ELSIF x = 6095 THEN
            sigmoid_f := 1948;
        ELSIF x = 6096 THEN
            sigmoid_f := 1948;
        ELSIF x = 6097 THEN
            sigmoid_f := 1948;
        ELSIF x = 6098 THEN
            sigmoid_f := 1948;
        ELSIF x = 6099 THEN
            sigmoid_f := 1948;
        ELSIF x = 6100 THEN
            sigmoid_f := 1948;
        ELSIF x = 6101 THEN
            sigmoid_f := 1948;
        ELSIF x = 6102 THEN
            sigmoid_f := 1948;
        ELSIF x = 6103 THEN
            sigmoid_f := 1948;
        ELSIF x = 6104 THEN
            sigmoid_f := 1949;
        ELSIF x = 6105 THEN
            sigmoid_f := 1949;
        ELSIF x = 6106 THEN
            sigmoid_f := 1949;
        ELSIF x = 6107 THEN
            sigmoid_f := 1949;
        ELSIF x = 6108 THEN
            sigmoid_f := 1949;
        ELSIF x = 6109 THEN
            sigmoid_f := 1949;
        ELSIF x = 6110 THEN
            sigmoid_f := 1949;
        ELSIF x = 6111 THEN
            sigmoid_f := 1949;
        ELSIF x = 6112 THEN
            sigmoid_f := 1949;
        ELSIF x = 6113 THEN
            sigmoid_f := 1949;
        ELSIF x = 6114 THEN
            sigmoid_f := 1949;
        ELSIF x = 6115 THEN
            sigmoid_f := 1949;
        ELSIF x = 6116 THEN
            sigmoid_f := 1949;
        ELSIF x = 6117 THEN
            sigmoid_f := 1949;
        ELSIF x = 6118 THEN
            sigmoid_f := 1949;
        ELSIF x = 6119 THEN
            sigmoid_f := 1949;
        ELSIF x = 6120 THEN
            sigmoid_f := 1949;
        ELSIF x = 6121 THEN
            sigmoid_f := 1949;
        ELSIF x = 6122 THEN
            sigmoid_f := 1949;
        ELSIF x = 6123 THEN
            sigmoid_f := 1949;
        ELSIF x = 6124 THEN
            sigmoid_f := 1950;
        ELSIF x = 6125 THEN
            sigmoid_f := 1950;
        ELSIF x = 6126 THEN
            sigmoid_f := 1950;
        ELSIF x = 6127 THEN
            sigmoid_f := 1950;
        ELSIF x = 6128 THEN
            sigmoid_f := 1950;
        ELSIF x = 6129 THEN
            sigmoid_f := 1950;
        ELSIF x = 6130 THEN
            sigmoid_f := 1950;
        ELSIF x = 6131 THEN
            sigmoid_f := 1950;
        ELSIF x = 6132 THEN
            sigmoid_f := 1950;
        ELSIF x = 6133 THEN
            sigmoid_f := 1950;
        ELSIF x = 6134 THEN
            sigmoid_f := 1950;
        ELSIF x = 6135 THEN
            sigmoid_f := 1950;
        ELSIF x = 6136 THEN
            sigmoid_f := 1950;
        ELSIF x = 6137 THEN
            sigmoid_f := 1950;
        ELSIF x = 6138 THEN
            sigmoid_f := 1950;
        ELSIF x = 6139 THEN
            sigmoid_f := 1950;
        ELSIF x = 6140 THEN
            sigmoid_f := 1950;
        ELSIF x = 6141 THEN
            sigmoid_f := 1950;
        ELSIF x = 6142 THEN
            sigmoid_f := 1950;
        ELSIF x = 6143 THEN
            sigmoid_f := 1950;
        ELSIF x = 6144 THEN
            sigmoid_f := 1951;
        ELSIF x = 6145 THEN
            sigmoid_f := 1951;
        ELSIF x = 6146 THEN
            sigmoid_f := 1951;
        ELSIF x = 6147 THEN
            sigmoid_f := 1951;
        ELSIF x = 6148 THEN
            sigmoid_f := 1951;
        ELSIF x = 6149 THEN
            sigmoid_f := 1951;
        ELSIF x = 6150 THEN
            sigmoid_f := 1951;
        ELSIF x = 6151 THEN
            sigmoid_f := 1951;
        ELSIF x = 6152 THEN
            sigmoid_f := 1951;
        ELSIF x = 6153 THEN
            sigmoid_f := 1951;
        ELSIF x = 6154 THEN
            sigmoid_f := 1951;
        ELSIF x = 6155 THEN
            sigmoid_f := 1951;
        ELSIF x = 6156 THEN
            sigmoid_f := 1951;
        ELSIF x = 6157 THEN
            sigmoid_f := 1951;
        ELSIF x = 6158 THEN
            sigmoid_f := 1951;
        ELSIF x = 6159 THEN
            sigmoid_f := 1951;
        ELSIF x = 6160 THEN
            sigmoid_f := 1951;
        ELSIF x = 6161 THEN
            sigmoid_f := 1951;
        ELSIF x = 6162 THEN
            sigmoid_f := 1951;
        ELSIF x = 6163 THEN
            sigmoid_f := 1951;
        ELSIF x = 6164 THEN
            sigmoid_f := 1951;
        ELSIF x = 6165 THEN
            sigmoid_f := 1951;
        ELSIF x = 6166 THEN
            sigmoid_f := 1951;
        ELSIF x = 6167 THEN
            sigmoid_f := 1951;
        ELSIF x = 6168 THEN
            sigmoid_f := 1951;
        ELSIF x = 6169 THEN
            sigmoid_f := 1952;
        ELSIF x = 6170 THEN
            sigmoid_f := 1952;
        ELSIF x = 6171 THEN
            sigmoid_f := 1952;
        ELSIF x = 6172 THEN
            sigmoid_f := 1952;
        ELSIF x = 6173 THEN
            sigmoid_f := 1952;
        ELSIF x = 6174 THEN
            sigmoid_f := 1952;
        ELSIF x = 6175 THEN
            sigmoid_f := 1952;
        ELSIF x = 6176 THEN
            sigmoid_f := 1952;
        ELSIF x = 6177 THEN
            sigmoid_f := 1952;
        ELSIF x = 6178 THEN
            sigmoid_f := 1952;
        ELSIF x = 6179 THEN
            sigmoid_f := 1952;
        ELSIF x = 6180 THEN
            sigmoid_f := 1952;
        ELSIF x = 6181 THEN
            sigmoid_f := 1952;
        ELSIF x = 6182 THEN
            sigmoid_f := 1952;
        ELSIF x = 6183 THEN
            sigmoid_f := 1952;
        ELSIF x = 6184 THEN
            sigmoid_f := 1952;
        ELSIF x = 6185 THEN
            sigmoid_f := 1952;
        ELSIF x = 6186 THEN
            sigmoid_f := 1952;
        ELSIF x = 6187 THEN
            sigmoid_f := 1952;
        ELSIF x = 6188 THEN
            sigmoid_f := 1952;
        ELSIF x = 6189 THEN
            sigmoid_f := 1952;
        ELSIF x = 6190 THEN
            sigmoid_f := 1952;
        ELSIF x = 6191 THEN
            sigmoid_f := 1952;
        ELSIF x = 6192 THEN
            sigmoid_f := 1952;
        ELSIF x = 6193 THEN
            sigmoid_f := 1953;
        ELSIF x = 6194 THEN
            sigmoid_f := 1953;
        ELSIF x = 6195 THEN
            sigmoid_f := 1953;
        ELSIF x = 6196 THEN
            sigmoid_f := 1953;
        ELSIF x = 6197 THEN
            sigmoid_f := 1953;
        ELSIF x = 6198 THEN
            sigmoid_f := 1953;
        ELSIF x = 6199 THEN
            sigmoid_f := 1953;
        ELSIF x = 6200 THEN
            sigmoid_f := 1953;
        ELSIF x = 6201 THEN
            sigmoid_f := 1953;
        ELSIF x = 6202 THEN
            sigmoid_f := 1953;
        ELSIF x = 6203 THEN
            sigmoid_f := 1953;
        ELSIF x = 6204 THEN
            sigmoid_f := 1953;
        ELSIF x = 6205 THEN
            sigmoid_f := 1953;
        ELSIF x = 6206 THEN
            sigmoid_f := 1953;
        ELSIF x = 6207 THEN
            sigmoid_f := 1953;
        ELSIF x = 6208 THEN
            sigmoid_f := 1953;
        ELSIF x = 6209 THEN
            sigmoid_f := 1953;
        ELSIF x = 6210 THEN
            sigmoid_f := 1953;
        ELSIF x = 6211 THEN
            sigmoid_f := 1953;
        ELSIF x = 6212 THEN
            sigmoid_f := 1953;
        ELSIF x = 6213 THEN
            sigmoid_f := 1953;
        ELSIF x = 6214 THEN
            sigmoid_f := 1953;
        ELSIF x = 6215 THEN
            sigmoid_f := 1953;
        ELSIF x = 6216 THEN
            sigmoid_f := 1953;
        ELSIF x = 6217 THEN
            sigmoid_f := 1953;
        ELSIF x = 6218 THEN
            sigmoid_f := 1954;
        ELSIF x = 6219 THEN
            sigmoid_f := 1954;
        ELSIF x = 6220 THEN
            sigmoid_f := 1954;
        ELSIF x = 6221 THEN
            sigmoid_f := 1954;
        ELSIF x = 6222 THEN
            sigmoid_f := 1954;
        ELSIF x = 6223 THEN
            sigmoid_f := 1954;
        ELSIF x = 6224 THEN
            sigmoid_f := 1954;
        ELSIF x = 6225 THEN
            sigmoid_f := 1954;
        ELSIF x = 6226 THEN
            sigmoid_f := 1954;
        ELSIF x = 6227 THEN
            sigmoid_f := 1954;
        ELSIF x = 6228 THEN
            sigmoid_f := 1954;
        ELSIF x = 6229 THEN
            sigmoid_f := 1954;
        ELSIF x = 6230 THEN
            sigmoid_f := 1954;
        ELSIF x = 6231 THEN
            sigmoid_f := 1954;
        ELSIF x = 6232 THEN
            sigmoid_f := 1954;
        ELSIF x = 6233 THEN
            sigmoid_f := 1954;
        ELSIF x = 6234 THEN
            sigmoid_f := 1954;
        ELSIF x = 6235 THEN
            sigmoid_f := 1954;
        ELSIF x = 6236 THEN
            sigmoid_f := 1954;
        ELSIF x = 6237 THEN
            sigmoid_f := 1954;
        ELSIF x = 6238 THEN
            sigmoid_f := 1954;
        ELSIF x = 6239 THEN
            sigmoid_f := 1954;
        ELSIF x = 6240 THEN
            sigmoid_f := 1954;
        ELSIF x = 6241 THEN
            sigmoid_f := 1954;
        ELSIF x = 6242 THEN
            sigmoid_f := 1955;
        ELSIF x = 6243 THEN
            sigmoid_f := 1955;
        ELSIF x = 6244 THEN
            sigmoid_f := 1955;
        ELSIF x = 6245 THEN
            sigmoid_f := 1955;
        ELSIF x = 6246 THEN
            sigmoid_f := 1955;
        ELSIF x = 6247 THEN
            sigmoid_f := 1955;
        ELSIF x = 6248 THEN
            sigmoid_f := 1955;
        ELSIF x = 6249 THEN
            sigmoid_f := 1955;
        ELSIF x = 6250 THEN
            sigmoid_f := 1955;
        ELSIF x = 6251 THEN
            sigmoid_f := 1955;
        ELSIF x = 6252 THEN
            sigmoid_f := 1955;
        ELSIF x = 6253 THEN
            sigmoid_f := 1955;
        ELSIF x = 6254 THEN
            sigmoid_f := 1955;
        ELSIF x = 6255 THEN
            sigmoid_f := 1955;
        ELSIF x = 6256 THEN
            sigmoid_f := 1955;
        ELSIF x = 6257 THEN
            sigmoid_f := 1955;
        ELSIF x = 6258 THEN
            sigmoid_f := 1955;
        ELSIF x = 6259 THEN
            sigmoid_f := 1955;
        ELSIF x = 6260 THEN
            sigmoid_f := 1955;
        ELSIF x = 6261 THEN
            sigmoid_f := 1955;
        ELSIF x = 6262 THEN
            sigmoid_f := 1955;
        ELSIF x = 6263 THEN
            sigmoid_f := 1955;
        ELSIF x = 6264 THEN
            sigmoid_f := 1955;
        ELSIF x = 6265 THEN
            sigmoid_f := 1955;
        ELSIF x = 6266 THEN
            sigmoid_f := 1956;
        ELSIF x = 6267 THEN
            sigmoid_f := 1956;
        ELSIF x = 6268 THEN
            sigmoid_f := 1956;
        ELSIF x = 6269 THEN
            sigmoid_f := 1956;
        ELSIF x = 6270 THEN
            sigmoid_f := 1956;
        ELSIF x = 6271 THEN
            sigmoid_f := 1956;
        ELSIF x = 6272 THEN
            sigmoid_f := 1956;
        ELSIF x = 6273 THEN
            sigmoid_f := 1956;
        ELSIF x = 6274 THEN
            sigmoid_f := 1956;
        ELSIF x = 6275 THEN
            sigmoid_f := 1956;
        ELSIF x = 6276 THEN
            sigmoid_f := 1956;
        ELSIF x = 6277 THEN
            sigmoid_f := 1956;
        ELSIF x = 6278 THEN
            sigmoid_f := 1956;
        ELSIF x = 6279 THEN
            sigmoid_f := 1956;
        ELSIF x = 6280 THEN
            sigmoid_f := 1956;
        ELSIF x = 6281 THEN
            sigmoid_f := 1956;
        ELSIF x = 6282 THEN
            sigmoid_f := 1956;
        ELSIF x = 6283 THEN
            sigmoid_f := 1956;
        ELSIF x = 6284 THEN
            sigmoid_f := 1956;
        ELSIF x = 6285 THEN
            sigmoid_f := 1956;
        ELSIF x = 6286 THEN
            sigmoid_f := 1956;
        ELSIF x = 6287 THEN
            sigmoid_f := 1956;
        ELSIF x = 6288 THEN
            sigmoid_f := 1956;
        ELSIF x = 6289 THEN
            sigmoid_f := 1956;
        ELSIF x = 6290 THEN
            sigmoid_f := 1956;
        ELSIF x = 6291 THEN
            sigmoid_f := 1957;
        ELSIF x = 6292 THEN
            sigmoid_f := 1957;
        ELSIF x = 6293 THEN
            sigmoid_f := 1957;
        ELSIF x = 6294 THEN
            sigmoid_f := 1957;
        ELSIF x = 6295 THEN
            sigmoid_f := 1957;
        ELSIF x = 6296 THEN
            sigmoid_f := 1957;
        ELSIF x = 6297 THEN
            sigmoid_f := 1957;
        ELSIF x = 6298 THEN
            sigmoid_f := 1957;
        ELSIF x = 6299 THEN
            sigmoid_f := 1957;
        ELSIF x = 6300 THEN
            sigmoid_f := 1957;
        ELSIF x = 6301 THEN
            sigmoid_f := 1957;
        ELSIF x = 6302 THEN
            sigmoid_f := 1957;
        ELSIF x = 6303 THEN
            sigmoid_f := 1957;
        ELSIF x = 6304 THEN
            sigmoid_f := 1957;
        ELSIF x = 6305 THEN
            sigmoid_f := 1957;
        ELSIF x = 6306 THEN
            sigmoid_f := 1957;
        ELSIF x = 6307 THEN
            sigmoid_f := 1957;
        ELSIF x = 6308 THEN
            sigmoid_f := 1957;
        ELSIF x = 6309 THEN
            sigmoid_f := 1957;
        ELSIF x = 6310 THEN
            sigmoid_f := 1957;
        ELSIF x = 6311 THEN
            sigmoid_f := 1957;
        ELSIF x = 6312 THEN
            sigmoid_f := 1957;
        ELSIF x = 6313 THEN
            sigmoid_f := 1957;
        ELSIF x = 6314 THEN
            sigmoid_f := 1957;
        ELSIF x = 6315 THEN
            sigmoid_f := 1958;
        ELSIF x = 6316 THEN
            sigmoid_f := 1958;
        ELSIF x = 6317 THEN
            sigmoid_f := 1958;
        ELSIF x = 6318 THEN
            sigmoid_f := 1958;
        ELSIF x = 6319 THEN
            sigmoid_f := 1958;
        ELSIF x = 6320 THEN
            sigmoid_f := 1958;
        ELSIF x = 6321 THEN
            sigmoid_f := 1958;
        ELSIF x = 6322 THEN
            sigmoid_f := 1958;
        ELSIF x = 6323 THEN
            sigmoid_f := 1958;
        ELSIF x = 6324 THEN
            sigmoid_f := 1958;
        ELSIF x = 6325 THEN
            sigmoid_f := 1958;
        ELSIF x = 6326 THEN
            sigmoid_f := 1958;
        ELSIF x = 6327 THEN
            sigmoid_f := 1958;
        ELSIF x = 6328 THEN
            sigmoid_f := 1958;
        ELSIF x = 6329 THEN
            sigmoid_f := 1958;
        ELSIF x = 6330 THEN
            sigmoid_f := 1958;
        ELSIF x = 6331 THEN
            sigmoid_f := 1958;
        ELSIF x = 6332 THEN
            sigmoid_f := 1958;
        ELSIF x = 6333 THEN
            sigmoid_f := 1958;
        ELSIF x = 6334 THEN
            sigmoid_f := 1958;
        ELSIF x = 6335 THEN
            sigmoid_f := 1958;
        ELSIF x = 6336 THEN
            sigmoid_f := 1958;
        ELSIF x = 6337 THEN
            sigmoid_f := 1958;
        ELSIF x = 6338 THEN
            sigmoid_f := 1958;
        ELSIF x = 6339 THEN
            sigmoid_f := 1958;
        ELSIF x = 6340 THEN
            sigmoid_f := 1959;
        ELSIF x = 6341 THEN
            sigmoid_f := 1959;
        ELSIF x = 6342 THEN
            sigmoid_f := 1959;
        ELSIF x = 6343 THEN
            sigmoid_f := 1959;
        ELSIF x = 6344 THEN
            sigmoid_f := 1959;
        ELSIF x = 6345 THEN
            sigmoid_f := 1959;
        ELSIF x = 6346 THEN
            sigmoid_f := 1959;
        ELSIF x = 6347 THEN
            sigmoid_f := 1959;
        ELSIF x = 6348 THEN
            sigmoid_f := 1959;
        ELSIF x = 6349 THEN
            sigmoid_f := 1959;
        ELSIF x = 6350 THEN
            sigmoid_f := 1959;
        ELSIF x = 6351 THEN
            sigmoid_f := 1959;
        ELSIF x = 6352 THEN
            sigmoid_f := 1959;
        ELSIF x = 6353 THEN
            sigmoid_f := 1959;
        ELSIF x = 6354 THEN
            sigmoid_f := 1959;
        ELSIF x = 6355 THEN
            sigmoid_f := 1959;
        ELSIF x = 6356 THEN
            sigmoid_f := 1959;
        ELSIF x = 6357 THEN
            sigmoid_f := 1959;
        ELSIF x = 6358 THEN
            sigmoid_f := 1959;
        ELSIF x = 6359 THEN
            sigmoid_f := 1959;
        ELSIF x = 6360 THEN
            sigmoid_f := 1959;
        ELSIF x = 6361 THEN
            sigmoid_f := 1959;
        ELSIF x = 6362 THEN
            sigmoid_f := 1959;
        ELSIF x = 6363 THEN
            sigmoid_f := 1959;
        ELSIF x = 6364 THEN
            sigmoid_f := 1960;
        ELSIF x = 6365 THEN
            sigmoid_f := 1960;
        ELSIF x = 6366 THEN
            sigmoid_f := 1960;
        ELSIF x = 6367 THEN
            sigmoid_f := 1960;
        ELSIF x = 6368 THEN
            sigmoid_f := 1960;
        ELSIF x = 6369 THEN
            sigmoid_f := 1960;
        ELSIF x = 6370 THEN
            sigmoid_f := 1960;
        ELSIF x = 6371 THEN
            sigmoid_f := 1960;
        ELSIF x = 6372 THEN
            sigmoid_f := 1960;
        ELSIF x = 6373 THEN
            sigmoid_f := 1960;
        ELSIF x = 6374 THEN
            sigmoid_f := 1960;
        ELSIF x = 6375 THEN
            sigmoid_f := 1960;
        ELSIF x = 6376 THEN
            sigmoid_f := 1960;
        ELSIF x = 6377 THEN
            sigmoid_f := 1960;
        ELSIF x = 6378 THEN
            sigmoid_f := 1960;
        ELSIF x = 6379 THEN
            sigmoid_f := 1960;
        ELSIF x = 6380 THEN
            sigmoid_f := 1960;
        ELSIF x = 6381 THEN
            sigmoid_f := 1960;
        ELSIF x = 6382 THEN
            sigmoid_f := 1960;
        ELSIF x = 6383 THEN
            sigmoid_f := 1960;
        ELSIF x = 6384 THEN
            sigmoid_f := 1960;
        ELSIF x = 6385 THEN
            sigmoid_f := 1960;
        ELSIF x = 6386 THEN
            sigmoid_f := 1960;
        ELSIF x = 6387 THEN
            sigmoid_f := 1960;
        ELSIF x = 6388 THEN
            sigmoid_f := 1961;
        ELSIF x = 6389 THEN
            sigmoid_f := 1961;
        ELSIF x = 6390 THEN
            sigmoid_f := 1961;
        ELSIF x = 6391 THEN
            sigmoid_f := 1961;
        ELSIF x = 6392 THEN
            sigmoid_f := 1961;
        ELSIF x = 6393 THEN
            sigmoid_f := 1961;
        ELSIF x = 6394 THEN
            sigmoid_f := 1961;
        ELSIF x = 6395 THEN
            sigmoid_f := 1961;
        ELSIF x = 6396 THEN
            sigmoid_f := 1961;
        ELSIF x = 6397 THEN
            sigmoid_f := 1961;
        ELSIF x = 6398 THEN
            sigmoid_f := 1961;
        ELSIF x = 6399 THEN
            sigmoid_f := 1961;
        ELSIF x = 6400 THEN
            sigmoid_f := 1961;
        ELSIF x = 6401 THEN
            sigmoid_f := 1961;
        ELSIF x = 6402 THEN
            sigmoid_f := 1961;
        ELSIF x = 6403 THEN
            sigmoid_f := 1961;
        ELSIF x = 6404 THEN
            sigmoid_f := 1961;
        ELSIF x = 6405 THEN
            sigmoid_f := 1961;
        ELSIF x = 6406 THEN
            sigmoid_f := 1961;
        ELSIF x = 6407 THEN
            sigmoid_f := 1961;
        ELSIF x = 6408 THEN
            sigmoid_f := 1961;
        ELSIF x = 6409 THEN
            sigmoid_f := 1961;
        ELSIF x = 6410 THEN
            sigmoid_f := 1961;
        ELSIF x = 6411 THEN
            sigmoid_f := 1961;
        ELSIF x = 6412 THEN
            sigmoid_f := 1961;
        ELSIF x = 6413 THEN
            sigmoid_f := 1962;
        ELSIF x = 6414 THEN
            sigmoid_f := 1962;
        ELSIF x = 6415 THEN
            sigmoid_f := 1962;
        ELSIF x = 6416 THEN
            sigmoid_f := 1962;
        ELSIF x = 6417 THEN
            sigmoid_f := 1962;
        ELSIF x = 6418 THEN
            sigmoid_f := 1962;
        ELSIF x = 6419 THEN
            sigmoid_f := 1962;
        ELSIF x = 6420 THEN
            sigmoid_f := 1962;
        ELSIF x = 6421 THEN
            sigmoid_f := 1962;
        ELSIF x = 6422 THEN
            sigmoid_f := 1962;
        ELSIF x = 6423 THEN
            sigmoid_f := 1962;
        ELSIF x = 6424 THEN
            sigmoid_f := 1962;
        ELSIF x = 6425 THEN
            sigmoid_f := 1962;
        ELSIF x = 6426 THEN
            sigmoid_f := 1962;
        ELSIF x = 6427 THEN
            sigmoid_f := 1962;
        ELSIF x = 6428 THEN
            sigmoid_f := 1962;
        ELSIF x = 6429 THEN
            sigmoid_f := 1962;
        ELSIF x = 6430 THEN
            sigmoid_f := 1962;
        ELSIF x = 6431 THEN
            sigmoid_f := 1962;
        ELSIF x = 6432 THEN
            sigmoid_f := 1962;
        ELSIF x = 6433 THEN
            sigmoid_f := 1962;
        ELSIF x = 6434 THEN
            sigmoid_f := 1962;
        ELSIF x = 6435 THEN
            sigmoid_f := 1962;
        ELSIF x = 6436 THEN
            sigmoid_f := 1962;
        ELSIF x = 6437 THEN
            sigmoid_f := 1963;
        ELSIF x = 6438 THEN
            sigmoid_f := 1963;
        ELSIF x = 6439 THEN
            sigmoid_f := 1963;
        ELSIF x = 6440 THEN
            sigmoid_f := 1963;
        ELSIF x = 6441 THEN
            sigmoid_f := 1963;
        ELSIF x = 6442 THEN
            sigmoid_f := 1963;
        ELSIF x = 6443 THEN
            sigmoid_f := 1963;
        ELSIF x = 6444 THEN
            sigmoid_f := 1963;
        ELSIF x = 6445 THEN
            sigmoid_f := 1963;
        ELSIF x = 6446 THEN
            sigmoid_f := 1963;
        ELSIF x = 6447 THEN
            sigmoid_f := 1963;
        ELSIF x = 6448 THEN
            sigmoid_f := 1963;
        ELSIF x = 6449 THEN
            sigmoid_f := 1963;
        ELSIF x = 6450 THEN
            sigmoid_f := 1963;
        ELSIF x = 6451 THEN
            sigmoid_f := 1963;
        ELSIF x = 6452 THEN
            sigmoid_f := 1963;
        ELSIF x = 6453 THEN
            sigmoid_f := 1963;
        ELSIF x = 6454 THEN
            sigmoid_f := 1963;
        ELSIF x = 6455 THEN
            sigmoid_f := 1963;
        ELSIF x = 6456 THEN
            sigmoid_f := 1963;
        ELSIF x = 6457 THEN
            sigmoid_f := 1963;
        ELSIF x = 6458 THEN
            sigmoid_f := 1963;
        ELSIF x = 6459 THEN
            sigmoid_f := 1963;
        ELSIF x = 6460 THEN
            sigmoid_f := 1963;
        ELSIF x = 6461 THEN
            sigmoid_f := 1964;
        ELSIF x = 6462 THEN
            sigmoid_f := 1964;
        ELSIF x = 6463 THEN
            sigmoid_f := 1964;
        ELSIF x = 6464 THEN
            sigmoid_f := 1964;
        ELSIF x = 6465 THEN
            sigmoid_f := 1964;
        ELSIF x = 6466 THEN
            sigmoid_f := 1964;
        ELSIF x = 6467 THEN
            sigmoid_f := 1964;
        ELSIF x = 6468 THEN
            sigmoid_f := 1964;
        ELSIF x = 6469 THEN
            sigmoid_f := 1964;
        ELSIF x = 6470 THEN
            sigmoid_f := 1964;
        ELSIF x = 6471 THEN
            sigmoid_f := 1964;
        ELSIF x = 6472 THEN
            sigmoid_f := 1964;
        ELSIF x = 6473 THEN
            sigmoid_f := 1964;
        ELSIF x = 6474 THEN
            sigmoid_f := 1964;
        ELSIF x = 6475 THEN
            sigmoid_f := 1964;
        ELSIF x = 6476 THEN
            sigmoid_f := 1964;
        ELSIF x = 6477 THEN
            sigmoid_f := 1964;
        ELSIF x = 6478 THEN
            sigmoid_f := 1964;
        ELSIF x = 6479 THEN
            sigmoid_f := 1964;
        ELSIF x = 6480 THEN
            sigmoid_f := 1964;
        ELSIF x = 6481 THEN
            sigmoid_f := 1964;
        ELSIF x = 6482 THEN
            sigmoid_f := 1964;
        ELSIF x = 6483 THEN
            sigmoid_f := 1964;
        ELSIF x = 6484 THEN
            sigmoid_f := 1964;
        ELSIF x = 6485 THEN
            sigmoid_f := 1964;
        ELSIF x = 6486 THEN
            sigmoid_f := 1965;
        ELSIF x = 6487 THEN
            sigmoid_f := 1965;
        ELSIF x = 6488 THEN
            sigmoid_f := 1965;
        ELSIF x = 6489 THEN
            sigmoid_f := 1965;
        ELSIF x = 6490 THEN
            sigmoid_f := 1965;
        ELSIF x = 6491 THEN
            sigmoid_f := 1965;
        ELSIF x = 6492 THEN
            sigmoid_f := 1965;
        ELSIF x = 6493 THEN
            sigmoid_f := 1965;
        ELSIF x = 6494 THEN
            sigmoid_f := 1965;
        ELSIF x = 6495 THEN
            sigmoid_f := 1965;
        ELSIF x = 6496 THEN
            sigmoid_f := 1965;
        ELSIF x = 6497 THEN
            sigmoid_f := 1965;
        ELSIF x = 6498 THEN
            sigmoid_f := 1965;
        ELSIF x = 6499 THEN
            sigmoid_f := 1965;
        ELSIF x = 6500 THEN
            sigmoid_f := 1965;
        ELSIF x = 6501 THEN
            sigmoid_f := 1965;
        ELSIF x = 6502 THEN
            sigmoid_f := 1965;
        ELSIF x = 6503 THEN
            sigmoid_f := 1965;
        ELSIF x = 6504 THEN
            sigmoid_f := 1965;
        ELSIF x = 6505 THEN
            sigmoid_f := 1965;
        ELSIF x = 6506 THEN
            sigmoid_f := 1965;
        ELSIF x = 6507 THEN
            sigmoid_f := 1965;
        ELSIF x = 6508 THEN
            sigmoid_f := 1965;
        ELSIF x = 6509 THEN
            sigmoid_f := 1965;
        ELSIF x = 6510 THEN
            sigmoid_f := 1966;
        ELSIF x = 6511 THEN
            sigmoid_f := 1966;
        ELSIF x = 6512 THEN
            sigmoid_f := 1966;
        ELSIF x = 6513 THEN
            sigmoid_f := 1966;
        ELSIF x = 6514 THEN
            sigmoid_f := 1966;
        ELSIF x = 6515 THEN
            sigmoid_f := 1966;
        ELSIF x = 6516 THEN
            sigmoid_f := 1966;
        ELSIF x = 6517 THEN
            sigmoid_f := 1966;
        ELSIF x = 6518 THEN
            sigmoid_f := 1966;
        ELSIF x = 6519 THEN
            sigmoid_f := 1966;
        ELSIF x = 6520 THEN
            sigmoid_f := 1966;
        ELSIF x = 6521 THEN
            sigmoid_f := 1966;
        ELSIF x = 6522 THEN
            sigmoid_f := 1966;
        ELSIF x = 6523 THEN
            sigmoid_f := 1966;
        ELSIF x = 6524 THEN
            sigmoid_f := 1966;
        ELSIF x = 6525 THEN
            sigmoid_f := 1966;
        ELSIF x = 6526 THEN
            sigmoid_f := 1966;
        ELSIF x = 6527 THEN
            sigmoid_f := 1966;
        ELSIF x = 6528 THEN
            sigmoid_f := 1966;
        ELSIF x = 6529 THEN
            sigmoid_f := 1966;
        ELSIF x = 6530 THEN
            sigmoid_f := 1966;
        ELSIF x = 6531 THEN
            sigmoid_f := 1966;
        ELSIF x = 6532 THEN
            sigmoid_f := 1966;
        ELSIF x = 6533 THEN
            sigmoid_f := 1966;
        ELSIF x = 6534 THEN
            sigmoid_f := 1966;
        ELSIF x = 6535 THEN
            sigmoid_f := 1967;
        ELSIF x = 6536 THEN
            sigmoid_f := 1967;
        ELSIF x = 6537 THEN
            sigmoid_f := 1967;
        ELSIF x = 6538 THEN
            sigmoid_f := 1967;
        ELSIF x = 6539 THEN
            sigmoid_f := 1967;
        ELSIF x = 6540 THEN
            sigmoid_f := 1967;
        ELSIF x = 6541 THEN
            sigmoid_f := 1967;
        ELSIF x = 6542 THEN
            sigmoid_f := 1967;
        ELSIF x = 6543 THEN
            sigmoid_f := 1967;
        ELSIF x = 6544 THEN
            sigmoid_f := 1967;
        ELSIF x = 6545 THEN
            sigmoid_f := 1967;
        ELSIF x = 6546 THEN
            sigmoid_f := 1967;
        ELSIF x = 6547 THEN
            sigmoid_f := 1967;
        ELSIF x = 6548 THEN
            sigmoid_f := 1967;
        ELSIF x = 6549 THEN
            sigmoid_f := 1967;
        ELSIF x = 6550 THEN
            sigmoid_f := 1967;
        ELSIF x = 6551 THEN
            sigmoid_f := 1967;
        ELSIF x = 6552 THEN
            sigmoid_f := 1967;
        ELSIF x = 6553 THEN
            sigmoid_f := 1967;
        ELSIF x = 6554 THEN
            sigmoid_f := 1967;
        ELSIF x = 6555 THEN
            sigmoid_f := 1967;
        ELSIF x = 6556 THEN
            sigmoid_f := 1967;
        ELSIF x = 6557 THEN
            sigmoid_f := 1967;
        ELSIF x = 6558 THEN
            sigmoid_f := 1967;
        ELSIF x = 6559 THEN
            sigmoid_f := 1968;
        ELSIF x = 6560 THEN
            sigmoid_f := 1968;
        ELSIF x = 6561 THEN
            sigmoid_f := 1968;
        ELSIF x = 6562 THEN
            sigmoid_f := 1968;
        ELSIF x = 6563 THEN
            sigmoid_f := 1968;
        ELSIF x = 6564 THEN
            sigmoid_f := 1968;
        ELSIF x = 6565 THEN
            sigmoid_f := 1968;
        ELSIF x = 6566 THEN
            sigmoid_f := 1968;
        ELSIF x = 6567 THEN
            sigmoid_f := 1968;
        ELSIF x = 6568 THEN
            sigmoid_f := 1968;
        ELSIF x = 6569 THEN
            sigmoid_f := 1968;
        ELSIF x = 6570 THEN
            sigmoid_f := 1968;
        ELSIF x = 6571 THEN
            sigmoid_f := 1968;
        ELSIF x = 6572 THEN
            sigmoid_f := 1968;
        ELSIF x = 6573 THEN
            sigmoid_f := 1968;
        ELSIF x = 6574 THEN
            sigmoid_f := 1968;
        ELSIF x = 6575 THEN
            sigmoid_f := 1968;
        ELSIF x = 6576 THEN
            sigmoid_f := 1968;
        ELSIF x = 6577 THEN
            sigmoid_f := 1968;
        ELSIF x = 6578 THEN
            sigmoid_f := 1968;
        ELSIF x = 6579 THEN
            sigmoid_f := 1968;
        ELSIF x = 6580 THEN
            sigmoid_f := 1968;
        ELSIF x = 6581 THEN
            sigmoid_f := 1968;
        ELSIF x = 6582 THEN
            sigmoid_f := 1968;
        ELSIF x = 6583 THEN
            sigmoid_f := 1969;
        ELSIF x = 6584 THEN
            sigmoid_f := 1969;
        ELSIF x = 6585 THEN
            sigmoid_f := 1969;
        ELSIF x = 6586 THEN
            sigmoid_f := 1969;
        ELSIF x = 6587 THEN
            sigmoid_f := 1969;
        ELSIF x = 6588 THEN
            sigmoid_f := 1969;
        ELSIF x = 6589 THEN
            sigmoid_f := 1969;
        ELSIF x = 6590 THEN
            sigmoid_f := 1969;
        ELSIF x = 6591 THEN
            sigmoid_f := 1969;
        ELSIF x = 6592 THEN
            sigmoid_f := 1969;
        ELSIF x = 6593 THEN
            sigmoid_f := 1969;
        ELSIF x = 6594 THEN
            sigmoid_f := 1969;
        ELSIF x = 6595 THEN
            sigmoid_f := 1969;
        ELSIF x = 6596 THEN
            sigmoid_f := 1969;
        ELSIF x = 6597 THEN
            sigmoid_f := 1969;
        ELSIF x = 6598 THEN
            sigmoid_f := 1969;
        ELSIF x = 6599 THEN
            sigmoid_f := 1969;
        ELSIF x = 6600 THEN
            sigmoid_f := 1969;
        ELSIF x = 6601 THEN
            sigmoid_f := 1969;
        ELSIF x = 6602 THEN
            sigmoid_f := 1969;
        ELSIF x = 6603 THEN
            sigmoid_f := 1969;
        ELSIF x = 6604 THEN
            sigmoid_f := 1969;
        ELSIF x = 6605 THEN
            sigmoid_f := 1969;
        ELSIF x = 6606 THEN
            sigmoid_f := 1969;
        ELSIF x = 6607 THEN
            sigmoid_f := 1969;
        ELSIF x = 6608 THEN
            sigmoid_f := 1970;
        ELSIF x = 6609 THEN
            sigmoid_f := 1970;
        ELSIF x = 6610 THEN
            sigmoid_f := 1970;
        ELSIF x = 6611 THEN
            sigmoid_f := 1970;
        ELSIF x = 6612 THEN
            sigmoid_f := 1970;
        ELSIF x = 6613 THEN
            sigmoid_f := 1970;
        ELSIF x = 6614 THEN
            sigmoid_f := 1970;
        ELSIF x = 6615 THEN
            sigmoid_f := 1970;
        ELSIF x = 6616 THEN
            sigmoid_f := 1970;
        ELSIF x = 6617 THEN
            sigmoid_f := 1970;
        ELSIF x = 6618 THEN
            sigmoid_f := 1970;
        ELSIF x = 6619 THEN
            sigmoid_f := 1970;
        ELSIF x = 6620 THEN
            sigmoid_f := 1970;
        ELSIF x = 6621 THEN
            sigmoid_f := 1970;
        ELSIF x = 6622 THEN
            sigmoid_f := 1970;
        ELSIF x = 6623 THEN
            sigmoid_f := 1970;
        ELSIF x = 6624 THEN
            sigmoid_f := 1970;
        ELSIF x = 6625 THEN
            sigmoid_f := 1970;
        ELSIF x = 6626 THEN
            sigmoid_f := 1970;
        ELSIF x = 6627 THEN
            sigmoid_f := 1970;
        ELSIF x = 6628 THEN
            sigmoid_f := 1970;
        ELSIF x = 6629 THEN
            sigmoid_f := 1970;
        ELSIF x = 6630 THEN
            sigmoid_f := 1970;
        ELSIF x = 6631 THEN
            sigmoid_f := 1970;
        ELSIF x = 6632 THEN
            sigmoid_f := 1971;
        ELSIF x = 6633 THEN
            sigmoid_f := 1971;
        ELSIF x = 6634 THEN
            sigmoid_f := 1971;
        ELSIF x = 6635 THEN
            sigmoid_f := 1971;
        ELSIF x = 6636 THEN
            sigmoid_f := 1971;
        ELSIF x = 6637 THEN
            sigmoid_f := 1971;
        ELSIF x = 6638 THEN
            sigmoid_f := 1971;
        ELSIF x = 6639 THEN
            sigmoid_f := 1971;
        ELSIF x = 6640 THEN
            sigmoid_f := 1971;
        ELSIF x = 6641 THEN
            sigmoid_f := 1971;
        ELSIF x = 6642 THEN
            sigmoid_f := 1971;
        ELSIF x = 6643 THEN
            sigmoid_f := 1971;
        ELSIF x = 6644 THEN
            sigmoid_f := 1971;
        ELSIF x = 6645 THEN
            sigmoid_f := 1971;
        ELSIF x = 6646 THEN
            sigmoid_f := 1971;
        ELSIF x = 6647 THEN
            sigmoid_f := 1971;
        ELSIF x = 6648 THEN
            sigmoid_f := 1971;
        ELSIF x = 6649 THEN
            sigmoid_f := 1971;
        ELSIF x = 6650 THEN
            sigmoid_f := 1971;
        ELSIF x = 6651 THEN
            sigmoid_f := 1971;
        ELSIF x = 6652 THEN
            sigmoid_f := 1971;
        ELSIF x = 6653 THEN
            sigmoid_f := 1971;
        ELSIF x = 6654 THEN
            sigmoid_f := 1971;
        ELSIF x = 6655 THEN
            sigmoid_f := 1971;
        ELSIF x = 6656 THEN
            sigmoid_f := 1972;
        ELSIF x = 6657 THEN
            sigmoid_f := 1972;
        ELSIF x = 6658 THEN
            sigmoid_f := 1972;
        ELSIF x = 6659 THEN
            sigmoid_f := 1972;
        ELSIF x = 6660 THEN
            sigmoid_f := 1972;
        ELSIF x = 6661 THEN
            sigmoid_f := 1972;
        ELSIF x = 6662 THEN
            sigmoid_f := 1972;
        ELSIF x = 6663 THEN
            sigmoid_f := 1972;
        ELSIF x = 6664 THEN
            sigmoid_f := 1972;
        ELSIF x = 6665 THEN
            sigmoid_f := 1972;
        ELSIF x = 6666 THEN
            sigmoid_f := 1972;
        ELSIF x = 6667 THEN
            sigmoid_f := 1972;
        ELSIF x = 6668 THEN
            sigmoid_f := 1972;
        ELSIF x = 6669 THEN
            sigmoid_f := 1972;
        ELSIF x = 6670 THEN
            sigmoid_f := 1972;
        ELSIF x = 6671 THEN
            sigmoid_f := 1972;
        ELSIF x = 6672 THEN
            sigmoid_f := 1972;
        ELSIF x = 6673 THEN
            sigmoid_f := 1972;
        ELSIF x = 6674 THEN
            sigmoid_f := 1972;
        ELSIF x = 6675 THEN
            sigmoid_f := 1972;
        ELSIF x = 6676 THEN
            sigmoid_f := 1972;
        ELSIF x = 6677 THEN
            sigmoid_f := 1972;
        ELSIF x = 6678 THEN
            sigmoid_f := 1972;
        ELSIF x = 6679 THEN
            sigmoid_f := 1972;
        ELSIF x = 6680 THEN
            sigmoid_f := 1972;
        ELSIF x = 6681 THEN
            sigmoid_f := 1972;
        ELSIF x = 6682 THEN
            sigmoid_f := 1972;
        ELSIF x = 6683 THEN
            sigmoid_f := 1972;
        ELSIF x = 6684 THEN
            sigmoid_f := 1972;
        ELSIF x = 6685 THEN
            sigmoid_f := 1972;
        ELSIF x = 6686 THEN
            sigmoid_f := 1972;
        ELSIF x = 6687 THEN
            sigmoid_f := 1972;
        ELSIF x = 6688 THEN
            sigmoid_f := 1973;
        ELSIF x = 6689 THEN
            sigmoid_f := 1973;
        ELSIF x = 6690 THEN
            sigmoid_f := 1973;
        ELSIF x = 6691 THEN
            sigmoid_f := 1973;
        ELSIF x = 6692 THEN
            sigmoid_f := 1973;
        ELSIF x = 6693 THEN
            sigmoid_f := 1973;
        ELSIF x = 6694 THEN
            sigmoid_f := 1973;
        ELSIF x = 6695 THEN
            sigmoid_f := 1973;
        ELSIF x = 6696 THEN
            sigmoid_f := 1973;
        ELSIF x = 6697 THEN
            sigmoid_f := 1973;
        ELSIF x = 6698 THEN
            sigmoid_f := 1973;
        ELSIF x = 6699 THEN
            sigmoid_f := 1973;
        ELSIF x = 6700 THEN
            sigmoid_f := 1973;
        ELSIF x = 6701 THEN
            sigmoid_f := 1973;
        ELSIF x = 6702 THEN
            sigmoid_f := 1973;
        ELSIF x = 6703 THEN
            sigmoid_f := 1973;
        ELSIF x = 6704 THEN
            sigmoid_f := 1973;
        ELSIF x = 6705 THEN
            sigmoid_f := 1973;
        ELSIF x = 6706 THEN
            sigmoid_f := 1973;
        ELSIF x = 6707 THEN
            sigmoid_f := 1973;
        ELSIF x = 6708 THEN
            sigmoid_f := 1973;
        ELSIF x = 6709 THEN
            sigmoid_f := 1973;
        ELSIF x = 6710 THEN
            sigmoid_f := 1973;
        ELSIF x = 6711 THEN
            sigmoid_f := 1973;
        ELSIF x = 6712 THEN
            sigmoid_f := 1973;
        ELSIF x = 6713 THEN
            sigmoid_f := 1973;
        ELSIF x = 6714 THEN
            sigmoid_f := 1973;
        ELSIF x = 6715 THEN
            sigmoid_f := 1973;
        ELSIF x = 6716 THEN
            sigmoid_f := 1973;
        ELSIF x = 6717 THEN
            sigmoid_f := 1973;
        ELSIF x = 6718 THEN
            sigmoid_f := 1973;
        ELSIF x = 6719 THEN
            sigmoid_f := 1973;
        ELSIF x = 6720 THEN
            sigmoid_f := 1974;
        ELSIF x = 6721 THEN
            sigmoid_f := 1974;
        ELSIF x = 6722 THEN
            sigmoid_f := 1974;
        ELSIF x = 6723 THEN
            sigmoid_f := 1974;
        ELSIF x = 6724 THEN
            sigmoid_f := 1974;
        ELSIF x = 6725 THEN
            sigmoid_f := 1974;
        ELSIF x = 6726 THEN
            sigmoid_f := 1974;
        ELSIF x = 6727 THEN
            sigmoid_f := 1974;
        ELSIF x = 6728 THEN
            sigmoid_f := 1974;
        ELSIF x = 6729 THEN
            sigmoid_f := 1974;
        ELSIF x = 6730 THEN
            sigmoid_f := 1974;
        ELSIF x = 6731 THEN
            sigmoid_f := 1974;
        ELSIF x = 6732 THEN
            sigmoid_f := 1974;
        ELSIF x = 6733 THEN
            sigmoid_f := 1974;
        ELSIF x = 6734 THEN
            sigmoid_f := 1974;
        ELSIF x = 6735 THEN
            sigmoid_f := 1974;
        ELSIF x = 6736 THEN
            sigmoid_f := 1974;
        ELSIF x = 6737 THEN
            sigmoid_f := 1974;
        ELSIF x = 6738 THEN
            sigmoid_f := 1974;
        ELSIF x = 6739 THEN
            sigmoid_f := 1974;
        ELSIF x = 6740 THEN
            sigmoid_f := 1974;
        ELSIF x = 6741 THEN
            sigmoid_f := 1974;
        ELSIF x = 6742 THEN
            sigmoid_f := 1974;
        ELSIF x = 6743 THEN
            sigmoid_f := 1974;
        ELSIF x = 6744 THEN
            sigmoid_f := 1974;
        ELSIF x = 6745 THEN
            sigmoid_f := 1974;
        ELSIF x = 6746 THEN
            sigmoid_f := 1974;
        ELSIF x = 6747 THEN
            sigmoid_f := 1974;
        ELSIF x = 6748 THEN
            sigmoid_f := 1974;
        ELSIF x = 6749 THEN
            sigmoid_f := 1974;
        ELSIF x = 6750 THEN
            sigmoid_f := 1974;
        ELSIF x = 6751 THEN
            sigmoid_f := 1974;
        ELSIF x = 6752 THEN
            sigmoid_f := 1975;
        ELSIF x = 6753 THEN
            sigmoid_f := 1975;
        ELSIF x = 6754 THEN
            sigmoid_f := 1975;
        ELSIF x = 6755 THEN
            sigmoid_f := 1975;
        ELSIF x = 6756 THEN
            sigmoid_f := 1975;
        ELSIF x = 6757 THEN
            sigmoid_f := 1975;
        ELSIF x = 6758 THEN
            sigmoid_f := 1975;
        ELSIF x = 6759 THEN
            sigmoid_f := 1975;
        ELSIF x = 6760 THEN
            sigmoid_f := 1975;
        ELSIF x = 6761 THEN
            sigmoid_f := 1975;
        ELSIF x = 6762 THEN
            sigmoid_f := 1975;
        ELSIF x = 6763 THEN
            sigmoid_f := 1975;
        ELSIF x = 6764 THEN
            sigmoid_f := 1975;
        ELSIF x = 6765 THEN
            sigmoid_f := 1975;
        ELSIF x = 6766 THEN
            sigmoid_f := 1975;
        ELSIF x = 6767 THEN
            sigmoid_f := 1975;
        ELSIF x = 6768 THEN
            sigmoid_f := 1975;
        ELSIF x = 6769 THEN
            sigmoid_f := 1975;
        ELSIF x = 6770 THEN
            sigmoid_f := 1975;
        ELSIF x = 6771 THEN
            sigmoid_f := 1975;
        ELSIF x = 6772 THEN
            sigmoid_f := 1975;
        ELSIF x = 6773 THEN
            sigmoid_f := 1975;
        ELSIF x = 6774 THEN
            sigmoid_f := 1975;
        ELSIF x = 6775 THEN
            sigmoid_f := 1975;
        ELSIF x = 6776 THEN
            sigmoid_f := 1975;
        ELSIF x = 6777 THEN
            sigmoid_f := 1975;
        ELSIF x = 6778 THEN
            sigmoid_f := 1975;
        ELSIF x = 6779 THEN
            sigmoid_f := 1975;
        ELSIF x = 6780 THEN
            sigmoid_f := 1975;
        ELSIF x = 6781 THEN
            sigmoid_f := 1975;
        ELSIF x = 6782 THEN
            sigmoid_f := 1975;
        ELSIF x = 6783 THEN
            sigmoid_f := 1975;
        ELSIF x = 6784 THEN
            sigmoid_f := 1976;
        ELSIF x = 6785 THEN
            sigmoid_f := 1976;
        ELSIF x = 6786 THEN
            sigmoid_f := 1976;
        ELSIF x = 6787 THEN
            sigmoid_f := 1976;
        ELSIF x = 6788 THEN
            sigmoid_f := 1976;
        ELSIF x = 6789 THEN
            sigmoid_f := 1976;
        ELSIF x = 6790 THEN
            sigmoid_f := 1976;
        ELSIF x = 6791 THEN
            sigmoid_f := 1976;
        ELSIF x = 6792 THEN
            sigmoid_f := 1976;
        ELSIF x = 6793 THEN
            sigmoid_f := 1976;
        ELSIF x = 6794 THEN
            sigmoid_f := 1976;
        ELSIF x = 6795 THEN
            sigmoid_f := 1976;
        ELSIF x = 6796 THEN
            sigmoid_f := 1976;
        ELSIF x = 6797 THEN
            sigmoid_f := 1976;
        ELSIF x = 6798 THEN
            sigmoid_f := 1976;
        ELSIF x = 6799 THEN
            sigmoid_f := 1976;
        ELSIF x = 6800 THEN
            sigmoid_f := 1976;
        ELSIF x = 6801 THEN
            sigmoid_f := 1976;
        ELSIF x = 6802 THEN
            sigmoid_f := 1976;
        ELSIF x = 6803 THEN
            sigmoid_f := 1976;
        ELSIF x = 6804 THEN
            sigmoid_f := 1976;
        ELSIF x = 6805 THEN
            sigmoid_f := 1976;
        ELSIF x = 6806 THEN
            sigmoid_f := 1976;
        ELSIF x = 6807 THEN
            sigmoid_f := 1976;
        ELSIF x = 6808 THEN
            sigmoid_f := 1976;
        ELSIF x = 6809 THEN
            sigmoid_f := 1976;
        ELSIF x = 6810 THEN
            sigmoid_f := 1976;
        ELSIF x = 6811 THEN
            sigmoid_f := 1976;
        ELSIF x = 6812 THEN
            sigmoid_f := 1976;
        ELSIF x = 6813 THEN
            sigmoid_f := 1976;
        ELSIF x = 6814 THEN
            sigmoid_f := 1976;
        ELSIF x = 6815 THEN
            sigmoid_f := 1976;
        ELSIF x = 6816 THEN
            sigmoid_f := 1977;
        ELSIF x = 6817 THEN
            sigmoid_f := 1977;
        ELSIF x = 6818 THEN
            sigmoid_f := 1977;
        ELSIF x = 6819 THEN
            sigmoid_f := 1977;
        ELSIF x = 6820 THEN
            sigmoid_f := 1977;
        ELSIF x = 6821 THEN
            sigmoid_f := 1977;
        ELSIF x = 6822 THEN
            sigmoid_f := 1977;
        ELSIF x = 6823 THEN
            sigmoid_f := 1977;
        ELSIF x = 6824 THEN
            sigmoid_f := 1977;
        ELSIF x = 6825 THEN
            sigmoid_f := 1977;
        ELSIF x = 6826 THEN
            sigmoid_f := 1977;
        ELSIF x = 6827 THEN
            sigmoid_f := 1977;
        ELSIF x = 6828 THEN
            sigmoid_f := 1977;
        ELSIF x = 6829 THEN
            sigmoid_f := 1977;
        ELSIF x = 6830 THEN
            sigmoid_f := 1977;
        ELSIF x = 6831 THEN
            sigmoid_f := 1977;
        ELSIF x = 6832 THEN
            sigmoid_f := 1977;
        ELSIF x = 6833 THEN
            sigmoid_f := 1977;
        ELSIF x = 6834 THEN
            sigmoid_f := 1977;
        ELSIF x = 6835 THEN
            sigmoid_f := 1977;
        ELSIF x = 6836 THEN
            sigmoid_f := 1977;
        ELSIF x = 6837 THEN
            sigmoid_f := 1977;
        ELSIF x = 6838 THEN
            sigmoid_f := 1977;
        ELSIF x = 6839 THEN
            sigmoid_f := 1977;
        ELSIF x = 6840 THEN
            sigmoid_f := 1977;
        ELSIF x = 6841 THEN
            sigmoid_f := 1977;
        ELSIF x = 6842 THEN
            sigmoid_f := 1977;
        ELSIF x = 6843 THEN
            sigmoid_f := 1977;
        ELSIF x = 6844 THEN
            sigmoid_f := 1977;
        ELSIF x = 6845 THEN
            sigmoid_f := 1977;
        ELSIF x = 6846 THEN
            sigmoid_f := 1977;
        ELSIF x = 6847 THEN
            sigmoid_f := 1977;
        ELSIF x = 6848 THEN
            sigmoid_f := 1978;
        ELSIF x = 6849 THEN
            sigmoid_f := 1978;
        ELSIF x = 6850 THEN
            sigmoid_f := 1978;
        ELSIF x = 6851 THEN
            sigmoid_f := 1978;
        ELSIF x = 6852 THEN
            sigmoid_f := 1978;
        ELSIF x = 6853 THEN
            sigmoid_f := 1978;
        ELSIF x = 6854 THEN
            sigmoid_f := 1978;
        ELSIF x = 6855 THEN
            sigmoid_f := 1978;
        ELSIF x = 6856 THEN
            sigmoid_f := 1978;
        ELSIF x = 6857 THEN
            sigmoid_f := 1978;
        ELSIF x = 6858 THEN
            sigmoid_f := 1978;
        ELSIF x = 6859 THEN
            sigmoid_f := 1978;
        ELSIF x = 6860 THEN
            sigmoid_f := 1978;
        ELSIF x = 6861 THEN
            sigmoid_f := 1978;
        ELSIF x = 6862 THEN
            sigmoid_f := 1978;
        ELSIF x = 6863 THEN
            sigmoid_f := 1978;
        ELSIF x = 6864 THEN
            sigmoid_f := 1978;
        ELSIF x = 6865 THEN
            sigmoid_f := 1978;
        ELSIF x = 6866 THEN
            sigmoid_f := 1978;
        ELSIF x = 6867 THEN
            sigmoid_f := 1978;
        ELSIF x = 6868 THEN
            sigmoid_f := 1978;
        ELSIF x = 6869 THEN
            sigmoid_f := 1978;
        ELSIF x = 6870 THEN
            sigmoid_f := 1978;
        ELSIF x = 6871 THEN
            sigmoid_f := 1978;
        ELSIF x = 6872 THEN
            sigmoid_f := 1978;
        ELSIF x = 6873 THEN
            sigmoid_f := 1978;
        ELSIF x = 6874 THEN
            sigmoid_f := 1978;
        ELSIF x = 6875 THEN
            sigmoid_f := 1978;
        ELSIF x = 6876 THEN
            sigmoid_f := 1978;
        ELSIF x = 6877 THEN
            sigmoid_f := 1978;
        ELSIF x = 6878 THEN
            sigmoid_f := 1978;
        ELSIF x = 6879 THEN
            sigmoid_f := 1978;
        ELSIF x = 6880 THEN
            sigmoid_f := 1979;
        ELSIF x = 6881 THEN
            sigmoid_f := 1979;
        ELSIF x = 6882 THEN
            sigmoid_f := 1979;
        ELSIF x = 6883 THEN
            sigmoid_f := 1979;
        ELSIF x = 6884 THEN
            sigmoid_f := 1979;
        ELSIF x = 6885 THEN
            sigmoid_f := 1979;
        ELSIF x = 6886 THEN
            sigmoid_f := 1979;
        ELSIF x = 6887 THEN
            sigmoid_f := 1979;
        ELSIF x = 6888 THEN
            sigmoid_f := 1979;
        ELSIF x = 6889 THEN
            sigmoid_f := 1979;
        ELSIF x = 6890 THEN
            sigmoid_f := 1979;
        ELSIF x = 6891 THEN
            sigmoid_f := 1979;
        ELSIF x = 6892 THEN
            sigmoid_f := 1979;
        ELSIF x = 6893 THEN
            sigmoid_f := 1979;
        ELSIF x = 6894 THEN
            sigmoid_f := 1979;
        ELSIF x = 6895 THEN
            sigmoid_f := 1979;
        ELSIF x = 6896 THEN
            sigmoid_f := 1979;
        ELSIF x = 6897 THEN
            sigmoid_f := 1979;
        ELSIF x = 6898 THEN
            sigmoid_f := 1979;
        ELSIF x = 6899 THEN
            sigmoid_f := 1979;
        ELSIF x = 6900 THEN
            sigmoid_f := 1979;
        ELSIF x = 6901 THEN
            sigmoid_f := 1979;
        ELSIF x = 6902 THEN
            sigmoid_f := 1979;
        ELSIF x = 6903 THEN
            sigmoid_f := 1979;
        ELSIF x = 6904 THEN
            sigmoid_f := 1979;
        ELSIF x = 6905 THEN
            sigmoid_f := 1979;
        ELSIF x = 6906 THEN
            sigmoid_f := 1979;
        ELSIF x = 6907 THEN
            sigmoid_f := 1979;
        ELSIF x = 6908 THEN
            sigmoid_f := 1979;
        ELSIF x = 6909 THEN
            sigmoid_f := 1979;
        ELSIF x = 6910 THEN
            sigmoid_f := 1979;
        ELSIF x = 6911 THEN
            sigmoid_f := 1979;
        ELSIF x = 6912 THEN
            sigmoid_f := 1980;
        ELSIF x = 6913 THEN
            sigmoid_f := 1980;
        ELSIF x = 6914 THEN
            sigmoid_f := 1980;
        ELSIF x = 6915 THEN
            sigmoid_f := 1980;
        ELSIF x = 6916 THEN
            sigmoid_f := 1980;
        ELSIF x = 6917 THEN
            sigmoid_f := 1980;
        ELSIF x = 6918 THEN
            sigmoid_f := 1980;
        ELSIF x = 6919 THEN
            sigmoid_f := 1980;
        ELSIF x = 6920 THEN
            sigmoid_f := 1980;
        ELSIF x = 6921 THEN
            sigmoid_f := 1980;
        ELSIF x = 6922 THEN
            sigmoid_f := 1980;
        ELSIF x = 6923 THEN
            sigmoid_f := 1980;
        ELSIF x = 6924 THEN
            sigmoid_f := 1980;
        ELSIF x = 6925 THEN
            sigmoid_f := 1980;
        ELSIF x = 6926 THEN
            sigmoid_f := 1980;
        ELSIF x = 6927 THEN
            sigmoid_f := 1980;
        ELSIF x = 6928 THEN
            sigmoid_f := 1980;
        ELSIF x = 6929 THEN
            sigmoid_f := 1980;
        ELSIF x = 6930 THEN
            sigmoid_f := 1980;
        ELSIF x = 6931 THEN
            sigmoid_f := 1980;
        ELSIF x = 6932 THEN
            sigmoid_f := 1980;
        ELSIF x = 6933 THEN
            sigmoid_f := 1980;
        ELSIF x = 6934 THEN
            sigmoid_f := 1980;
        ELSIF x = 6935 THEN
            sigmoid_f := 1980;
        ELSIF x = 6936 THEN
            sigmoid_f := 1980;
        ELSIF x = 6937 THEN
            sigmoid_f := 1980;
        ELSIF x = 6938 THEN
            sigmoid_f := 1980;
        ELSIF x = 6939 THEN
            sigmoid_f := 1980;
        ELSIF x = 6940 THEN
            sigmoid_f := 1980;
        ELSIF x = 6941 THEN
            sigmoid_f := 1980;
        ELSIF x = 6942 THEN
            sigmoid_f := 1980;
        ELSIF x = 6943 THEN
            sigmoid_f := 1980;
        ELSIF x = 6944 THEN
            sigmoid_f := 1981;
        ELSIF x = 6945 THEN
            sigmoid_f := 1981;
        ELSIF x = 6946 THEN
            sigmoid_f := 1981;
        ELSIF x = 6947 THEN
            sigmoid_f := 1981;
        ELSIF x = 6948 THEN
            sigmoid_f := 1981;
        ELSIF x = 6949 THEN
            sigmoid_f := 1981;
        ELSIF x = 6950 THEN
            sigmoid_f := 1981;
        ELSIF x = 6951 THEN
            sigmoid_f := 1981;
        ELSIF x = 6952 THEN
            sigmoid_f := 1981;
        ELSIF x = 6953 THEN
            sigmoid_f := 1981;
        ELSIF x = 6954 THEN
            sigmoid_f := 1981;
        ELSIF x = 6955 THEN
            sigmoid_f := 1981;
        ELSIF x = 6956 THEN
            sigmoid_f := 1981;
        ELSIF x = 6957 THEN
            sigmoid_f := 1981;
        ELSIF x = 6958 THEN
            sigmoid_f := 1981;
        ELSIF x = 6959 THEN
            sigmoid_f := 1981;
        ELSIF x = 6960 THEN
            sigmoid_f := 1981;
        ELSIF x = 6961 THEN
            sigmoid_f := 1981;
        ELSIF x = 6962 THEN
            sigmoid_f := 1981;
        ELSIF x = 6963 THEN
            sigmoid_f := 1981;
        ELSIF x = 6964 THEN
            sigmoid_f := 1981;
        ELSIF x = 6965 THEN
            sigmoid_f := 1981;
        ELSIF x = 6966 THEN
            sigmoid_f := 1981;
        ELSIF x = 6967 THEN
            sigmoid_f := 1981;
        ELSIF x = 6968 THEN
            sigmoid_f := 1981;
        ELSIF x = 6969 THEN
            sigmoid_f := 1981;
        ELSIF x = 6970 THEN
            sigmoid_f := 1981;
        ELSIF x = 6971 THEN
            sigmoid_f := 1981;
        ELSIF x = 6972 THEN
            sigmoid_f := 1981;
        ELSIF x = 6973 THEN
            sigmoid_f := 1981;
        ELSIF x = 6974 THEN
            sigmoid_f := 1981;
        ELSIF x = 6975 THEN
            sigmoid_f := 1981;
        ELSIF x = 6976 THEN
            sigmoid_f := 1982;
        ELSIF x = 6977 THEN
            sigmoid_f := 1982;
        ELSIF x = 6978 THEN
            sigmoid_f := 1982;
        ELSIF x = 6979 THEN
            sigmoid_f := 1982;
        ELSIF x = 6980 THEN
            sigmoid_f := 1982;
        ELSIF x = 6981 THEN
            sigmoid_f := 1982;
        ELSIF x = 6982 THEN
            sigmoid_f := 1982;
        ELSIF x = 6983 THEN
            sigmoid_f := 1982;
        ELSIF x = 6984 THEN
            sigmoid_f := 1982;
        ELSIF x = 6985 THEN
            sigmoid_f := 1982;
        ELSIF x = 6986 THEN
            sigmoid_f := 1982;
        ELSIF x = 6987 THEN
            sigmoid_f := 1982;
        ELSIF x = 6988 THEN
            sigmoid_f := 1982;
        ELSIF x = 6989 THEN
            sigmoid_f := 1982;
        ELSIF x = 6990 THEN
            sigmoid_f := 1982;
        ELSIF x = 6991 THEN
            sigmoid_f := 1982;
        ELSIF x = 6992 THEN
            sigmoid_f := 1982;
        ELSIF x = 6993 THEN
            sigmoid_f := 1982;
        ELSIF x = 6994 THEN
            sigmoid_f := 1982;
        ELSIF x = 6995 THEN
            sigmoid_f := 1982;
        ELSIF x = 6996 THEN
            sigmoid_f := 1982;
        ELSIF x = 6997 THEN
            sigmoid_f := 1982;
        ELSIF x = 6998 THEN
            sigmoid_f := 1982;
        ELSIF x = 6999 THEN
            sigmoid_f := 1982;
        ELSIF x = 7000 THEN
            sigmoid_f := 1982;
        ELSIF x = 7001 THEN
            sigmoid_f := 1982;
        ELSIF x = 7002 THEN
            sigmoid_f := 1982;
        ELSIF x = 7003 THEN
            sigmoid_f := 1982;
        ELSIF x = 7004 THEN
            sigmoid_f := 1982;
        ELSIF x = 7005 THEN
            sigmoid_f := 1982;
        ELSIF x = 7006 THEN
            sigmoid_f := 1982;
        ELSIF x = 7007 THEN
            sigmoid_f := 1982;
        ELSIF x = 7008 THEN
            sigmoid_f := 1983;
        ELSIF x = 7009 THEN
            sigmoid_f := 1983;
        ELSIF x = 7010 THEN
            sigmoid_f := 1983;
        ELSIF x = 7011 THEN
            sigmoid_f := 1983;
        ELSIF x = 7012 THEN
            sigmoid_f := 1983;
        ELSIF x = 7013 THEN
            sigmoid_f := 1983;
        ELSIF x = 7014 THEN
            sigmoid_f := 1983;
        ELSIF x = 7015 THEN
            sigmoid_f := 1983;
        ELSIF x = 7016 THEN
            sigmoid_f := 1983;
        ELSIF x = 7017 THEN
            sigmoid_f := 1983;
        ELSIF x = 7018 THEN
            sigmoid_f := 1983;
        ELSIF x = 7019 THEN
            sigmoid_f := 1983;
        ELSIF x = 7020 THEN
            sigmoid_f := 1983;
        ELSIF x = 7021 THEN
            sigmoid_f := 1983;
        ELSIF x = 7022 THEN
            sigmoid_f := 1983;
        ELSIF x = 7023 THEN
            sigmoid_f := 1983;
        ELSIF x = 7024 THEN
            sigmoid_f := 1983;
        ELSIF x = 7025 THEN
            sigmoid_f := 1983;
        ELSIF x = 7026 THEN
            sigmoid_f := 1983;
        ELSIF x = 7027 THEN
            sigmoid_f := 1983;
        ELSIF x = 7028 THEN
            sigmoid_f := 1983;
        ELSIF x = 7029 THEN
            sigmoid_f := 1983;
        ELSIF x = 7030 THEN
            sigmoid_f := 1983;
        ELSIF x = 7031 THEN
            sigmoid_f := 1983;
        ELSIF x = 7032 THEN
            sigmoid_f := 1983;
        ELSIF x = 7033 THEN
            sigmoid_f := 1983;
        ELSIF x = 7034 THEN
            sigmoid_f := 1983;
        ELSIF x = 7035 THEN
            sigmoid_f := 1983;
        ELSIF x = 7036 THEN
            sigmoid_f := 1983;
        ELSIF x = 7037 THEN
            sigmoid_f := 1983;
        ELSIF x = 7038 THEN
            sigmoid_f := 1983;
        ELSIF x = 7039 THEN
            sigmoid_f := 1983;
        ELSIF x = 7040 THEN
            sigmoid_f := 1984;
        ELSIF x = 7041 THEN
            sigmoid_f := 1984;
        ELSIF x = 7042 THEN
            sigmoid_f := 1984;
        ELSIF x = 7043 THEN
            sigmoid_f := 1984;
        ELSIF x = 7044 THEN
            sigmoid_f := 1984;
        ELSIF x = 7045 THEN
            sigmoid_f := 1984;
        ELSIF x = 7046 THEN
            sigmoid_f := 1984;
        ELSIF x = 7047 THEN
            sigmoid_f := 1984;
        ELSIF x = 7048 THEN
            sigmoid_f := 1984;
        ELSIF x = 7049 THEN
            sigmoid_f := 1984;
        ELSIF x = 7050 THEN
            sigmoid_f := 1984;
        ELSIF x = 7051 THEN
            sigmoid_f := 1984;
        ELSIF x = 7052 THEN
            sigmoid_f := 1984;
        ELSIF x = 7053 THEN
            sigmoid_f := 1984;
        ELSIF x = 7054 THEN
            sigmoid_f := 1984;
        ELSIF x = 7055 THEN
            sigmoid_f := 1984;
        ELSIF x = 7056 THEN
            sigmoid_f := 1984;
        ELSIF x = 7057 THEN
            sigmoid_f := 1984;
        ELSIF x = 7058 THEN
            sigmoid_f := 1984;
        ELSIF x = 7059 THEN
            sigmoid_f := 1984;
        ELSIF x = 7060 THEN
            sigmoid_f := 1984;
        ELSIF x = 7061 THEN
            sigmoid_f := 1984;
        ELSIF x = 7062 THEN
            sigmoid_f := 1984;
        ELSIF x = 7063 THEN
            sigmoid_f := 1984;
        ELSIF x = 7064 THEN
            sigmoid_f := 1984;
        ELSIF x = 7065 THEN
            sigmoid_f := 1984;
        ELSIF x = 7066 THEN
            sigmoid_f := 1984;
        ELSIF x = 7067 THEN
            sigmoid_f := 1984;
        ELSIF x = 7068 THEN
            sigmoid_f := 1984;
        ELSIF x = 7069 THEN
            sigmoid_f := 1984;
        ELSIF x = 7070 THEN
            sigmoid_f := 1984;
        ELSIF x = 7071 THEN
            sigmoid_f := 1984;
        ELSIF x = 7072 THEN
            sigmoid_f := 1985;
        ELSIF x = 7073 THEN
            sigmoid_f := 1985;
        ELSIF x = 7074 THEN
            sigmoid_f := 1985;
        ELSIF x = 7075 THEN
            sigmoid_f := 1985;
        ELSIF x = 7076 THEN
            sigmoid_f := 1985;
        ELSIF x = 7077 THEN
            sigmoid_f := 1985;
        ELSIF x = 7078 THEN
            sigmoid_f := 1985;
        ELSIF x = 7079 THEN
            sigmoid_f := 1985;
        ELSIF x = 7080 THEN
            sigmoid_f := 1985;
        ELSIF x = 7081 THEN
            sigmoid_f := 1985;
        ELSIF x = 7082 THEN
            sigmoid_f := 1985;
        ELSIF x = 7083 THEN
            sigmoid_f := 1985;
        ELSIF x = 7084 THEN
            sigmoid_f := 1985;
        ELSIF x = 7085 THEN
            sigmoid_f := 1985;
        ELSIF x = 7086 THEN
            sigmoid_f := 1985;
        ELSIF x = 7087 THEN
            sigmoid_f := 1985;
        ELSIF x = 7088 THEN
            sigmoid_f := 1985;
        ELSIF x = 7089 THEN
            sigmoid_f := 1985;
        ELSIF x = 7090 THEN
            sigmoid_f := 1985;
        ELSIF x = 7091 THEN
            sigmoid_f := 1985;
        ELSIF x = 7092 THEN
            sigmoid_f := 1985;
        ELSIF x = 7093 THEN
            sigmoid_f := 1985;
        ELSIF x = 7094 THEN
            sigmoid_f := 1985;
        ELSIF x = 7095 THEN
            sigmoid_f := 1985;
        ELSIF x = 7096 THEN
            sigmoid_f := 1985;
        ELSIF x = 7097 THEN
            sigmoid_f := 1985;
        ELSIF x = 7098 THEN
            sigmoid_f := 1985;
        ELSIF x = 7099 THEN
            sigmoid_f := 1985;
        ELSIF x = 7100 THEN
            sigmoid_f := 1985;
        ELSIF x = 7101 THEN
            sigmoid_f := 1985;
        ELSIF x = 7102 THEN
            sigmoid_f := 1985;
        ELSIF x = 7103 THEN
            sigmoid_f := 1985;
        ELSIF x = 7104 THEN
            sigmoid_f := 1986;
        ELSIF x = 7105 THEN
            sigmoid_f := 1986;
        ELSIF x = 7106 THEN
            sigmoid_f := 1986;
        ELSIF x = 7107 THEN
            sigmoid_f := 1986;
        ELSIF x = 7108 THEN
            sigmoid_f := 1986;
        ELSIF x = 7109 THEN
            sigmoid_f := 1986;
        ELSIF x = 7110 THEN
            sigmoid_f := 1986;
        ELSIF x = 7111 THEN
            sigmoid_f := 1986;
        ELSIF x = 7112 THEN
            sigmoid_f := 1986;
        ELSIF x = 7113 THEN
            sigmoid_f := 1986;
        ELSIF x = 7114 THEN
            sigmoid_f := 1986;
        ELSIF x = 7115 THEN
            sigmoid_f := 1986;
        ELSIF x = 7116 THEN
            sigmoid_f := 1986;
        ELSIF x = 7117 THEN
            sigmoid_f := 1986;
        ELSIF x = 7118 THEN
            sigmoid_f := 1986;
        ELSIF x = 7119 THEN
            sigmoid_f := 1986;
        ELSIF x = 7120 THEN
            sigmoid_f := 1986;
        ELSIF x = 7121 THEN
            sigmoid_f := 1986;
        ELSIF x = 7122 THEN
            sigmoid_f := 1986;
        ELSIF x = 7123 THEN
            sigmoid_f := 1986;
        ELSIF x = 7124 THEN
            sigmoid_f := 1986;
        ELSIF x = 7125 THEN
            sigmoid_f := 1986;
        ELSIF x = 7126 THEN
            sigmoid_f := 1986;
        ELSIF x = 7127 THEN
            sigmoid_f := 1986;
        ELSIF x = 7128 THEN
            sigmoid_f := 1986;
        ELSIF x = 7129 THEN
            sigmoid_f := 1986;
        ELSIF x = 7130 THEN
            sigmoid_f := 1986;
        ELSIF x = 7131 THEN
            sigmoid_f := 1986;
        ELSIF x = 7132 THEN
            sigmoid_f := 1986;
        ELSIF x = 7133 THEN
            sigmoid_f := 1986;
        ELSIF x = 7134 THEN
            sigmoid_f := 1986;
        ELSIF x = 7135 THEN
            sigmoid_f := 1986;
        ELSIF x = 7136 THEN
            sigmoid_f := 1987;
        ELSIF x = 7137 THEN
            sigmoid_f := 1987;
        ELSIF x = 7138 THEN
            sigmoid_f := 1987;
        ELSIF x = 7139 THEN
            sigmoid_f := 1987;
        ELSIF x = 7140 THEN
            sigmoid_f := 1987;
        ELSIF x = 7141 THEN
            sigmoid_f := 1987;
        ELSIF x = 7142 THEN
            sigmoid_f := 1987;
        ELSIF x = 7143 THEN
            sigmoid_f := 1987;
        ELSIF x = 7144 THEN
            sigmoid_f := 1987;
        ELSIF x = 7145 THEN
            sigmoid_f := 1987;
        ELSIF x = 7146 THEN
            sigmoid_f := 1987;
        ELSIF x = 7147 THEN
            sigmoid_f := 1987;
        ELSIF x = 7148 THEN
            sigmoid_f := 1987;
        ELSIF x = 7149 THEN
            sigmoid_f := 1987;
        ELSIF x = 7150 THEN
            sigmoid_f := 1987;
        ELSIF x = 7151 THEN
            sigmoid_f := 1987;
        ELSIF x = 7152 THEN
            sigmoid_f := 1987;
        ELSIF x = 7153 THEN
            sigmoid_f := 1987;
        ELSIF x = 7154 THEN
            sigmoid_f := 1987;
        ELSIF x = 7155 THEN
            sigmoid_f := 1987;
        ELSIF x = 7156 THEN
            sigmoid_f := 1987;
        ELSIF x = 7157 THEN
            sigmoid_f := 1987;
        ELSIF x = 7158 THEN
            sigmoid_f := 1987;
        ELSIF x = 7159 THEN
            sigmoid_f := 1987;
        ELSIF x = 7160 THEN
            sigmoid_f := 1987;
        ELSIF x = 7161 THEN
            sigmoid_f := 1987;
        ELSIF x = 7162 THEN
            sigmoid_f := 1987;
        ELSIF x = 7163 THEN
            sigmoid_f := 1987;
        ELSIF x = 7164 THEN
            sigmoid_f := 1987;
        ELSIF x = 7165 THEN
            sigmoid_f := 1987;
        ELSIF x = 7166 THEN
            sigmoid_f := 1987;
        ELSIF x = 7167 THEN
            sigmoid_f := 1987;
        ELSIF x = 7168 THEN
            sigmoid_f := 1988;
        ELSIF x = 7169 THEN
            sigmoid_f := 1988;
        ELSIF x = 7170 THEN
            sigmoid_f := 1988;
        ELSIF x = 7171 THEN
            sigmoid_f := 1988;
        ELSIF x = 7172 THEN
            sigmoid_f := 1988;
        ELSIF x = 7173 THEN
            sigmoid_f := 1988;
        ELSIF x = 7174 THEN
            sigmoid_f := 1988;
        ELSIF x = 7175 THEN
            sigmoid_f := 1988;
        ELSIF x = 7176 THEN
            sigmoid_f := 1988;
        ELSIF x = 7177 THEN
            sigmoid_f := 1988;
        ELSIF x = 7178 THEN
            sigmoid_f := 1988;
        ELSIF x = 7179 THEN
            sigmoid_f := 1988;
        ELSIF x = 7180 THEN
            sigmoid_f := 1988;
        ELSIF x = 7181 THEN
            sigmoid_f := 1988;
        ELSIF x = 7182 THEN
            sigmoid_f := 1988;
        ELSIF x = 7183 THEN
            sigmoid_f := 1988;
        ELSIF x = 7184 THEN
            sigmoid_f := 1988;
        ELSIF x = 7185 THEN
            sigmoid_f := 1988;
        ELSIF x = 7186 THEN
            sigmoid_f := 1988;
        ELSIF x = 7187 THEN
            sigmoid_f := 1988;
        ELSIF x = 7188 THEN
            sigmoid_f := 1988;
        ELSIF x = 7189 THEN
            sigmoid_f := 1988;
        ELSIF x = 7190 THEN
            sigmoid_f := 1988;
        ELSIF x = 7191 THEN
            sigmoid_f := 1988;
        ELSIF x = 7192 THEN
            sigmoid_f := 1988;
        ELSIF x = 7193 THEN
            sigmoid_f := 1988;
        ELSIF x = 7194 THEN
            sigmoid_f := 1988;
        ELSIF x = 7195 THEN
            sigmoid_f := 1988;
        ELSIF x = 7196 THEN
            sigmoid_f := 1988;
        ELSIF x = 7197 THEN
            sigmoid_f := 1988;
        ELSIF x = 7198 THEN
            sigmoid_f := 1988;
        ELSIF x = 7199 THEN
            sigmoid_f := 1988;
        ELSIF x = 7200 THEN
            sigmoid_f := 1988;
        ELSIF x = 7201 THEN
            sigmoid_f := 1988;
        ELSIF x = 7202 THEN
            sigmoid_f := 1988;
        ELSIF x = 7203 THEN
            sigmoid_f := 1988;
        ELSIF x = 7204 THEN
            sigmoid_f := 1988;
        ELSIF x = 7205 THEN
            sigmoid_f := 1988;
        ELSIF x = 7206 THEN
            sigmoid_f := 1989;
        ELSIF x = 7207 THEN
            sigmoid_f := 1989;
        ELSIF x = 7208 THEN
            sigmoid_f := 1989;
        ELSIF x = 7209 THEN
            sigmoid_f := 1989;
        ELSIF x = 7210 THEN
            sigmoid_f := 1989;
        ELSIF x = 7211 THEN
            sigmoid_f := 1989;
        ELSIF x = 7212 THEN
            sigmoid_f := 1989;
        ELSIF x = 7213 THEN
            sigmoid_f := 1989;
        ELSIF x = 7214 THEN
            sigmoid_f := 1989;
        ELSIF x = 7215 THEN
            sigmoid_f := 1989;
        ELSIF x = 7216 THEN
            sigmoid_f := 1989;
        ELSIF x = 7217 THEN
            sigmoid_f := 1989;
        ELSIF x = 7218 THEN
            sigmoid_f := 1989;
        ELSIF x = 7219 THEN
            sigmoid_f := 1989;
        ELSIF x = 7220 THEN
            sigmoid_f := 1989;
        ELSIF x = 7221 THEN
            sigmoid_f := 1989;
        ELSIF x = 7222 THEN
            sigmoid_f := 1989;
        ELSIF x = 7223 THEN
            sigmoid_f := 1989;
        ELSIF x = 7224 THEN
            sigmoid_f := 1989;
        ELSIF x = 7225 THEN
            sigmoid_f := 1989;
        ELSIF x = 7226 THEN
            sigmoid_f := 1989;
        ELSIF x = 7227 THEN
            sigmoid_f := 1989;
        ELSIF x = 7228 THEN
            sigmoid_f := 1989;
        ELSIF x = 7229 THEN
            sigmoid_f := 1989;
        ELSIF x = 7230 THEN
            sigmoid_f := 1989;
        ELSIF x = 7231 THEN
            sigmoid_f := 1989;
        ELSIF x = 7232 THEN
            sigmoid_f := 1989;
        ELSIF x = 7233 THEN
            sigmoid_f := 1989;
        ELSIF x = 7234 THEN
            sigmoid_f := 1989;
        ELSIF x = 7235 THEN
            sigmoid_f := 1989;
        ELSIF x = 7236 THEN
            sigmoid_f := 1989;
        ELSIF x = 7237 THEN
            sigmoid_f := 1989;
        ELSIF x = 7238 THEN
            sigmoid_f := 1989;
        ELSIF x = 7239 THEN
            sigmoid_f := 1989;
        ELSIF x = 7240 THEN
            sigmoid_f := 1989;
        ELSIF x = 7241 THEN
            sigmoid_f := 1989;
        ELSIF x = 7242 THEN
            sigmoid_f := 1989;
        ELSIF x = 7243 THEN
            sigmoid_f := 1989;
        ELSIF x = 7244 THEN
            sigmoid_f := 1990;
        ELSIF x = 7245 THEN
            sigmoid_f := 1990;
        ELSIF x = 7246 THEN
            sigmoid_f := 1990;
        ELSIF x = 7247 THEN
            sigmoid_f := 1990;
        ELSIF x = 7248 THEN
            sigmoid_f := 1990;
        ELSIF x = 7249 THEN
            sigmoid_f := 1990;
        ELSIF x = 7250 THEN
            sigmoid_f := 1990;
        ELSIF x = 7251 THEN
            sigmoid_f := 1990;
        ELSIF x = 7252 THEN
            sigmoid_f := 1990;
        ELSIF x = 7253 THEN
            sigmoid_f := 1990;
        ELSIF x = 7254 THEN
            sigmoid_f := 1990;
        ELSIF x = 7255 THEN
            sigmoid_f := 1990;
        ELSIF x = 7256 THEN
            sigmoid_f := 1990;
        ELSIF x = 7257 THEN
            sigmoid_f := 1990;
        ELSIF x = 7258 THEN
            sigmoid_f := 1990;
        ELSIF x = 7259 THEN
            sigmoid_f := 1990;
        ELSIF x = 7260 THEN
            sigmoid_f := 1990;
        ELSIF x = 7261 THEN
            sigmoid_f := 1990;
        ELSIF x = 7262 THEN
            sigmoid_f := 1990;
        ELSIF x = 7263 THEN
            sigmoid_f := 1990;
        ELSIF x = 7264 THEN
            sigmoid_f := 1990;
        ELSIF x = 7265 THEN
            sigmoid_f := 1990;
        ELSIF x = 7266 THEN
            sigmoid_f := 1990;
        ELSIF x = 7267 THEN
            sigmoid_f := 1990;
        ELSIF x = 7268 THEN
            sigmoid_f := 1990;
        ELSIF x = 7269 THEN
            sigmoid_f := 1990;
        ELSIF x = 7270 THEN
            sigmoid_f := 1990;
        ELSIF x = 7271 THEN
            sigmoid_f := 1990;
        ELSIF x = 7272 THEN
            sigmoid_f := 1990;
        ELSIF x = 7273 THEN
            sigmoid_f := 1990;
        ELSIF x = 7274 THEN
            sigmoid_f := 1990;
        ELSIF x = 7275 THEN
            sigmoid_f := 1990;
        ELSIF x = 7276 THEN
            sigmoid_f := 1990;
        ELSIF x = 7277 THEN
            sigmoid_f := 1990;
        ELSIF x = 7278 THEN
            sigmoid_f := 1990;
        ELSIF x = 7279 THEN
            sigmoid_f := 1990;
        ELSIF x = 7280 THEN
            sigmoid_f := 1990;
        ELSIF x = 7281 THEN
            sigmoid_f := 1990;
        ELSIF x = 7282 THEN
            sigmoid_f := 1991;
        ELSIF x = 7283 THEN
            sigmoid_f := 1991;
        ELSIF x = 7284 THEN
            sigmoid_f := 1991;
        ELSIF x = 7285 THEN
            sigmoid_f := 1991;
        ELSIF x = 7286 THEN
            sigmoid_f := 1991;
        ELSIF x = 7287 THEN
            sigmoid_f := 1991;
        ELSIF x = 7288 THEN
            sigmoid_f := 1991;
        ELSIF x = 7289 THEN
            sigmoid_f := 1991;
        ELSIF x = 7290 THEN
            sigmoid_f := 1991;
        ELSIF x = 7291 THEN
            sigmoid_f := 1991;
        ELSIF x = 7292 THEN
            sigmoid_f := 1991;
        ELSIF x = 7293 THEN
            sigmoid_f := 1991;
        ELSIF x = 7294 THEN
            sigmoid_f := 1991;
        ELSIF x = 7295 THEN
            sigmoid_f := 1991;
        ELSIF x = 7296 THEN
            sigmoid_f := 1991;
        ELSIF x = 7297 THEN
            sigmoid_f := 1991;
        ELSIF x = 7298 THEN
            sigmoid_f := 1991;
        ELSIF x = 7299 THEN
            sigmoid_f := 1991;
        ELSIF x = 7300 THEN
            sigmoid_f := 1991;
        ELSIF x = 7301 THEN
            sigmoid_f := 1991;
        ELSIF x = 7302 THEN
            sigmoid_f := 1991;
        ELSIF x = 7303 THEN
            sigmoid_f := 1991;
        ELSIF x = 7304 THEN
            sigmoid_f := 1991;
        ELSIF x = 7305 THEN
            sigmoid_f := 1991;
        ELSIF x = 7306 THEN
            sigmoid_f := 1991;
        ELSIF x = 7307 THEN
            sigmoid_f := 1991;
        ELSIF x = 7308 THEN
            sigmoid_f := 1991;
        ELSIF x = 7309 THEN
            sigmoid_f := 1991;
        ELSIF x = 7310 THEN
            sigmoid_f := 1991;
        ELSIF x = 7311 THEN
            sigmoid_f := 1991;
        ELSIF x = 7312 THEN
            sigmoid_f := 1991;
        ELSIF x = 7313 THEN
            sigmoid_f := 1991;
        ELSIF x = 7314 THEN
            sigmoid_f := 1991;
        ELSIF x = 7315 THEN
            sigmoid_f := 1991;
        ELSIF x = 7316 THEN
            sigmoid_f := 1991;
        ELSIF x = 7317 THEN
            sigmoid_f := 1991;
        ELSIF x = 7318 THEN
            sigmoid_f := 1991;
        ELSIF x = 7319 THEN
            sigmoid_f := 1991;
        ELSIF x = 7320 THEN
            sigmoid_f := 1992;
        ELSIF x = 7321 THEN
            sigmoid_f := 1992;
        ELSIF x = 7322 THEN
            sigmoid_f := 1992;
        ELSIF x = 7323 THEN
            sigmoid_f := 1992;
        ELSIF x = 7324 THEN
            sigmoid_f := 1992;
        ELSIF x = 7325 THEN
            sigmoid_f := 1992;
        ELSIF x = 7326 THEN
            sigmoid_f := 1992;
        ELSIF x = 7327 THEN
            sigmoid_f := 1992;
        ELSIF x = 7328 THEN
            sigmoid_f := 1992;
        ELSIF x = 7329 THEN
            sigmoid_f := 1992;
        ELSIF x = 7330 THEN
            sigmoid_f := 1992;
        ELSIF x = 7331 THEN
            sigmoid_f := 1992;
        ELSIF x = 7332 THEN
            sigmoid_f := 1992;
        ELSIF x = 7333 THEN
            sigmoid_f := 1992;
        ELSIF x = 7334 THEN
            sigmoid_f := 1992;
        ELSIF x = 7335 THEN
            sigmoid_f := 1992;
        ELSIF x = 7336 THEN
            sigmoid_f := 1992;
        ELSIF x = 7337 THEN
            sigmoid_f := 1992;
        ELSIF x = 7338 THEN
            sigmoid_f := 1992;
        ELSIF x = 7339 THEN
            sigmoid_f := 1992;
        ELSIF x = 7340 THEN
            sigmoid_f := 1992;
        ELSIF x = 7341 THEN
            sigmoid_f := 1992;
        ELSIF x = 7342 THEN
            sigmoid_f := 1992;
        ELSIF x = 7343 THEN
            sigmoid_f := 1992;
        ELSIF x = 7344 THEN
            sigmoid_f := 1992;
        ELSIF x = 7345 THEN
            sigmoid_f := 1992;
        ELSIF x = 7346 THEN
            sigmoid_f := 1992;
        ELSIF x = 7347 THEN
            sigmoid_f := 1992;
        ELSIF x = 7348 THEN
            sigmoid_f := 1992;
        ELSIF x = 7349 THEN
            sigmoid_f := 1992;
        ELSIF x = 7350 THEN
            sigmoid_f := 1992;
        ELSIF x = 7351 THEN
            sigmoid_f := 1992;
        ELSIF x = 7352 THEN
            sigmoid_f := 1992;
        ELSIF x = 7353 THEN
            sigmoid_f := 1992;
        ELSIF x = 7354 THEN
            sigmoid_f := 1992;
        ELSIF x = 7355 THEN
            sigmoid_f := 1992;
        ELSIF x = 7356 THEN
            sigmoid_f := 1992;
        ELSIF x = 7357 THEN
            sigmoid_f := 1992;
        ELSIF x = 7358 THEN
            sigmoid_f := 1993;
        ELSIF x = 7359 THEN
            sigmoid_f := 1993;
        ELSIF x = 7360 THEN
            sigmoid_f := 1993;
        ELSIF x = 7361 THEN
            sigmoid_f := 1993;
        ELSIF x = 7362 THEN
            sigmoid_f := 1993;
        ELSIF x = 7363 THEN
            sigmoid_f := 1993;
        ELSIF x = 7364 THEN
            sigmoid_f := 1993;
        ELSIF x = 7365 THEN
            sigmoid_f := 1993;
        ELSIF x = 7366 THEN
            sigmoid_f := 1993;
        ELSIF x = 7367 THEN
            sigmoid_f := 1993;
        ELSIF x = 7368 THEN
            sigmoid_f := 1993;
        ELSIF x = 7369 THEN
            sigmoid_f := 1993;
        ELSIF x = 7370 THEN
            sigmoid_f := 1993;
        ELSIF x = 7371 THEN
            sigmoid_f := 1993;
        ELSIF x = 7372 THEN
            sigmoid_f := 1993;
        ELSIF x = 7373 THEN
            sigmoid_f := 1993;
        ELSIF x = 7374 THEN
            sigmoid_f := 1993;
        ELSIF x = 7375 THEN
            sigmoid_f := 1993;
        ELSIF x = 7376 THEN
            sigmoid_f := 1993;
        ELSIF x = 7377 THEN
            sigmoid_f := 1993;
        ELSIF x = 7378 THEN
            sigmoid_f := 1993;
        ELSIF x = 7379 THEN
            sigmoid_f := 1993;
        ELSIF x = 7380 THEN
            sigmoid_f := 1993;
        ELSIF x = 7381 THEN
            sigmoid_f := 1993;
        ELSIF x = 7382 THEN
            sigmoid_f := 1993;
        ELSIF x = 7383 THEN
            sigmoid_f := 1993;
        ELSIF x = 7384 THEN
            sigmoid_f := 1993;
        ELSIF x = 7385 THEN
            sigmoid_f := 1993;
        ELSIF x = 7386 THEN
            sigmoid_f := 1993;
        ELSIF x = 7387 THEN
            sigmoid_f := 1993;
        ELSIF x = 7388 THEN
            sigmoid_f := 1993;
        ELSIF x = 7389 THEN
            sigmoid_f := 1993;
        ELSIF x = 7390 THEN
            sigmoid_f := 1993;
        ELSIF x = 7391 THEN
            sigmoid_f := 1993;
        ELSIF x = 7392 THEN
            sigmoid_f := 1993;
        ELSIF x = 7393 THEN
            sigmoid_f := 1993;
        ELSIF x = 7394 THEN
            sigmoid_f := 1993;
        ELSIF x = 7395 THEN
            sigmoid_f := 1993;
        ELSIF x = 7396 THEN
            sigmoid_f := 1994;
        ELSIF x = 7397 THEN
            sigmoid_f := 1994;
        ELSIF x = 7398 THEN
            sigmoid_f := 1994;
        ELSIF x = 7399 THEN
            sigmoid_f := 1994;
        ELSIF x = 7400 THEN
            sigmoid_f := 1994;
        ELSIF x = 7401 THEN
            sigmoid_f := 1994;
        ELSIF x = 7402 THEN
            sigmoid_f := 1994;
        ELSIF x = 7403 THEN
            sigmoid_f := 1994;
        ELSIF x = 7404 THEN
            sigmoid_f := 1994;
        ELSIF x = 7405 THEN
            sigmoid_f := 1994;
        ELSIF x = 7406 THEN
            sigmoid_f := 1994;
        ELSIF x = 7407 THEN
            sigmoid_f := 1994;
        ELSIF x = 7408 THEN
            sigmoid_f := 1994;
        ELSIF x = 7409 THEN
            sigmoid_f := 1994;
        ELSIF x = 7410 THEN
            sigmoid_f := 1994;
        ELSIF x = 7411 THEN
            sigmoid_f := 1994;
        ELSIF x = 7412 THEN
            sigmoid_f := 1994;
        ELSIF x = 7413 THEN
            sigmoid_f := 1994;
        ELSIF x = 7414 THEN
            sigmoid_f := 1994;
        ELSIF x = 7415 THEN
            sigmoid_f := 1994;
        ELSIF x = 7416 THEN
            sigmoid_f := 1994;
        ELSIF x = 7417 THEN
            sigmoid_f := 1994;
        ELSIF x = 7418 THEN
            sigmoid_f := 1994;
        ELSIF x = 7419 THEN
            sigmoid_f := 1994;
        ELSIF x = 7420 THEN
            sigmoid_f := 1994;
        ELSIF x = 7421 THEN
            sigmoid_f := 1994;
        ELSIF x = 7422 THEN
            sigmoid_f := 1994;
        ELSIF x = 7423 THEN
            sigmoid_f := 1994;
        ELSIF x = 7424 THEN
            sigmoid_f := 1994;
        ELSIF x = 7425 THEN
            sigmoid_f := 1994;
        ELSIF x = 7426 THEN
            sigmoid_f := 1994;
        ELSIF x = 7427 THEN
            sigmoid_f := 1994;
        ELSIF x = 7428 THEN
            sigmoid_f := 1994;
        ELSIF x = 7429 THEN
            sigmoid_f := 1994;
        ELSIF x = 7430 THEN
            sigmoid_f := 1994;
        ELSIF x = 7431 THEN
            sigmoid_f := 1994;
        ELSIF x = 7432 THEN
            sigmoid_f := 1994;
        ELSIF x = 7433 THEN
            sigmoid_f := 1994;
        ELSIF x = 7434 THEN
            sigmoid_f := 1995;
        ELSIF x = 7435 THEN
            sigmoid_f := 1995;
        ELSIF x = 7436 THEN
            sigmoid_f := 1995;
        ELSIF x = 7437 THEN
            sigmoid_f := 1995;
        ELSIF x = 7438 THEN
            sigmoid_f := 1995;
        ELSIF x = 7439 THEN
            sigmoid_f := 1995;
        ELSIF x = 7440 THEN
            sigmoid_f := 1995;
        ELSIF x = 7441 THEN
            sigmoid_f := 1995;
        ELSIF x = 7442 THEN
            sigmoid_f := 1995;
        ELSIF x = 7443 THEN
            sigmoid_f := 1995;
        ELSIF x = 7444 THEN
            sigmoid_f := 1995;
        ELSIF x = 7445 THEN
            sigmoid_f := 1995;
        ELSIF x = 7446 THEN
            sigmoid_f := 1995;
        ELSIF x = 7447 THEN
            sigmoid_f := 1995;
        ELSIF x = 7448 THEN
            sigmoid_f := 1995;
        ELSIF x = 7449 THEN
            sigmoid_f := 1995;
        ELSIF x = 7450 THEN
            sigmoid_f := 1995;
        ELSIF x = 7451 THEN
            sigmoid_f := 1995;
        ELSIF x = 7452 THEN
            sigmoid_f := 1995;
        ELSIF x = 7453 THEN
            sigmoid_f := 1995;
        ELSIF x = 7454 THEN
            sigmoid_f := 1995;
        ELSIF x = 7455 THEN
            sigmoid_f := 1995;
        ELSIF x = 7456 THEN
            sigmoid_f := 1995;
        ELSIF x = 7457 THEN
            sigmoid_f := 1995;
        ELSIF x = 7458 THEN
            sigmoid_f := 1995;
        ELSIF x = 7459 THEN
            sigmoid_f := 1995;
        ELSIF x = 7460 THEN
            sigmoid_f := 1995;
        ELSIF x = 7461 THEN
            sigmoid_f := 1995;
        ELSIF x = 7462 THEN
            sigmoid_f := 1995;
        ELSIF x = 7463 THEN
            sigmoid_f := 1995;
        ELSIF x = 7464 THEN
            sigmoid_f := 1995;
        ELSIF x = 7465 THEN
            sigmoid_f := 1995;
        ELSIF x = 7466 THEN
            sigmoid_f := 1995;
        ELSIF x = 7467 THEN
            sigmoid_f := 1995;
        ELSIF x = 7468 THEN
            sigmoid_f := 1995;
        ELSIF x = 7469 THEN
            sigmoid_f := 1995;
        ELSIF x = 7470 THEN
            sigmoid_f := 1995;
        ELSIF x = 7471 THEN
            sigmoid_f := 1995;
        ELSIF x = 7472 THEN
            sigmoid_f := 1996;
        ELSIF x = 7473 THEN
            sigmoid_f := 1996;
        ELSIF x = 7474 THEN
            sigmoid_f := 1996;
        ELSIF x = 7475 THEN
            sigmoid_f := 1996;
        ELSIF x = 7476 THEN
            sigmoid_f := 1996;
        ELSIF x = 7477 THEN
            sigmoid_f := 1996;
        ELSIF x = 7478 THEN
            sigmoid_f := 1996;
        ELSIF x = 7479 THEN
            sigmoid_f := 1996;
        ELSIF x = 7480 THEN
            sigmoid_f := 1996;
        ELSIF x = 7481 THEN
            sigmoid_f := 1996;
        ELSIF x = 7482 THEN
            sigmoid_f := 1996;
        ELSIF x = 7483 THEN
            sigmoid_f := 1996;
        ELSIF x = 7484 THEN
            sigmoid_f := 1996;
        ELSIF x = 7485 THEN
            sigmoid_f := 1996;
        ELSIF x = 7486 THEN
            sigmoid_f := 1996;
        ELSIF x = 7487 THEN
            sigmoid_f := 1996;
        ELSIF x = 7488 THEN
            sigmoid_f := 1996;
        ELSIF x = 7489 THEN
            sigmoid_f := 1996;
        ELSIF x = 7490 THEN
            sigmoid_f := 1996;
        ELSIF x = 7491 THEN
            sigmoid_f := 1996;
        ELSIF x = 7492 THEN
            sigmoid_f := 1996;
        ELSIF x = 7493 THEN
            sigmoid_f := 1996;
        ELSIF x = 7494 THEN
            sigmoid_f := 1996;
        ELSIF x = 7495 THEN
            sigmoid_f := 1996;
        ELSIF x = 7496 THEN
            sigmoid_f := 1996;
        ELSIF x = 7497 THEN
            sigmoid_f := 1996;
        ELSIF x = 7498 THEN
            sigmoid_f := 1996;
        ELSIF x = 7499 THEN
            sigmoid_f := 1996;
        ELSIF x = 7500 THEN
            sigmoid_f := 1996;
        ELSIF x = 7501 THEN
            sigmoid_f := 1996;
        ELSIF x = 7502 THEN
            sigmoid_f := 1996;
        ELSIF x = 7503 THEN
            sigmoid_f := 1996;
        ELSIF x = 7504 THEN
            sigmoid_f := 1996;
        ELSIF x = 7505 THEN
            sigmoid_f := 1996;
        ELSIF x = 7506 THEN
            sigmoid_f := 1996;
        ELSIF x = 7507 THEN
            sigmoid_f := 1996;
        ELSIF x = 7508 THEN
            sigmoid_f := 1996;
        ELSIF x = 7509 THEN
            sigmoid_f := 1996;
        ELSIF x = 7510 THEN
            sigmoid_f := 1997;
        ELSIF x = 7511 THEN
            sigmoid_f := 1997;
        ELSIF x = 7512 THEN
            sigmoid_f := 1997;
        ELSIF x = 7513 THEN
            sigmoid_f := 1997;
        ELSIF x = 7514 THEN
            sigmoid_f := 1997;
        ELSIF x = 7515 THEN
            sigmoid_f := 1997;
        ELSIF x = 7516 THEN
            sigmoid_f := 1997;
        ELSIF x = 7517 THEN
            sigmoid_f := 1997;
        ELSIF x = 7518 THEN
            sigmoid_f := 1997;
        ELSIF x = 7519 THEN
            sigmoid_f := 1997;
        ELSIF x = 7520 THEN
            sigmoid_f := 1997;
        ELSIF x = 7521 THEN
            sigmoid_f := 1997;
        ELSIF x = 7522 THEN
            sigmoid_f := 1997;
        ELSIF x = 7523 THEN
            sigmoid_f := 1997;
        ELSIF x = 7524 THEN
            sigmoid_f := 1997;
        ELSIF x = 7525 THEN
            sigmoid_f := 1997;
        ELSIF x = 7526 THEN
            sigmoid_f := 1997;
        ELSIF x = 7527 THEN
            sigmoid_f := 1997;
        ELSIF x = 7528 THEN
            sigmoid_f := 1997;
        ELSIF x = 7529 THEN
            sigmoid_f := 1997;
        ELSIF x = 7530 THEN
            sigmoid_f := 1997;
        ELSIF x = 7531 THEN
            sigmoid_f := 1997;
        ELSIF x = 7532 THEN
            sigmoid_f := 1997;
        ELSIF x = 7533 THEN
            sigmoid_f := 1997;
        ELSIF x = 7534 THEN
            sigmoid_f := 1997;
        ELSIF x = 7535 THEN
            sigmoid_f := 1997;
        ELSIF x = 7536 THEN
            sigmoid_f := 1997;
        ELSIF x = 7537 THEN
            sigmoid_f := 1997;
        ELSIF x = 7538 THEN
            sigmoid_f := 1997;
        ELSIF x = 7539 THEN
            sigmoid_f := 1997;
        ELSIF x = 7540 THEN
            sigmoid_f := 1997;
        ELSIF x = 7541 THEN
            sigmoid_f := 1997;
        ELSIF x = 7542 THEN
            sigmoid_f := 1997;
        ELSIF x = 7543 THEN
            sigmoid_f := 1997;
        ELSIF x = 7544 THEN
            sigmoid_f := 1997;
        ELSIF x = 7545 THEN
            sigmoid_f := 1997;
        ELSIF x = 7546 THEN
            sigmoid_f := 1997;
        ELSIF x = 7547 THEN
            sigmoid_f := 1997;
        ELSIF x = 7548 THEN
            sigmoid_f := 1998;
        ELSIF x = 7549 THEN
            sigmoid_f := 1998;
        ELSIF x = 7550 THEN
            sigmoid_f := 1998;
        ELSIF x = 7551 THEN
            sigmoid_f := 1998;
        ELSIF x = 7552 THEN
            sigmoid_f := 1998;
        ELSIF x = 7553 THEN
            sigmoid_f := 1998;
        ELSIF x = 7554 THEN
            sigmoid_f := 1998;
        ELSIF x = 7555 THEN
            sigmoid_f := 1998;
        ELSIF x = 7556 THEN
            sigmoid_f := 1998;
        ELSIF x = 7557 THEN
            sigmoid_f := 1998;
        ELSIF x = 7558 THEN
            sigmoid_f := 1998;
        ELSIF x = 7559 THEN
            sigmoid_f := 1998;
        ELSIF x = 7560 THEN
            sigmoid_f := 1998;
        ELSIF x = 7561 THEN
            sigmoid_f := 1998;
        ELSIF x = 7562 THEN
            sigmoid_f := 1998;
        ELSIF x = 7563 THEN
            sigmoid_f := 1998;
        ELSIF x = 7564 THEN
            sigmoid_f := 1998;
        ELSIF x = 7565 THEN
            sigmoid_f := 1998;
        ELSIF x = 7566 THEN
            sigmoid_f := 1998;
        ELSIF x = 7567 THEN
            sigmoid_f := 1998;
        ELSIF x = 7568 THEN
            sigmoid_f := 1998;
        ELSIF x = 7569 THEN
            sigmoid_f := 1998;
        ELSIF x = 7570 THEN
            sigmoid_f := 1998;
        ELSIF x = 7571 THEN
            sigmoid_f := 1998;
        ELSIF x = 7572 THEN
            sigmoid_f := 1998;
        ELSIF x = 7573 THEN
            sigmoid_f := 1998;
        ELSIF x = 7574 THEN
            sigmoid_f := 1998;
        ELSIF x = 7575 THEN
            sigmoid_f := 1998;
        ELSIF x = 7576 THEN
            sigmoid_f := 1998;
        ELSIF x = 7577 THEN
            sigmoid_f := 1998;
        ELSIF x = 7578 THEN
            sigmoid_f := 1998;
        ELSIF x = 7579 THEN
            sigmoid_f := 1998;
        ELSIF x = 7580 THEN
            sigmoid_f := 1998;
        ELSIF x = 7581 THEN
            sigmoid_f := 1998;
        ELSIF x = 7582 THEN
            sigmoid_f := 1998;
        ELSIF x = 7583 THEN
            sigmoid_f := 1998;
        ELSIF x = 7584 THEN
            sigmoid_f := 1998;
        ELSIF x = 7585 THEN
            sigmoid_f := 1998;
        ELSIF x = 7586 THEN
            sigmoid_f := 1999;
        ELSIF x = 7587 THEN
            sigmoid_f := 1999;
        ELSIF x = 7588 THEN
            sigmoid_f := 1999;
        ELSIF x = 7589 THEN
            sigmoid_f := 1999;
        ELSIF x = 7590 THEN
            sigmoid_f := 1999;
        ELSIF x = 7591 THEN
            sigmoid_f := 1999;
        ELSIF x = 7592 THEN
            sigmoid_f := 1999;
        ELSIF x = 7593 THEN
            sigmoid_f := 1999;
        ELSIF x = 7594 THEN
            sigmoid_f := 1999;
        ELSIF x = 7595 THEN
            sigmoid_f := 1999;
        ELSIF x = 7596 THEN
            sigmoid_f := 1999;
        ELSIF x = 7597 THEN
            sigmoid_f := 1999;
        ELSIF x = 7598 THEN
            sigmoid_f := 1999;
        ELSIF x = 7599 THEN
            sigmoid_f := 1999;
        ELSIF x = 7600 THEN
            sigmoid_f := 1999;
        ELSIF x = 7601 THEN
            sigmoid_f := 1999;
        ELSIF x = 7602 THEN
            sigmoid_f := 1999;
        ELSIF x = 7603 THEN
            sigmoid_f := 1999;
        ELSIF x = 7604 THEN
            sigmoid_f := 1999;
        ELSIF x = 7605 THEN
            sigmoid_f := 1999;
        ELSIF x = 7606 THEN
            sigmoid_f := 1999;
        ELSIF x = 7607 THEN
            sigmoid_f := 1999;
        ELSIF x = 7608 THEN
            sigmoid_f := 1999;
        ELSIF x = 7609 THEN
            sigmoid_f := 1999;
        ELSIF x = 7610 THEN
            sigmoid_f := 1999;
        ELSIF x = 7611 THEN
            sigmoid_f := 1999;
        ELSIF x = 7612 THEN
            sigmoid_f := 1999;
        ELSIF x = 7613 THEN
            sigmoid_f := 1999;
        ELSIF x = 7614 THEN
            sigmoid_f := 1999;
        ELSIF x = 7615 THEN
            sigmoid_f := 1999;
        ELSIF x = 7616 THEN
            sigmoid_f := 1999;
        ELSIF x = 7617 THEN
            sigmoid_f := 1999;
        ELSIF x = 7618 THEN
            sigmoid_f := 1999;
        ELSIF x = 7619 THEN
            sigmoid_f := 1999;
        ELSIF x = 7620 THEN
            sigmoid_f := 1999;
        ELSIF x = 7621 THEN
            sigmoid_f := 1999;
        ELSIF x = 7622 THEN
            sigmoid_f := 1999;
        ELSIF x = 7623 THEN
            sigmoid_f := 1999;
        ELSIF x = 7624 THEN
            sigmoid_f := 2000;
        ELSIF x = 7625 THEN
            sigmoid_f := 2000;
        ELSIF x = 7626 THEN
            sigmoid_f := 2000;
        ELSIF x = 7627 THEN
            sigmoid_f := 2000;
        ELSIF x = 7628 THEN
            sigmoid_f := 2000;
        ELSIF x = 7629 THEN
            sigmoid_f := 2000;
        ELSIF x = 7630 THEN
            sigmoid_f := 2000;
        ELSIF x = 7631 THEN
            sigmoid_f := 2000;
        ELSIF x = 7632 THEN
            sigmoid_f := 2000;
        ELSIF x = 7633 THEN
            sigmoid_f := 2000;
        ELSIF x = 7634 THEN
            sigmoid_f := 2000;
        ELSIF x = 7635 THEN
            sigmoid_f := 2000;
        ELSIF x = 7636 THEN
            sigmoid_f := 2000;
        ELSIF x = 7637 THEN
            sigmoid_f := 2000;
        ELSIF x = 7638 THEN
            sigmoid_f := 2000;
        ELSIF x = 7639 THEN
            sigmoid_f := 2000;
        ELSIF x = 7640 THEN
            sigmoid_f := 2000;
        ELSIF x = 7641 THEN
            sigmoid_f := 2000;
        ELSIF x = 7642 THEN
            sigmoid_f := 2000;
        ELSIF x = 7643 THEN
            sigmoid_f := 2000;
        ELSIF x = 7644 THEN
            sigmoid_f := 2000;
        ELSIF x = 7645 THEN
            sigmoid_f := 2000;
        ELSIF x = 7646 THEN
            sigmoid_f := 2000;
        ELSIF x = 7647 THEN
            sigmoid_f := 2000;
        ELSIF x = 7648 THEN
            sigmoid_f := 2000;
        ELSIF x = 7649 THEN
            sigmoid_f := 2000;
        ELSIF x = 7650 THEN
            sigmoid_f := 2000;
        ELSIF x = 7651 THEN
            sigmoid_f := 2000;
        ELSIF x = 7652 THEN
            sigmoid_f := 2000;
        ELSIF x = 7653 THEN
            sigmoid_f := 2000;
        ELSIF x = 7654 THEN
            sigmoid_f := 2000;
        ELSIF x = 7655 THEN
            sigmoid_f := 2000;
        ELSIF x = 7656 THEN
            sigmoid_f := 2000;
        ELSIF x = 7657 THEN
            sigmoid_f := 2000;
        ELSIF x = 7658 THEN
            sigmoid_f := 2000;
        ELSIF x = 7659 THEN
            sigmoid_f := 2000;
        ELSIF x = 7660 THEN
            sigmoid_f := 2000;
        ELSIF x = 7661 THEN
            sigmoid_f := 2000;
        ELSIF x = 7662 THEN
            sigmoid_f := 2001;
        ELSIF x = 7663 THEN
            sigmoid_f := 2001;
        ELSIF x = 7664 THEN
            sigmoid_f := 2001;
        ELSIF x = 7665 THEN
            sigmoid_f := 2001;
        ELSIF x = 7666 THEN
            sigmoid_f := 2001;
        ELSIF x = 7667 THEN
            sigmoid_f := 2001;
        ELSIF x = 7668 THEN
            sigmoid_f := 2001;
        ELSIF x = 7669 THEN
            sigmoid_f := 2001;
        ELSIF x = 7670 THEN
            sigmoid_f := 2001;
        ELSIF x = 7671 THEN
            sigmoid_f := 2001;
        ELSIF x = 7672 THEN
            sigmoid_f := 2001;
        ELSIF x = 7673 THEN
            sigmoid_f := 2001;
        ELSIF x = 7674 THEN
            sigmoid_f := 2001;
        ELSIF x = 7675 THEN
            sigmoid_f := 2001;
        ELSIF x = 7676 THEN
            sigmoid_f := 2001;
        ELSIF x = 7677 THEN
            sigmoid_f := 2001;
        ELSIF x = 7678 THEN
            sigmoid_f := 2001;
        ELSIF x = 7679 THEN
            sigmoid_f := 2001;
        ELSIF x = 7680 THEN
            sigmoid_f := 2001;
        ELSIF x = 7681 THEN
            sigmoid_f := 2001;
        ELSIF x = 7682 THEN
            sigmoid_f := 2001;
        ELSIF x = 7683 THEN
            sigmoid_f := 2001;
        ELSIF x = 7684 THEN
            sigmoid_f := 2001;
        ELSIF x = 7685 THEN
            sigmoid_f := 2001;
        ELSIF x = 7686 THEN
            sigmoid_f := 2001;
        ELSIF x = 7687 THEN
            sigmoid_f := 2001;
        ELSIF x = 7688 THEN
            sigmoid_f := 2001;
        ELSIF x = 7689 THEN
            sigmoid_f := 2001;
        ELSIF x = 7690 THEN
            sigmoid_f := 2001;
        ELSIF x = 7691 THEN
            sigmoid_f := 2001;
        ELSIF x = 7692 THEN
            sigmoid_f := 2001;
        ELSIF x = 7693 THEN
            sigmoid_f := 2001;
        ELSIF x = 7694 THEN
            sigmoid_f := 2001;
        ELSIF x = 7695 THEN
            sigmoid_f := 2001;
        ELSIF x = 7696 THEN
            sigmoid_f := 2001;
        ELSIF x = 7697 THEN
            sigmoid_f := 2001;
        ELSIF x = 7698 THEN
            sigmoid_f := 2001;
        ELSIF x = 7699 THEN
            sigmoid_f := 2001;
        ELSIF x = 7700 THEN
            sigmoid_f := 2001;
        ELSIF x = 7701 THEN
            sigmoid_f := 2001;
        ELSIF x = 7702 THEN
            sigmoid_f := 2001;
        ELSIF x = 7703 THEN
            sigmoid_f := 2001;
        ELSIF x = 7704 THEN
            sigmoid_f := 2001;
        ELSIF x = 7705 THEN
            sigmoid_f := 2001;
        ELSIF x = 7706 THEN
            sigmoid_f := 2001;
        ELSIF x = 7707 THEN
            sigmoid_f := 2001;
        ELSIF x = 7708 THEN
            sigmoid_f := 2001;
        ELSIF x = 7709 THEN
            sigmoid_f := 2001;
        ELSIF x = 7710 THEN
            sigmoid_f := 2001;
        ELSIF x = 7711 THEN
            sigmoid_f := 2001;
        ELSIF x = 7712 THEN
            sigmoid_f := 2001;
        ELSIF x = 7713 THEN
            sigmoid_f := 2001;
        ELSIF x = 7714 THEN
            sigmoid_f := 2001;
        ELSIF x = 7715 THEN
            sigmoid_f := 2001;
        ELSIF x = 7716 THEN
            sigmoid_f := 2001;
        ELSIF x = 7717 THEN
            sigmoid_f := 2001;
        ELSIF x = 7718 THEN
            sigmoid_f := 2001;
        ELSIF x = 7719 THEN
            sigmoid_f := 2001;
        ELSIF x = 7720 THEN
            sigmoid_f := 2002;
        ELSIF x = 7721 THEN
            sigmoid_f := 2002;
        ELSIF x = 7722 THEN
            sigmoid_f := 2002;
        ELSIF x = 7723 THEN
            sigmoid_f := 2002;
        ELSIF x = 7724 THEN
            sigmoid_f := 2002;
        ELSIF x = 7725 THEN
            sigmoid_f := 2002;
        ELSIF x = 7726 THEN
            sigmoid_f := 2002;
        ELSIF x = 7727 THEN
            sigmoid_f := 2002;
        ELSIF x = 7728 THEN
            sigmoid_f := 2002;
        ELSIF x = 7729 THEN
            sigmoid_f := 2002;
        ELSIF x = 7730 THEN
            sigmoid_f := 2002;
        ELSIF x = 7731 THEN
            sigmoid_f := 2002;
        ELSIF x = 7732 THEN
            sigmoid_f := 2002;
        ELSIF x = 7733 THEN
            sigmoid_f := 2002;
        ELSIF x = 7734 THEN
            sigmoid_f := 2002;
        ELSIF x = 7735 THEN
            sigmoid_f := 2002;
        ELSIF x = 7736 THEN
            sigmoid_f := 2002;
        ELSIF x = 7737 THEN
            sigmoid_f := 2002;
        ELSIF x = 7738 THEN
            sigmoid_f := 2002;
        ELSIF x = 7739 THEN
            sigmoid_f := 2002;
        ELSIF x = 7740 THEN
            sigmoid_f := 2002;
        ELSIF x = 7741 THEN
            sigmoid_f := 2002;
        ELSIF x = 7742 THEN
            sigmoid_f := 2002;
        ELSIF x = 7743 THEN
            sigmoid_f := 2002;
        ELSIF x = 7744 THEN
            sigmoid_f := 2002;
        ELSIF x = 7745 THEN
            sigmoid_f := 2002;
        ELSIF x = 7746 THEN
            sigmoid_f := 2002;
        ELSIF x = 7747 THEN
            sigmoid_f := 2002;
        ELSIF x = 7748 THEN
            sigmoid_f := 2002;
        ELSIF x = 7749 THEN
            sigmoid_f := 2002;
        ELSIF x = 7750 THEN
            sigmoid_f := 2002;
        ELSIF x = 7751 THEN
            sigmoid_f := 2002;
        ELSIF x = 7752 THEN
            sigmoid_f := 2002;
        ELSIF x = 7753 THEN
            sigmoid_f := 2002;
        ELSIF x = 7754 THEN
            sigmoid_f := 2002;
        ELSIF x = 7755 THEN
            sigmoid_f := 2002;
        ELSIF x = 7756 THEN
            sigmoid_f := 2002;
        ELSIF x = 7757 THEN
            sigmoid_f := 2002;
        ELSIF x = 7758 THEN
            sigmoid_f := 2002;
        ELSIF x = 7759 THEN
            sigmoid_f := 2002;
        ELSIF x = 7760 THEN
            sigmoid_f := 2002;
        ELSIF x = 7761 THEN
            sigmoid_f := 2002;
        ELSIF x = 7762 THEN
            sigmoid_f := 2002;
        ELSIF x = 7763 THEN
            sigmoid_f := 2002;
        ELSIF x = 7764 THEN
            sigmoid_f := 2002;
        ELSIF x = 7765 THEN
            sigmoid_f := 2002;
        ELSIF x = 7766 THEN
            sigmoid_f := 2002;
        ELSIF x = 7767 THEN
            sigmoid_f := 2002;
        ELSIF x = 7768 THEN
            sigmoid_f := 2002;
        ELSIF x = 7769 THEN
            sigmoid_f := 2002;
        ELSIF x = 7770 THEN
            sigmoid_f := 2002;
        ELSIF x = 7771 THEN
            sigmoid_f := 2002;
        ELSIF x = 7772 THEN
            sigmoid_f := 2003;
        ELSIF x = 7773 THEN
            sigmoid_f := 2003;
        ELSIF x = 7774 THEN
            sigmoid_f := 2003;
        ELSIF x = 7775 THEN
            sigmoid_f := 2003;
        ELSIF x = 7776 THEN
            sigmoid_f := 2003;
        ELSIF x = 7777 THEN
            sigmoid_f := 2003;
        ELSIF x = 7778 THEN
            sigmoid_f := 2003;
        ELSIF x = 7779 THEN
            sigmoid_f := 2003;
        ELSIF x = 7780 THEN
            sigmoid_f := 2003;
        ELSIF x = 7781 THEN
            sigmoid_f := 2003;
        ELSIF x = 7782 THEN
            sigmoid_f := 2003;
        ELSIF x = 7783 THEN
            sigmoid_f := 2003;
        ELSIF x = 7784 THEN
            sigmoid_f := 2003;
        ELSIF x = 7785 THEN
            sigmoid_f := 2003;
        ELSIF x = 7786 THEN
            sigmoid_f := 2003;
        ELSIF x = 7787 THEN
            sigmoid_f := 2003;
        ELSIF x = 7788 THEN
            sigmoid_f := 2003;
        ELSIF x = 7789 THEN
            sigmoid_f := 2003;
        ELSIF x = 7790 THEN
            sigmoid_f := 2003;
        ELSIF x = 7791 THEN
            sigmoid_f := 2003;
        ELSIF x = 7792 THEN
            sigmoid_f := 2003;
        ELSIF x = 7793 THEN
            sigmoid_f := 2003;
        ELSIF x = 7794 THEN
            sigmoid_f := 2003;
        ELSIF x = 7795 THEN
            sigmoid_f := 2003;
        ELSIF x = 7796 THEN
            sigmoid_f := 2003;
        ELSIF x = 7797 THEN
            sigmoid_f := 2003;
        ELSIF x = 7798 THEN
            sigmoid_f := 2003;
        ELSIF x = 7799 THEN
            sigmoid_f := 2003;
        ELSIF x = 7800 THEN
            sigmoid_f := 2003;
        ELSIF x = 7801 THEN
            sigmoid_f := 2003;
        ELSIF x = 7802 THEN
            sigmoid_f := 2003;
        ELSIF x = 7803 THEN
            sigmoid_f := 2003;
        ELSIF x = 7804 THEN
            sigmoid_f := 2003;
        ELSIF x = 7805 THEN
            sigmoid_f := 2003;
        ELSIF x = 7806 THEN
            sigmoid_f := 2003;
        ELSIF x = 7807 THEN
            sigmoid_f := 2003;
        ELSIF x = 7808 THEN
            sigmoid_f := 2003;
        ELSIF x = 7809 THEN
            sigmoid_f := 2003;
        ELSIF x = 7810 THEN
            sigmoid_f := 2003;
        ELSIF x = 7811 THEN
            sigmoid_f := 2003;
        ELSIF x = 7812 THEN
            sigmoid_f := 2003;
        ELSIF x = 7813 THEN
            sigmoid_f := 2003;
        ELSIF x = 7814 THEN
            sigmoid_f := 2003;
        ELSIF x = 7815 THEN
            sigmoid_f := 2003;
        ELSIF x = 7816 THEN
            sigmoid_f := 2003;
        ELSIF x = 7817 THEN
            sigmoid_f := 2003;
        ELSIF x = 7818 THEN
            sigmoid_f := 2003;
        ELSIF x = 7819 THEN
            sigmoid_f := 2003;
        ELSIF x = 7820 THEN
            sigmoid_f := 2003;
        ELSIF x = 7821 THEN
            sigmoid_f := 2003;
        ELSIF x = 7822 THEN
            sigmoid_f := 2003;
        ELSIF x = 7823 THEN
            sigmoid_f := 2003;
        ELSIF x = 7824 THEN
            sigmoid_f := 2003;
        ELSIF x = 7825 THEN
            sigmoid_f := 2004;
        ELSIF x = 7826 THEN
            sigmoid_f := 2004;
        ELSIF x = 7827 THEN
            sigmoid_f := 2004;
        ELSIF x = 7828 THEN
            sigmoid_f := 2004;
        ELSIF x = 7829 THEN
            sigmoid_f := 2004;
        ELSIF x = 7830 THEN
            sigmoid_f := 2004;
        ELSIF x = 7831 THEN
            sigmoid_f := 2004;
        ELSIF x = 7832 THEN
            sigmoid_f := 2004;
        ELSIF x = 7833 THEN
            sigmoid_f := 2004;
        ELSIF x = 7834 THEN
            sigmoid_f := 2004;
        ELSIF x = 7835 THEN
            sigmoid_f := 2004;
        ELSIF x = 7836 THEN
            sigmoid_f := 2004;
        ELSIF x = 7837 THEN
            sigmoid_f := 2004;
        ELSIF x = 7838 THEN
            sigmoid_f := 2004;
        ELSIF x = 7839 THEN
            sigmoid_f := 2004;
        ELSIF x = 7840 THEN
            sigmoid_f := 2004;
        ELSIF x = 7841 THEN
            sigmoid_f := 2004;
        ELSIF x = 7842 THEN
            sigmoid_f := 2004;
        ELSIF x = 7843 THEN
            sigmoid_f := 2004;
        ELSIF x = 7844 THEN
            sigmoid_f := 2004;
        ELSIF x = 7845 THEN
            sigmoid_f := 2004;
        ELSIF x = 7846 THEN
            sigmoid_f := 2004;
        ELSIF x = 7847 THEN
            sigmoid_f := 2004;
        ELSIF x = 7848 THEN
            sigmoid_f := 2004;
        ELSIF x = 7849 THEN
            sigmoid_f := 2004;
        ELSIF x = 7850 THEN
            sigmoid_f := 2004;
        ELSIF x = 7851 THEN
            sigmoid_f := 2004;
        ELSIF x = 7852 THEN
            sigmoid_f := 2004;
        ELSIF x = 7853 THEN
            sigmoid_f := 2004;
        ELSIF x = 7854 THEN
            sigmoid_f := 2004;
        ELSIF x = 7855 THEN
            sigmoid_f := 2004;
        ELSIF x = 7856 THEN
            sigmoid_f := 2004;
        ELSIF x = 7857 THEN
            sigmoid_f := 2004;
        ELSIF x = 7858 THEN
            sigmoid_f := 2004;
        ELSIF x = 7859 THEN
            sigmoid_f := 2004;
        ELSIF x = 7860 THEN
            sigmoid_f := 2004;
        ELSIF x = 7861 THEN
            sigmoid_f := 2004;
        ELSIF x = 7862 THEN
            sigmoid_f := 2004;
        ELSIF x = 7863 THEN
            sigmoid_f := 2004;
        ELSIF x = 7864 THEN
            sigmoid_f := 2004;
        ELSIF x = 7865 THEN
            sigmoid_f := 2004;
        ELSIF x = 7866 THEN
            sigmoid_f := 2004;
        ELSIF x = 7867 THEN
            sigmoid_f := 2004;
        ELSIF x = 7868 THEN
            sigmoid_f := 2004;
        ELSIF x = 7869 THEN
            sigmoid_f := 2004;
        ELSIF x = 7870 THEN
            sigmoid_f := 2004;
        ELSIF x = 7871 THEN
            sigmoid_f := 2004;
        ELSIF x = 7872 THEN
            sigmoid_f := 2004;
        ELSIF x = 7873 THEN
            sigmoid_f := 2004;
        ELSIF x = 7874 THEN
            sigmoid_f := 2004;
        ELSIF x = 7875 THEN
            sigmoid_f := 2004;
        ELSIF x = 7876 THEN
            sigmoid_f := 2004;
        ELSIF x = 7877 THEN
            sigmoid_f := 2005;
        ELSIF x = 7878 THEN
            sigmoid_f := 2005;
        ELSIF x = 7879 THEN
            sigmoid_f := 2005;
        ELSIF x = 7880 THEN
            sigmoid_f := 2005;
        ELSIF x = 7881 THEN
            sigmoid_f := 2005;
        ELSIF x = 7882 THEN
            sigmoid_f := 2005;
        ELSIF x = 7883 THEN
            sigmoid_f := 2005;
        ELSIF x = 7884 THEN
            sigmoid_f := 2005;
        ELSIF x = 7885 THEN
            sigmoid_f := 2005;
        ELSIF x = 7886 THEN
            sigmoid_f := 2005;
        ELSIF x = 7887 THEN
            sigmoid_f := 2005;
        ELSIF x = 7888 THEN
            sigmoid_f := 2005;
        ELSIF x = 7889 THEN
            sigmoid_f := 2005;
        ELSIF x = 7890 THEN
            sigmoid_f := 2005;
        ELSIF x = 7891 THEN
            sigmoid_f := 2005;
        ELSIF x = 7892 THEN
            sigmoid_f := 2005;
        ELSIF x = 7893 THEN
            sigmoid_f := 2005;
        ELSIF x = 7894 THEN
            sigmoid_f := 2005;
        ELSIF x = 7895 THEN
            sigmoid_f := 2005;
        ELSIF x = 7896 THEN
            sigmoid_f := 2005;
        ELSIF x = 7897 THEN
            sigmoid_f := 2005;
        ELSIF x = 7898 THEN
            sigmoid_f := 2005;
        ELSIF x = 7899 THEN
            sigmoid_f := 2005;
        ELSIF x = 7900 THEN
            sigmoid_f := 2005;
        ELSIF x = 7901 THEN
            sigmoid_f := 2005;
        ELSIF x = 7902 THEN
            sigmoid_f := 2005;
        ELSIF x = 7903 THEN
            sigmoid_f := 2005;
        ELSIF x = 7904 THEN
            sigmoid_f := 2005;
        ELSIF x = 7905 THEN
            sigmoid_f := 2005;
        ELSIF x = 7906 THEN
            sigmoid_f := 2005;
        ELSIF x = 7907 THEN
            sigmoid_f := 2005;
        ELSIF x = 7908 THEN
            sigmoid_f := 2005;
        ELSIF x = 7909 THEN
            sigmoid_f := 2005;
        ELSIF x = 7910 THEN
            sigmoid_f := 2005;
        ELSIF x = 7911 THEN
            sigmoid_f := 2005;
        ELSIF x = 7912 THEN
            sigmoid_f := 2005;
        ELSIF x = 7913 THEN
            sigmoid_f := 2005;
        ELSIF x = 7914 THEN
            sigmoid_f := 2005;
        ELSIF x = 7915 THEN
            sigmoid_f := 2005;
        ELSIF x = 7916 THEN
            sigmoid_f := 2005;
        ELSIF x = 7917 THEN
            sigmoid_f := 2005;
        ELSIF x = 7918 THEN
            sigmoid_f := 2005;
        ELSIF x = 7919 THEN
            sigmoid_f := 2005;
        ELSIF x = 7920 THEN
            sigmoid_f := 2005;
        ELSIF x = 7921 THEN
            sigmoid_f := 2005;
        ELSIF x = 7922 THEN
            sigmoid_f := 2005;
        ELSIF x = 7923 THEN
            sigmoid_f := 2005;
        ELSIF x = 7924 THEN
            sigmoid_f := 2005;
        ELSIF x = 7925 THEN
            sigmoid_f := 2005;
        ELSIF x = 7926 THEN
            sigmoid_f := 2005;
        ELSIF x = 7927 THEN
            sigmoid_f := 2005;
        ELSIF x = 7928 THEN
            sigmoid_f := 2005;
        ELSIF x = 7929 THEN
            sigmoid_f := 2005;
        ELSIF x = 7930 THEN
            sigmoid_f := 2006;
        ELSIF x = 7931 THEN
            sigmoid_f := 2006;
        ELSIF x = 7932 THEN
            sigmoid_f := 2006;
        ELSIF x = 7933 THEN
            sigmoid_f := 2006;
        ELSIF x = 7934 THEN
            sigmoid_f := 2006;
        ELSIF x = 7935 THEN
            sigmoid_f := 2006;
        ELSIF x = 7936 THEN
            sigmoid_f := 2006;
        ELSIF x = 7937 THEN
            sigmoid_f := 2006;
        ELSIF x = 7938 THEN
            sigmoid_f := 2006;
        ELSIF x = 7939 THEN
            sigmoid_f := 2006;
        ELSIF x = 7940 THEN
            sigmoid_f := 2006;
        ELSIF x = 7941 THEN
            sigmoid_f := 2006;
        ELSIF x = 7942 THEN
            sigmoid_f := 2006;
        ELSIF x = 7943 THEN
            sigmoid_f := 2006;
        ELSIF x = 7944 THEN
            sigmoid_f := 2006;
        ELSIF x = 7945 THEN
            sigmoid_f := 2006;
        ELSIF x = 7946 THEN
            sigmoid_f := 2006;
        ELSIF x = 7947 THEN
            sigmoid_f := 2006;
        ELSIF x = 7948 THEN
            sigmoid_f := 2006;
        ELSIF x = 7949 THEN
            sigmoid_f := 2006;
        ELSIF x = 7950 THEN
            sigmoid_f := 2006;
        ELSIF x = 7951 THEN
            sigmoid_f := 2006;
        ELSIF x = 7952 THEN
            sigmoid_f := 2006;
        ELSIF x = 7953 THEN
            sigmoid_f := 2006;
        ELSIF x = 7954 THEN
            sigmoid_f := 2006;
        ELSIF x = 7955 THEN
            sigmoid_f := 2006;
        ELSIF x = 7956 THEN
            sigmoid_f := 2006;
        ELSIF x = 7957 THEN
            sigmoid_f := 2006;
        ELSIF x = 7958 THEN
            sigmoid_f := 2006;
        ELSIF x = 7959 THEN
            sigmoid_f := 2006;
        ELSIF x = 7960 THEN
            sigmoid_f := 2006;
        ELSIF x = 7961 THEN
            sigmoid_f := 2006;
        ELSIF x = 7962 THEN
            sigmoid_f := 2006;
        ELSIF x = 7963 THEN
            sigmoid_f := 2006;
        ELSIF x = 7964 THEN
            sigmoid_f := 2006;
        ELSIF x = 7965 THEN
            sigmoid_f := 2006;
        ELSIF x = 7966 THEN
            sigmoid_f := 2006;
        ELSIF x = 7967 THEN
            sigmoid_f := 2006;
        ELSIF x = 7968 THEN
            sigmoid_f := 2006;
        ELSIF x = 7969 THEN
            sigmoid_f := 2006;
        ELSIF x = 7970 THEN
            sigmoid_f := 2006;
        ELSIF x = 7971 THEN
            sigmoid_f := 2006;
        ELSIF x = 7972 THEN
            sigmoid_f := 2006;
        ELSIF x = 7973 THEN
            sigmoid_f := 2006;
        ELSIF x = 7974 THEN
            sigmoid_f := 2006;
        ELSIF x = 7975 THEN
            sigmoid_f := 2006;
        ELSIF x = 7976 THEN
            sigmoid_f := 2006;
        ELSIF x = 7977 THEN
            sigmoid_f := 2006;
        ELSIF x = 7978 THEN
            sigmoid_f := 2006;
        ELSIF x = 7979 THEN
            sigmoid_f := 2006;
        ELSIF x = 7980 THEN
            sigmoid_f := 2006;
        ELSIF x = 7981 THEN
            sigmoid_f := 2006;
        ELSIF x = 7982 THEN
            sigmoid_f := 2007;
        ELSIF x = 7983 THEN
            sigmoid_f := 2007;
        ELSIF x = 7984 THEN
            sigmoid_f := 2007;
        ELSIF x = 7985 THEN
            sigmoid_f := 2007;
        ELSIF x = 7986 THEN
            sigmoid_f := 2007;
        ELSIF x = 7987 THEN
            sigmoid_f := 2007;
        ELSIF x = 7988 THEN
            sigmoid_f := 2007;
        ELSIF x = 7989 THEN
            sigmoid_f := 2007;
        ELSIF x = 7990 THEN
            sigmoid_f := 2007;
        ELSIF x = 7991 THEN
            sigmoid_f := 2007;
        ELSIF x = 7992 THEN
            sigmoid_f := 2007;
        ELSIF x = 7993 THEN
            sigmoid_f := 2007;
        ELSIF x = 7994 THEN
            sigmoid_f := 2007;
        ELSIF x = 7995 THEN
            sigmoid_f := 2007;
        ELSIF x = 7996 THEN
            sigmoid_f := 2007;
        ELSIF x = 7997 THEN
            sigmoid_f := 2007;
        ELSIF x = 7998 THEN
            sigmoid_f := 2007;
        ELSIF x = 7999 THEN
            sigmoid_f := 2007;
        ELSIF x = 8000 THEN
            sigmoid_f := 2007;
        ELSIF x = 8001 THEN
            sigmoid_f := 2007;
        ELSIF x = 8002 THEN
            sigmoid_f := 2007;
        ELSIF x = 8003 THEN
            sigmoid_f := 2007;
        ELSIF x = 8004 THEN
            sigmoid_f := 2007;
        ELSIF x = 8005 THEN
            sigmoid_f := 2007;
        ELSIF x = 8006 THEN
            sigmoid_f := 2007;
        ELSIF x = 8007 THEN
            sigmoid_f := 2007;
        ELSIF x = 8008 THEN
            sigmoid_f := 2007;
        ELSIF x = 8009 THEN
            sigmoid_f := 2007;
        ELSIF x = 8010 THEN
            sigmoid_f := 2007;
        ELSIF x = 8011 THEN
            sigmoid_f := 2007;
        ELSIF x = 8012 THEN
            sigmoid_f := 2007;
        ELSIF x = 8013 THEN
            sigmoid_f := 2007;
        ELSIF x = 8014 THEN
            sigmoid_f := 2007;
        ELSIF x = 8015 THEN
            sigmoid_f := 2007;
        ELSIF x = 8016 THEN
            sigmoid_f := 2007;
        ELSIF x = 8017 THEN
            sigmoid_f := 2007;
        ELSIF x = 8018 THEN
            sigmoid_f := 2007;
        ELSIF x = 8019 THEN
            sigmoid_f := 2007;
        ELSIF x = 8020 THEN
            sigmoid_f := 2007;
        ELSIF x = 8021 THEN
            sigmoid_f := 2007;
        ELSIF x = 8022 THEN
            sigmoid_f := 2007;
        ELSIF x = 8023 THEN
            sigmoid_f := 2007;
        ELSIF x = 8024 THEN
            sigmoid_f := 2007;
        ELSIF x = 8025 THEN
            sigmoid_f := 2007;
        ELSIF x = 8026 THEN
            sigmoid_f := 2007;
        ELSIF x = 8027 THEN
            sigmoid_f := 2007;
        ELSIF x = 8028 THEN
            sigmoid_f := 2007;
        ELSIF x = 8029 THEN
            sigmoid_f := 2007;
        ELSIF x = 8030 THEN
            sigmoid_f := 2007;
        ELSIF x = 8031 THEN
            sigmoid_f := 2007;
        ELSIF x = 8032 THEN
            sigmoid_f := 2007;
        ELSIF x = 8033 THEN
            sigmoid_f := 2007;
        ELSIF x = 8034 THEN
            sigmoid_f := 2007;
        ELSIF x = 8035 THEN
            sigmoid_f := 2008;
        ELSIF x = 8036 THEN
            sigmoid_f := 2008;
        ELSIF x = 8037 THEN
            sigmoid_f := 2008;
        ELSIF x = 8038 THEN
            sigmoid_f := 2008;
        ELSIF x = 8039 THEN
            sigmoid_f := 2008;
        ELSIF x = 8040 THEN
            sigmoid_f := 2008;
        ELSIF x = 8041 THEN
            sigmoid_f := 2008;
        ELSIF x = 8042 THEN
            sigmoid_f := 2008;
        ELSIF x = 8043 THEN
            sigmoid_f := 2008;
        ELSIF x = 8044 THEN
            sigmoid_f := 2008;
        ELSIF x = 8045 THEN
            sigmoid_f := 2008;
        ELSIF x = 8046 THEN
            sigmoid_f := 2008;
        ELSIF x = 8047 THEN
            sigmoid_f := 2008;
        ELSIF x = 8048 THEN
            sigmoid_f := 2008;
        ELSIF x = 8049 THEN
            sigmoid_f := 2008;
        ELSIF x = 8050 THEN
            sigmoid_f := 2008;
        ELSIF x = 8051 THEN
            sigmoid_f := 2008;
        ELSIF x = 8052 THEN
            sigmoid_f := 2008;
        ELSIF x = 8053 THEN
            sigmoid_f := 2008;
        ELSIF x = 8054 THEN
            sigmoid_f := 2008;
        ELSIF x = 8055 THEN
            sigmoid_f := 2008;
        ELSIF x = 8056 THEN
            sigmoid_f := 2008;
        ELSIF x = 8057 THEN
            sigmoid_f := 2008;
        ELSIF x = 8058 THEN
            sigmoid_f := 2008;
        ELSIF x = 8059 THEN
            sigmoid_f := 2008;
        ELSIF x = 8060 THEN
            sigmoid_f := 2008;
        ELSIF x = 8061 THEN
            sigmoid_f := 2008;
        ELSIF x = 8062 THEN
            sigmoid_f := 2008;
        ELSIF x = 8063 THEN
            sigmoid_f := 2008;
        ELSIF x = 8064 THEN
            sigmoid_f := 2008;
        ELSIF x = 8065 THEN
            sigmoid_f := 2008;
        ELSIF x = 8066 THEN
            sigmoid_f := 2008;
        ELSIF x = 8067 THEN
            sigmoid_f := 2008;
        ELSIF x = 8068 THEN
            sigmoid_f := 2008;
        ELSIF x = 8069 THEN
            sigmoid_f := 2008;
        ELSIF x = 8070 THEN
            sigmoid_f := 2008;
        ELSIF x = 8071 THEN
            sigmoid_f := 2008;
        ELSIF x = 8072 THEN
            sigmoid_f := 2008;
        ELSIF x = 8073 THEN
            sigmoid_f := 2008;
        ELSIF x = 8074 THEN
            sigmoid_f := 2008;
        ELSIF x = 8075 THEN
            sigmoid_f := 2008;
        ELSIF x = 8076 THEN
            sigmoid_f := 2008;
        ELSIF x = 8077 THEN
            sigmoid_f := 2008;
        ELSIF x = 8078 THEN
            sigmoid_f := 2008;
        ELSIF x = 8079 THEN
            sigmoid_f := 2008;
        ELSIF x = 8080 THEN
            sigmoid_f := 2008;
        ELSIF x = 8081 THEN
            sigmoid_f := 2008;
        ELSIF x = 8082 THEN
            sigmoid_f := 2008;
        ELSIF x = 8083 THEN
            sigmoid_f := 2008;
        ELSIF x = 8084 THEN
            sigmoid_f := 2008;
        ELSIF x = 8085 THEN
            sigmoid_f := 2008;
        ELSIF x = 8086 THEN
            sigmoid_f := 2008;
        ELSIF x = 8087 THEN
            sigmoid_f := 2009;
        ELSIF x = 8088 THEN
            sigmoid_f := 2009;
        ELSIF x = 8089 THEN
            sigmoid_f := 2009;
        ELSIF x = 8090 THEN
            sigmoid_f := 2009;
        ELSIF x = 8091 THEN
            sigmoid_f := 2009;
        ELSIF x = 8092 THEN
            sigmoid_f := 2009;
        ELSIF x = 8093 THEN
            sigmoid_f := 2009;
        ELSIF x = 8094 THEN
            sigmoid_f := 2009;
        ELSIF x = 8095 THEN
            sigmoid_f := 2009;
        ELSIF x = 8096 THEN
            sigmoid_f := 2009;
        ELSIF x = 8097 THEN
            sigmoid_f := 2009;
        ELSIF x = 8098 THEN
            sigmoid_f := 2009;
        ELSIF x = 8099 THEN
            sigmoid_f := 2009;
        ELSIF x = 8100 THEN
            sigmoid_f := 2009;
        ELSIF x = 8101 THEN
            sigmoid_f := 2009;
        ELSIF x = 8102 THEN
            sigmoid_f := 2009;
        ELSIF x = 8103 THEN
            sigmoid_f := 2009;
        ELSIF x = 8104 THEN
            sigmoid_f := 2009;
        ELSIF x = 8105 THEN
            sigmoid_f := 2009;
        ELSIF x = 8106 THEN
            sigmoid_f := 2009;
        ELSIF x = 8107 THEN
            sigmoid_f := 2009;
        ELSIF x = 8108 THEN
            sigmoid_f := 2009;
        ELSIF x = 8109 THEN
            sigmoid_f := 2009;
        ELSIF x = 8110 THEN
            sigmoid_f := 2009;
        ELSIF x = 8111 THEN
            sigmoid_f := 2009;
        ELSIF x = 8112 THEN
            sigmoid_f := 2009;
        ELSIF x = 8113 THEN
            sigmoid_f := 2009;
        ELSIF x = 8114 THEN
            sigmoid_f := 2009;
        ELSIF x = 8115 THEN
            sigmoid_f := 2009;
        ELSIF x = 8116 THEN
            sigmoid_f := 2009;
        ELSIF x = 8117 THEN
            sigmoid_f := 2009;
        ELSIF x = 8118 THEN
            sigmoid_f := 2009;
        ELSIF x = 8119 THEN
            sigmoid_f := 2009;
        ELSIF x = 8120 THEN
            sigmoid_f := 2009;
        ELSIF x = 8121 THEN
            sigmoid_f := 2009;
        ELSIF x = 8122 THEN
            sigmoid_f := 2009;
        ELSIF x = 8123 THEN
            sigmoid_f := 2009;
        ELSIF x = 8124 THEN
            sigmoid_f := 2009;
        ELSIF x = 8125 THEN
            sigmoid_f := 2009;
        ELSIF x = 8126 THEN
            sigmoid_f := 2009;
        ELSIF x = 8127 THEN
            sigmoid_f := 2009;
        ELSIF x = 8128 THEN
            sigmoid_f := 2009;
        ELSIF x = 8129 THEN
            sigmoid_f := 2009;
        ELSIF x = 8130 THEN
            sigmoid_f := 2009;
        ELSIF x = 8131 THEN
            sigmoid_f := 2009;
        ELSIF x = 8132 THEN
            sigmoid_f := 2009;
        ELSIF x = 8133 THEN
            sigmoid_f := 2009;
        ELSIF x = 8134 THEN
            sigmoid_f := 2009;
        ELSIF x = 8135 THEN
            sigmoid_f := 2009;
        ELSIF x = 8136 THEN
            sigmoid_f := 2009;
        ELSIF x = 8137 THEN
            sigmoid_f := 2009;
        ELSIF x = 8138 THEN
            sigmoid_f := 2009;
        ELSIF x = 8139 THEN
            sigmoid_f := 2009;
        ELSIF x = 8140 THEN
            sigmoid_f := 2010;
        ELSIF x = 8141 THEN
            sigmoid_f := 2010;
        ELSIF x = 8142 THEN
            sigmoid_f := 2010;
        ELSIF x = 8143 THEN
            sigmoid_f := 2010;
        ELSIF x = 8144 THEN
            sigmoid_f := 2010;
        ELSIF x = 8145 THEN
            sigmoid_f := 2010;
        ELSIF x = 8146 THEN
            sigmoid_f := 2010;
        ELSIF x = 8147 THEN
            sigmoid_f := 2010;
        ELSIF x = 8148 THEN
            sigmoid_f := 2010;
        ELSIF x = 8149 THEN
            sigmoid_f := 2010;
        ELSIF x = 8150 THEN
            sigmoid_f := 2010;
        ELSIF x = 8151 THEN
            sigmoid_f := 2010;
        ELSIF x = 8152 THEN
            sigmoid_f := 2010;
        ELSIF x = 8153 THEN
            sigmoid_f := 2010;
        ELSIF x = 8154 THEN
            sigmoid_f := 2010;
        ELSIF x = 8155 THEN
            sigmoid_f := 2010;
        ELSIF x = 8156 THEN
            sigmoid_f := 2010;
        ELSIF x = 8157 THEN
            sigmoid_f := 2010;
        ELSIF x = 8158 THEN
            sigmoid_f := 2010;
        ELSIF x = 8159 THEN
            sigmoid_f := 2010;
        ELSIF x = 8160 THEN
            sigmoid_f := 2010;
        ELSIF x = 8161 THEN
            sigmoid_f := 2010;
        ELSIF x = 8162 THEN
            sigmoid_f := 2010;
        ELSIF x = 8163 THEN
            sigmoid_f := 2010;
        ELSIF x = 8164 THEN
            sigmoid_f := 2010;
        ELSIF x = 8165 THEN
            sigmoid_f := 2010;
        ELSIF x = 8166 THEN
            sigmoid_f := 2010;
        ELSIF x = 8167 THEN
            sigmoid_f := 2010;
        ELSIF x = 8168 THEN
            sigmoid_f := 2010;
        ELSIF x = 8169 THEN
            sigmoid_f := 2010;
        ELSIF x = 8170 THEN
            sigmoid_f := 2010;
        ELSIF x = 8171 THEN
            sigmoid_f := 2010;
        ELSIF x = 8172 THEN
            sigmoid_f := 2010;
        ELSIF x = 8173 THEN
            sigmoid_f := 2010;
        ELSIF x = 8174 THEN
            sigmoid_f := 2010;
        ELSIF x = 8175 THEN
            sigmoid_f := 2010;
        ELSIF x = 8176 THEN
            sigmoid_f := 2010;
        ELSIF x = 8177 THEN
            sigmoid_f := 2010;
        ELSIF x = 8178 THEN
            sigmoid_f := 2010;
        ELSIF x = 8179 THEN
            sigmoid_f := 2010;
        ELSIF x = 8180 THEN
            sigmoid_f := 2010;
        ELSIF x = 8181 THEN
            sigmoid_f := 2010;
        ELSIF x = 8182 THEN
            sigmoid_f := 2010;
        ELSIF x = 8183 THEN
            sigmoid_f := 2010;
        ELSIF x = 8184 THEN
            sigmoid_f := 2010;
        ELSIF x = 8185 THEN
            sigmoid_f := 2010;
        ELSIF x = 8186 THEN
            sigmoid_f := 2010;
        ELSIF x = 8187 THEN
            sigmoid_f := 2010;
        ELSIF x = 8188 THEN
            sigmoid_f := 2010;
        ELSIF x = 8189 THEN
            sigmoid_f := 2010;
        ELSIF x = 8190 THEN
            sigmoid_f := 2010;
        ELSIF x = 8191 THEN
            sigmoid_f := 2010;
        ELSIF x = 8192 THEN
            sigmoid_f := 2011;
        ELSIF x = 8193 THEN
            sigmoid_f := 2011;
        ELSIF x = 8194 THEN
            sigmoid_f := 2011;
        ELSIF x = 8195 THEN
            sigmoid_f := 2011;
        ELSIF x = 8196 THEN
            sigmoid_f := 2011;
        ELSIF x = 8197 THEN
            sigmoid_f := 2011;
        ELSIF x = 8198 THEN
            sigmoid_f := 2011;
        ELSIF x = 8199 THEN
            sigmoid_f := 2011;
        ELSIF x = 8200 THEN
            sigmoid_f := 2011;
        ELSIF x = 8201 THEN
            sigmoid_f := 2011;
        ELSIF x = 8202 THEN
            sigmoid_f := 2011;
        ELSIF x = 8203 THEN
            sigmoid_f := 2011;
        ELSIF x = 8204 THEN
            sigmoid_f := 2011;
        ELSIF x = 8205 THEN
            sigmoid_f := 2011;
        ELSIF x = 8206 THEN
            sigmoid_f := 2011;
        ELSIF x = 8207 THEN
            sigmoid_f := 2011;
        ELSIF x = 8208 THEN
            sigmoid_f := 2011;
        ELSIF x = 8209 THEN
            sigmoid_f := 2011;
        ELSIF x = 8210 THEN
            sigmoid_f := 2011;
        ELSIF x = 8211 THEN
            sigmoid_f := 2011;
        ELSIF x = 8212 THEN
            sigmoid_f := 2011;
        ELSIF x = 8213 THEN
            sigmoid_f := 2011;
        ELSIF x = 8214 THEN
            sigmoid_f := 2011;
        ELSIF x = 8215 THEN
            sigmoid_f := 2011;
        ELSIF x = 8216 THEN
            sigmoid_f := 2011;
        ELSIF x = 8217 THEN
            sigmoid_f := 2011;
        ELSIF x = 8218 THEN
            sigmoid_f := 2011;
        ELSIF x = 8219 THEN
            sigmoid_f := 2011;
        ELSIF x = 8220 THEN
            sigmoid_f := 2011;
        ELSIF x = 8221 THEN
            sigmoid_f := 2011;
        ELSIF x = 8222 THEN
            sigmoid_f := 2011;
        ELSIF x = 8223 THEN
            sigmoid_f := 2011;
        ELSIF x = 8224 THEN
            sigmoid_f := 2011;
        ELSIF x = 8225 THEN
            sigmoid_f := 2011;
        ELSIF x = 8226 THEN
            sigmoid_f := 2011;
        ELSIF x = 8227 THEN
            sigmoid_f := 2011;
        ELSIF x = 8228 THEN
            sigmoid_f := 2011;
        ELSIF x = 8229 THEN
            sigmoid_f := 2011;
        ELSIF x = 8230 THEN
            sigmoid_f := 2011;
        ELSIF x = 8231 THEN
            sigmoid_f := 2011;
        ELSIF x = 8232 THEN
            sigmoid_f := 2011;
        ELSIF x = 8233 THEN
            sigmoid_f := 2011;
        ELSIF x = 8234 THEN
            sigmoid_f := 2011;
        ELSIF x = 8235 THEN
            sigmoid_f := 2011;
        ELSIF x = 8236 THEN
            sigmoid_f := 2011;
        ELSIF x = 8237 THEN
            sigmoid_f := 2011;
        ELSIF x = 8238 THEN
            sigmoid_f := 2011;
        ELSIF x = 8239 THEN
            sigmoid_f := 2011;
        ELSIF x = 8240 THEN
            sigmoid_f := 2011;
        ELSIF x = 8241 THEN
            sigmoid_f := 2011;
        ELSIF x = 8242 THEN
            sigmoid_f := 2011;
        ELSIF x = 8243 THEN
            sigmoid_f := 2011;
        ELSIF x = 8244 THEN
            sigmoid_f := 2011;
        ELSIF x = 8245 THEN
            sigmoid_f := 2011;
        ELSIF x = 8246 THEN
            sigmoid_f := 2011;
        ELSIF x = 8247 THEN
            sigmoid_f := 2011;
        ELSIF x = 8248 THEN
            sigmoid_f := 2011;
        ELSIF x = 8249 THEN
            sigmoid_f := 2011;
        ELSIF x = 8250 THEN
            sigmoid_f := 2011;
        ELSIF x = 8251 THEN
            sigmoid_f := 2011;
        ELSIF x = 8252 THEN
            sigmoid_f := 2011;
        ELSIF x = 8253 THEN
            sigmoid_f := 2012;
        ELSIF x = 8254 THEN
            sigmoid_f := 2012;
        ELSIF x = 8255 THEN
            sigmoid_f := 2012;
        ELSIF x = 8256 THEN
            sigmoid_f := 2012;
        ELSIF x = 8257 THEN
            sigmoid_f := 2012;
        ELSIF x = 8258 THEN
            sigmoid_f := 2012;
        ELSIF x = 8259 THEN
            sigmoid_f := 2012;
        ELSIF x = 8260 THEN
            sigmoid_f := 2012;
        ELSIF x = 8261 THEN
            sigmoid_f := 2012;
        ELSIF x = 8262 THEN
            sigmoid_f := 2012;
        ELSIF x = 8263 THEN
            sigmoid_f := 2012;
        ELSIF x = 8264 THEN
            sigmoid_f := 2012;
        ELSIF x = 8265 THEN
            sigmoid_f := 2012;
        ELSIF x = 8266 THEN
            sigmoid_f := 2012;
        ELSIF x = 8267 THEN
            sigmoid_f := 2012;
        ELSIF x = 8268 THEN
            sigmoid_f := 2012;
        ELSIF x = 8269 THEN
            sigmoid_f := 2012;
        ELSIF x = 8270 THEN
            sigmoid_f := 2012;
        ELSIF x = 8271 THEN
            sigmoid_f := 2012;
        ELSIF x = 8272 THEN
            sigmoid_f := 2012;
        ELSIF x = 8273 THEN
            sigmoid_f := 2012;
        ELSIF x = 8274 THEN
            sigmoid_f := 2012;
        ELSIF x = 8275 THEN
            sigmoid_f := 2012;
        ELSIF x = 8276 THEN
            sigmoid_f := 2012;
        ELSIF x = 8277 THEN
            sigmoid_f := 2012;
        ELSIF x = 8278 THEN
            sigmoid_f := 2012;
        ELSIF x = 8279 THEN
            sigmoid_f := 2012;
        ELSIF x = 8280 THEN
            sigmoid_f := 2012;
        ELSIF x = 8281 THEN
            sigmoid_f := 2012;
        ELSIF x = 8282 THEN
            sigmoid_f := 2012;
        ELSIF x = 8283 THEN
            sigmoid_f := 2012;
        ELSIF x = 8284 THEN
            sigmoid_f := 2012;
        ELSIF x = 8285 THEN
            sigmoid_f := 2012;
        ELSIF x = 8286 THEN
            sigmoid_f := 2012;
        ELSIF x = 8287 THEN
            sigmoid_f := 2012;
        ELSIF x = 8288 THEN
            sigmoid_f := 2012;
        ELSIF x = 8289 THEN
            sigmoid_f := 2012;
        ELSIF x = 8290 THEN
            sigmoid_f := 2012;
        ELSIF x = 8291 THEN
            sigmoid_f := 2012;
        ELSIF x = 8292 THEN
            sigmoid_f := 2012;
        ELSIF x = 8293 THEN
            sigmoid_f := 2012;
        ELSIF x = 8294 THEN
            sigmoid_f := 2012;
        ELSIF x = 8295 THEN
            sigmoid_f := 2012;
        ELSIF x = 8296 THEN
            sigmoid_f := 2012;
        ELSIF x = 8297 THEN
            sigmoid_f := 2012;
        ELSIF x = 8298 THEN
            sigmoid_f := 2012;
        ELSIF x = 8299 THEN
            sigmoid_f := 2012;
        ELSIF x = 8300 THEN
            sigmoid_f := 2012;
        ELSIF x = 8301 THEN
            sigmoid_f := 2012;
        ELSIF x = 8302 THEN
            sigmoid_f := 2012;
        ELSIF x = 8303 THEN
            sigmoid_f := 2012;
        ELSIF x = 8304 THEN
            sigmoid_f := 2012;
        ELSIF x = 8305 THEN
            sigmoid_f := 2012;
        ELSIF x = 8306 THEN
            sigmoid_f := 2012;
        ELSIF x = 8307 THEN
            sigmoid_f := 2012;
        ELSIF x = 8308 THEN
            sigmoid_f := 2012;
        ELSIF x = 8309 THEN
            sigmoid_f := 2012;
        ELSIF x = 8310 THEN
            sigmoid_f := 2012;
        ELSIF x = 8311 THEN
            sigmoid_f := 2012;
        ELSIF x = 8312 THEN
            sigmoid_f := 2012;
        ELSIF x = 8313 THEN
            sigmoid_f := 2013;
        ELSIF x = 8314 THEN
            sigmoid_f := 2013;
        ELSIF x = 8315 THEN
            sigmoid_f := 2013;
        ELSIF x = 8316 THEN
            sigmoid_f := 2013;
        ELSIF x = 8317 THEN
            sigmoid_f := 2013;
        ELSIF x = 8318 THEN
            sigmoid_f := 2013;
        ELSIF x = 8319 THEN
            sigmoid_f := 2013;
        ELSIF x = 8320 THEN
            sigmoid_f := 2013;
        ELSIF x = 8321 THEN
            sigmoid_f := 2013;
        ELSIF x = 8322 THEN
            sigmoid_f := 2013;
        ELSIF x = 8323 THEN
            sigmoid_f := 2013;
        ELSIF x = 8324 THEN
            sigmoid_f := 2013;
        ELSIF x = 8325 THEN
            sigmoid_f := 2013;
        ELSIF x = 8326 THEN
            sigmoid_f := 2013;
        ELSIF x = 8327 THEN
            sigmoid_f := 2013;
        ELSIF x = 8328 THEN
            sigmoid_f := 2013;
        ELSIF x = 8329 THEN
            sigmoid_f := 2013;
        ELSIF x = 8330 THEN
            sigmoid_f := 2013;
        ELSIF x = 8331 THEN
            sigmoid_f := 2013;
        ELSIF x = 8332 THEN
            sigmoid_f := 2013;
        ELSIF x = 8333 THEN
            sigmoid_f := 2013;
        ELSIF x = 8334 THEN
            sigmoid_f := 2013;
        ELSIF x = 8335 THEN
            sigmoid_f := 2013;
        ELSIF x = 8336 THEN
            sigmoid_f := 2013;
        ELSIF x = 8337 THEN
            sigmoid_f := 2013;
        ELSIF x = 8338 THEN
            sigmoid_f := 2013;
        ELSIF x = 8339 THEN
            sigmoid_f := 2013;
        ELSIF x = 8340 THEN
            sigmoid_f := 2013;
        ELSIF x = 8341 THEN
            sigmoid_f := 2013;
        ELSIF x = 8342 THEN
            sigmoid_f := 2013;
        ELSIF x = 8343 THEN
            sigmoid_f := 2013;
        ELSIF x = 8344 THEN
            sigmoid_f := 2013;
        ELSIF x = 8345 THEN
            sigmoid_f := 2013;
        ELSIF x = 8346 THEN
            sigmoid_f := 2013;
        ELSIF x = 8347 THEN
            sigmoid_f := 2013;
        ELSIF x = 8348 THEN
            sigmoid_f := 2013;
        ELSIF x = 8349 THEN
            sigmoid_f := 2013;
        ELSIF x = 8350 THEN
            sigmoid_f := 2013;
        ELSIF x = 8351 THEN
            sigmoid_f := 2013;
        ELSIF x = 8352 THEN
            sigmoid_f := 2013;
        ELSIF x = 8353 THEN
            sigmoid_f := 2013;
        ELSIF x = 8354 THEN
            sigmoid_f := 2013;
        ELSIF x = 8355 THEN
            sigmoid_f := 2013;
        ELSIF x = 8356 THEN
            sigmoid_f := 2013;
        ELSIF x = 8357 THEN
            sigmoid_f := 2013;
        ELSIF x = 8358 THEN
            sigmoid_f := 2013;
        ELSIF x = 8359 THEN
            sigmoid_f := 2013;
        ELSIF x = 8360 THEN
            sigmoid_f := 2013;
        ELSIF x = 8361 THEN
            sigmoid_f := 2013;
        ELSIF x = 8362 THEN
            sigmoid_f := 2013;
        ELSIF x = 8363 THEN
            sigmoid_f := 2013;
        ELSIF x = 8364 THEN
            sigmoid_f := 2013;
        ELSIF x = 8365 THEN
            sigmoid_f := 2013;
        ELSIF x = 8366 THEN
            sigmoid_f := 2013;
        ELSIF x = 8367 THEN
            sigmoid_f := 2013;
        ELSIF x = 8368 THEN
            sigmoid_f := 2013;
        ELSIF x = 8369 THEN
            sigmoid_f := 2013;
        ELSIF x = 8370 THEN
            sigmoid_f := 2013;
        ELSIF x = 8371 THEN
            sigmoid_f := 2013;
        ELSIF x = 8372 THEN
            sigmoid_f := 2013;
        ELSIF x = 8373 THEN
            sigmoid_f := 2014;
        ELSIF x = 8374 THEN
            sigmoid_f := 2014;
        ELSIF x = 8375 THEN
            sigmoid_f := 2014;
        ELSIF x = 8376 THEN
            sigmoid_f := 2014;
        ELSIF x = 8377 THEN
            sigmoid_f := 2014;
        ELSIF x = 8378 THEN
            sigmoid_f := 2014;
        ELSIF x = 8379 THEN
            sigmoid_f := 2014;
        ELSIF x = 8380 THEN
            sigmoid_f := 2014;
        ELSIF x = 8381 THEN
            sigmoid_f := 2014;
        ELSIF x = 8382 THEN
            sigmoid_f := 2014;
        ELSIF x = 8383 THEN
            sigmoid_f := 2014;
        ELSIF x = 8384 THEN
            sigmoid_f := 2014;
        ELSIF x = 8385 THEN
            sigmoid_f := 2014;
        ELSIF x = 8386 THEN
            sigmoid_f := 2014;
        ELSIF x = 8387 THEN
            sigmoid_f := 2014;
        ELSIF x = 8388 THEN
            sigmoid_f := 2014;
        ELSIF x = 8389 THEN
            sigmoid_f := 2014;
        ELSIF x = 8390 THEN
            sigmoid_f := 2014;
        ELSIF x = 8391 THEN
            sigmoid_f := 2014;
        ELSIF x = 8392 THEN
            sigmoid_f := 2014;
        ELSIF x = 8393 THEN
            sigmoid_f := 2014;
        ELSIF x = 8394 THEN
            sigmoid_f := 2014;
        ELSIF x = 8395 THEN
            sigmoid_f := 2014;
        ELSIF x = 8396 THEN
            sigmoid_f := 2014;
        ELSIF x = 8397 THEN
            sigmoid_f := 2014;
        ELSIF x = 8398 THEN
            sigmoid_f := 2014;
        ELSIF x = 8399 THEN
            sigmoid_f := 2014;
        ELSIF x = 8400 THEN
            sigmoid_f := 2014;
        ELSIF x = 8401 THEN
            sigmoid_f := 2014;
        ELSIF x = 8402 THEN
            sigmoid_f := 2014;
        ELSIF x = 8403 THEN
            sigmoid_f := 2014;
        ELSIF x = 8404 THEN
            sigmoid_f := 2014;
        ELSIF x = 8405 THEN
            sigmoid_f := 2014;
        ELSIF x = 8406 THEN
            sigmoid_f := 2014;
        ELSIF x = 8407 THEN
            sigmoid_f := 2014;
        ELSIF x = 8408 THEN
            sigmoid_f := 2014;
        ELSIF x = 8409 THEN
            sigmoid_f := 2014;
        ELSIF x = 8410 THEN
            sigmoid_f := 2014;
        ELSIF x = 8411 THEN
            sigmoid_f := 2014;
        ELSIF x = 8412 THEN
            sigmoid_f := 2014;
        ELSIF x = 8413 THEN
            sigmoid_f := 2014;
        ELSIF x = 8414 THEN
            sigmoid_f := 2014;
        ELSIF x = 8415 THEN
            sigmoid_f := 2014;
        ELSIF x = 8416 THEN
            sigmoid_f := 2014;
        ELSIF x = 8417 THEN
            sigmoid_f := 2014;
        ELSIF x = 8418 THEN
            sigmoid_f := 2014;
        ELSIF x = 8419 THEN
            sigmoid_f := 2014;
        ELSIF x = 8420 THEN
            sigmoid_f := 2014;
        ELSIF x = 8421 THEN
            sigmoid_f := 2014;
        ELSIF x = 8422 THEN
            sigmoid_f := 2014;
        ELSIF x = 8423 THEN
            sigmoid_f := 2014;
        ELSIF x = 8424 THEN
            sigmoid_f := 2014;
        ELSIF x = 8425 THEN
            sigmoid_f := 2014;
        ELSIF x = 8426 THEN
            sigmoid_f := 2014;
        ELSIF x = 8427 THEN
            sigmoid_f := 2014;
        ELSIF x = 8428 THEN
            sigmoid_f := 2014;
        ELSIF x = 8429 THEN
            sigmoid_f := 2014;
        ELSIF x = 8430 THEN
            sigmoid_f := 2014;
        ELSIF x = 8431 THEN
            sigmoid_f := 2014;
        ELSIF x = 8432 THEN
            sigmoid_f := 2014;
        ELSIF x = 8433 THEN
            sigmoid_f := 2015;
        ELSIF x = 8434 THEN
            sigmoid_f := 2015;
        ELSIF x = 8435 THEN
            sigmoid_f := 2015;
        ELSIF x = 8436 THEN
            sigmoid_f := 2015;
        ELSIF x = 8437 THEN
            sigmoid_f := 2015;
        ELSIF x = 8438 THEN
            sigmoid_f := 2015;
        ELSIF x = 8439 THEN
            sigmoid_f := 2015;
        ELSIF x = 8440 THEN
            sigmoid_f := 2015;
        ELSIF x = 8441 THEN
            sigmoid_f := 2015;
        ELSIF x = 8442 THEN
            sigmoid_f := 2015;
        ELSIF x = 8443 THEN
            sigmoid_f := 2015;
        ELSIF x = 8444 THEN
            sigmoid_f := 2015;
        ELSIF x = 8445 THEN
            sigmoid_f := 2015;
        ELSIF x = 8446 THEN
            sigmoid_f := 2015;
        ELSIF x = 8447 THEN
            sigmoid_f := 2015;
        ELSIF x = 8448 THEN
            sigmoid_f := 2015;
        ELSIF x = 8449 THEN
            sigmoid_f := 2015;
        ELSIF x = 8450 THEN
            sigmoid_f := 2015;
        ELSIF x = 8451 THEN
            sigmoid_f := 2015;
        ELSIF x = 8452 THEN
            sigmoid_f := 2015;
        ELSIF x = 8453 THEN
            sigmoid_f := 2015;
        ELSIF x = 8454 THEN
            sigmoid_f := 2015;
        ELSIF x = 8455 THEN
            sigmoid_f := 2015;
        ELSIF x = 8456 THEN
            sigmoid_f := 2015;
        ELSIF x = 8457 THEN
            sigmoid_f := 2015;
        ELSIF x = 8458 THEN
            sigmoid_f := 2015;
        ELSIF x = 8459 THEN
            sigmoid_f := 2015;
        ELSIF x = 8460 THEN
            sigmoid_f := 2015;
        ELSIF x = 8461 THEN
            sigmoid_f := 2015;
        ELSIF x = 8462 THEN
            sigmoid_f := 2015;
        ELSIF x = 8463 THEN
            sigmoid_f := 2015;
        ELSIF x = 8464 THEN
            sigmoid_f := 2015;
        ELSIF x = 8465 THEN
            sigmoid_f := 2015;
        ELSIF x = 8466 THEN
            sigmoid_f := 2015;
        ELSIF x = 8467 THEN
            sigmoid_f := 2015;
        ELSIF x = 8468 THEN
            sigmoid_f := 2015;
        ELSIF x = 8469 THEN
            sigmoid_f := 2015;
        ELSIF x = 8470 THEN
            sigmoid_f := 2015;
        ELSIF x = 8471 THEN
            sigmoid_f := 2015;
        ELSIF x = 8472 THEN
            sigmoid_f := 2015;
        ELSIF x = 8473 THEN
            sigmoid_f := 2015;
        ELSIF x = 8474 THEN
            sigmoid_f := 2015;
        ELSIF x = 8475 THEN
            sigmoid_f := 2015;
        ELSIF x = 8476 THEN
            sigmoid_f := 2015;
        ELSIF x = 8477 THEN
            sigmoid_f := 2015;
        ELSIF x = 8478 THEN
            sigmoid_f := 2015;
        ELSIF x = 8479 THEN
            sigmoid_f := 2015;
        ELSIF x = 8480 THEN
            sigmoid_f := 2015;
        ELSIF x = 8481 THEN
            sigmoid_f := 2015;
        ELSIF x = 8482 THEN
            sigmoid_f := 2015;
        ELSIF x = 8483 THEN
            sigmoid_f := 2015;
        ELSIF x = 8484 THEN
            sigmoid_f := 2015;
        ELSIF x = 8485 THEN
            sigmoid_f := 2015;
        ELSIF x = 8486 THEN
            sigmoid_f := 2015;
        ELSIF x = 8487 THEN
            sigmoid_f := 2015;
        ELSIF x = 8488 THEN
            sigmoid_f := 2015;
        ELSIF x = 8489 THEN
            sigmoid_f := 2015;
        ELSIF x = 8490 THEN
            sigmoid_f := 2015;
        ELSIF x = 8491 THEN
            sigmoid_f := 2015;
        ELSIF x = 8492 THEN
            sigmoid_f := 2015;
        ELSIF x = 8493 THEN
            sigmoid_f := 2015;
        ELSIF x = 8494 THEN
            sigmoid_f := 2016;
        ELSIF x = 8495 THEN
            sigmoid_f := 2016;
        ELSIF x = 8496 THEN
            sigmoid_f := 2016;
        ELSIF x = 8497 THEN
            sigmoid_f := 2016;
        ELSIF x = 8498 THEN
            sigmoid_f := 2016;
        ELSIF x = 8499 THEN
            sigmoid_f := 2016;
        ELSIF x = 8500 THEN
            sigmoid_f := 2016;
        ELSIF x = 8501 THEN
            sigmoid_f := 2016;
        ELSIF x = 8502 THEN
            sigmoid_f := 2016;
        ELSIF x = 8503 THEN
            sigmoid_f := 2016;
        ELSIF x = 8504 THEN
            sigmoid_f := 2016;
        ELSIF x = 8505 THEN
            sigmoid_f := 2016;
        ELSIF x = 8506 THEN
            sigmoid_f := 2016;
        ELSIF x = 8507 THEN
            sigmoid_f := 2016;
        ELSIF x = 8508 THEN
            sigmoid_f := 2016;
        ELSIF x = 8509 THEN
            sigmoid_f := 2016;
        ELSIF x = 8510 THEN
            sigmoid_f := 2016;
        ELSIF x = 8511 THEN
            sigmoid_f := 2016;
        ELSIF x = 8512 THEN
            sigmoid_f := 2016;
        ELSIF x = 8513 THEN
            sigmoid_f := 2016;
        ELSIF x = 8514 THEN
            sigmoid_f := 2016;
        ELSIF x = 8515 THEN
            sigmoid_f := 2016;
        ELSIF x = 8516 THEN
            sigmoid_f := 2016;
        ELSIF x = 8517 THEN
            sigmoid_f := 2016;
        ELSIF x = 8518 THEN
            sigmoid_f := 2016;
        ELSIF x = 8519 THEN
            sigmoid_f := 2016;
        ELSIF x = 8520 THEN
            sigmoid_f := 2016;
        ELSIF x = 8521 THEN
            sigmoid_f := 2016;
        ELSIF x = 8522 THEN
            sigmoid_f := 2016;
        ELSIF x = 8523 THEN
            sigmoid_f := 2016;
        ELSIF x = 8524 THEN
            sigmoid_f := 2016;
        ELSIF x = 8525 THEN
            sigmoid_f := 2016;
        ELSIF x = 8526 THEN
            sigmoid_f := 2016;
        ELSIF x = 8527 THEN
            sigmoid_f := 2016;
        ELSIF x = 8528 THEN
            sigmoid_f := 2016;
        ELSIF x = 8529 THEN
            sigmoid_f := 2016;
        ELSIF x = 8530 THEN
            sigmoid_f := 2016;
        ELSIF x = 8531 THEN
            sigmoid_f := 2016;
        ELSIF x = 8532 THEN
            sigmoid_f := 2016;
        ELSIF x = 8533 THEN
            sigmoid_f := 2016;
        ELSIF x = 8534 THEN
            sigmoid_f := 2016;
        ELSIF x = 8535 THEN
            sigmoid_f := 2016;
        ELSIF x = 8536 THEN
            sigmoid_f := 2016;
        ELSIF x = 8537 THEN
            sigmoid_f := 2016;
        ELSIF x = 8538 THEN
            sigmoid_f := 2016;
        ELSIF x = 8539 THEN
            sigmoid_f := 2016;
        ELSIF x = 8540 THEN
            sigmoid_f := 2016;
        ELSIF x = 8541 THEN
            sigmoid_f := 2016;
        ELSIF x = 8542 THEN
            sigmoid_f := 2016;
        ELSIF x = 8543 THEN
            sigmoid_f := 2016;
        ELSIF x = 8544 THEN
            sigmoid_f := 2016;
        ELSIF x = 8545 THEN
            sigmoid_f := 2016;
        ELSIF x = 8546 THEN
            sigmoid_f := 2016;
        ELSIF x = 8547 THEN
            sigmoid_f := 2016;
        ELSIF x = 8548 THEN
            sigmoid_f := 2016;
        ELSIF x = 8549 THEN
            sigmoid_f := 2016;
        ELSIF x = 8550 THEN
            sigmoid_f := 2016;
        ELSIF x = 8551 THEN
            sigmoid_f := 2016;
        ELSIF x = 8552 THEN
            sigmoid_f := 2016;
        ELSIF x = 8553 THEN
            sigmoid_f := 2016;
        ELSIF x = 8554 THEN
            sigmoid_f := 2017;
        ELSIF x = 8555 THEN
            sigmoid_f := 2017;
        ELSIF x = 8556 THEN
            sigmoid_f := 2017;
        ELSIF x = 8557 THEN
            sigmoid_f := 2017;
        ELSIF x = 8558 THEN
            sigmoid_f := 2017;
        ELSIF x = 8559 THEN
            sigmoid_f := 2017;
        ELSIF x = 8560 THEN
            sigmoid_f := 2017;
        ELSIF x = 8561 THEN
            sigmoid_f := 2017;
        ELSIF x = 8562 THEN
            sigmoid_f := 2017;
        ELSIF x = 8563 THEN
            sigmoid_f := 2017;
        ELSIF x = 8564 THEN
            sigmoid_f := 2017;
        ELSIF x = 8565 THEN
            sigmoid_f := 2017;
        ELSIF x = 8566 THEN
            sigmoid_f := 2017;
        ELSIF x = 8567 THEN
            sigmoid_f := 2017;
        ELSIF x = 8568 THEN
            sigmoid_f := 2017;
        ELSIF x = 8569 THEN
            sigmoid_f := 2017;
        ELSIF x = 8570 THEN
            sigmoid_f := 2017;
        ELSIF x = 8571 THEN
            sigmoid_f := 2017;
        ELSIF x = 8572 THEN
            sigmoid_f := 2017;
        ELSIF x = 8573 THEN
            sigmoid_f := 2017;
        ELSIF x = 8574 THEN
            sigmoid_f := 2017;
        ELSIF x = 8575 THEN
            sigmoid_f := 2017;
        ELSIF x = 8576 THEN
            sigmoid_f := 2017;
        ELSIF x = 8577 THEN
            sigmoid_f := 2017;
        ELSIF x = 8578 THEN
            sigmoid_f := 2017;
        ELSIF x = 8579 THEN
            sigmoid_f := 2017;
        ELSIF x = 8580 THEN
            sigmoid_f := 2017;
        ELSIF x = 8581 THEN
            sigmoid_f := 2017;
        ELSIF x = 8582 THEN
            sigmoid_f := 2017;
        ELSIF x = 8583 THEN
            sigmoid_f := 2017;
        ELSIF x = 8584 THEN
            sigmoid_f := 2017;
        ELSIF x = 8585 THEN
            sigmoid_f := 2017;
        ELSIF x = 8586 THEN
            sigmoid_f := 2017;
        ELSIF x = 8587 THEN
            sigmoid_f := 2017;
        ELSIF x = 8588 THEN
            sigmoid_f := 2017;
        ELSIF x = 8589 THEN
            sigmoid_f := 2017;
        ELSIF x = 8590 THEN
            sigmoid_f := 2017;
        ELSIF x = 8591 THEN
            sigmoid_f := 2017;
        ELSIF x = 8592 THEN
            sigmoid_f := 2017;
        ELSIF x = 8593 THEN
            sigmoid_f := 2017;
        ELSIF x = 8594 THEN
            sigmoid_f := 2017;
        ELSIF x = 8595 THEN
            sigmoid_f := 2017;
        ELSIF x = 8596 THEN
            sigmoid_f := 2017;
        ELSIF x = 8597 THEN
            sigmoid_f := 2017;
        ELSIF x = 8598 THEN
            sigmoid_f := 2017;
        ELSIF x = 8599 THEN
            sigmoid_f := 2017;
        ELSIF x = 8600 THEN
            sigmoid_f := 2017;
        ELSIF x = 8601 THEN
            sigmoid_f := 2017;
        ELSIF x = 8602 THEN
            sigmoid_f := 2017;
        ELSIF x = 8603 THEN
            sigmoid_f := 2017;
        ELSIF x = 8604 THEN
            sigmoid_f := 2017;
        ELSIF x = 8605 THEN
            sigmoid_f := 2017;
        ELSIF x = 8606 THEN
            sigmoid_f := 2017;
        ELSIF x = 8607 THEN
            sigmoid_f := 2017;
        ELSIF x = 8608 THEN
            sigmoid_f := 2017;
        ELSIF x = 8609 THEN
            sigmoid_f := 2017;
        ELSIF x = 8610 THEN
            sigmoid_f := 2017;
        ELSIF x = 8611 THEN
            sigmoid_f := 2017;
        ELSIF x = 8612 THEN
            sigmoid_f := 2017;
        ELSIF x = 8613 THEN
            sigmoid_f := 2017;
        ELSIF x = 8614 THEN
            sigmoid_f := 2018;
        ELSIF x = 8615 THEN
            sigmoid_f := 2018;
        ELSIF x = 8616 THEN
            sigmoid_f := 2018;
        ELSIF x = 8617 THEN
            sigmoid_f := 2018;
        ELSIF x = 8618 THEN
            sigmoid_f := 2018;
        ELSIF x = 8619 THEN
            sigmoid_f := 2018;
        ELSIF x = 8620 THEN
            sigmoid_f := 2018;
        ELSIF x = 8621 THEN
            sigmoid_f := 2018;
        ELSIF x = 8622 THEN
            sigmoid_f := 2018;
        ELSIF x = 8623 THEN
            sigmoid_f := 2018;
        ELSIF x = 8624 THEN
            sigmoid_f := 2018;
        ELSIF x = 8625 THEN
            sigmoid_f := 2018;
        ELSIF x = 8626 THEN
            sigmoid_f := 2018;
        ELSIF x = 8627 THEN
            sigmoid_f := 2018;
        ELSIF x = 8628 THEN
            sigmoid_f := 2018;
        ELSIF x = 8629 THEN
            sigmoid_f := 2018;
        ELSIF x = 8630 THEN
            sigmoid_f := 2018;
        ELSIF x = 8631 THEN
            sigmoid_f := 2018;
        ELSIF x = 8632 THEN
            sigmoid_f := 2018;
        ELSIF x = 8633 THEN
            sigmoid_f := 2018;
        ELSIF x = 8634 THEN
            sigmoid_f := 2018;
        ELSIF x = 8635 THEN
            sigmoid_f := 2018;
        ELSIF x = 8636 THEN
            sigmoid_f := 2018;
        ELSIF x = 8637 THEN
            sigmoid_f := 2018;
        ELSIF x = 8638 THEN
            sigmoid_f := 2018;
        ELSIF x = 8639 THEN
            sigmoid_f := 2018;
        ELSIF x = 8640 THEN
            sigmoid_f := 2018;
        ELSIF x = 8641 THEN
            sigmoid_f := 2018;
        ELSIF x = 8642 THEN
            sigmoid_f := 2018;
        ELSIF x = 8643 THEN
            sigmoid_f := 2018;
        ELSIF x = 8644 THEN
            sigmoid_f := 2018;
        ELSIF x = 8645 THEN
            sigmoid_f := 2018;
        ELSIF x = 8646 THEN
            sigmoid_f := 2018;
        ELSIF x = 8647 THEN
            sigmoid_f := 2018;
        ELSIF x = 8648 THEN
            sigmoid_f := 2018;
        ELSIF x = 8649 THEN
            sigmoid_f := 2018;
        ELSIF x = 8650 THEN
            sigmoid_f := 2018;
        ELSIF x = 8651 THEN
            sigmoid_f := 2018;
        ELSIF x = 8652 THEN
            sigmoid_f := 2018;
        ELSIF x = 8653 THEN
            sigmoid_f := 2018;
        ELSIF x = 8654 THEN
            sigmoid_f := 2018;
        ELSIF x = 8655 THEN
            sigmoid_f := 2018;
        ELSIF x = 8656 THEN
            sigmoid_f := 2018;
        ELSIF x = 8657 THEN
            sigmoid_f := 2018;
        ELSIF x = 8658 THEN
            sigmoid_f := 2018;
        ELSIF x = 8659 THEN
            sigmoid_f := 2018;
        ELSIF x = 8660 THEN
            sigmoid_f := 2018;
        ELSIF x = 8661 THEN
            sigmoid_f := 2018;
        ELSIF x = 8662 THEN
            sigmoid_f := 2018;
        ELSIF x = 8663 THEN
            sigmoid_f := 2018;
        ELSIF x = 8664 THEN
            sigmoid_f := 2018;
        ELSIF x = 8665 THEN
            sigmoid_f := 2018;
        ELSIF x = 8666 THEN
            sigmoid_f := 2018;
        ELSIF x = 8667 THEN
            sigmoid_f := 2018;
        ELSIF x = 8668 THEN
            sigmoid_f := 2018;
        ELSIF x = 8669 THEN
            sigmoid_f := 2018;
        ELSIF x = 8670 THEN
            sigmoid_f := 2018;
        ELSIF x = 8671 THEN
            sigmoid_f := 2018;
        ELSIF x = 8672 THEN
            sigmoid_f := 2018;
        ELSIF x = 8673 THEN
            sigmoid_f := 2018;
        ELSIF x = 8674 THEN
            sigmoid_f := 2019;
        ELSIF x = 8675 THEN
            sigmoid_f := 2019;
        ELSIF x = 8676 THEN
            sigmoid_f := 2019;
        ELSIF x = 8677 THEN
            sigmoid_f := 2019;
        ELSIF x = 8678 THEN
            sigmoid_f := 2019;
        ELSIF x = 8679 THEN
            sigmoid_f := 2019;
        ELSIF x = 8680 THEN
            sigmoid_f := 2019;
        ELSIF x = 8681 THEN
            sigmoid_f := 2019;
        ELSIF x = 8682 THEN
            sigmoid_f := 2019;
        ELSIF x = 8683 THEN
            sigmoid_f := 2019;
        ELSIF x = 8684 THEN
            sigmoid_f := 2019;
        ELSIF x = 8685 THEN
            sigmoid_f := 2019;
        ELSIF x = 8686 THEN
            sigmoid_f := 2019;
        ELSIF x = 8687 THEN
            sigmoid_f := 2019;
        ELSIF x = 8688 THEN
            sigmoid_f := 2019;
        ELSIF x = 8689 THEN
            sigmoid_f := 2019;
        ELSIF x = 8690 THEN
            sigmoid_f := 2019;
        ELSIF x = 8691 THEN
            sigmoid_f := 2019;
        ELSIF x = 8692 THEN
            sigmoid_f := 2019;
        ELSIF x = 8693 THEN
            sigmoid_f := 2019;
        ELSIF x = 8694 THEN
            sigmoid_f := 2019;
        ELSIF x = 8695 THEN
            sigmoid_f := 2019;
        ELSIF x = 8696 THEN
            sigmoid_f := 2019;
        ELSIF x = 8697 THEN
            sigmoid_f := 2019;
        ELSIF x = 8698 THEN
            sigmoid_f := 2019;
        ELSIF x = 8699 THEN
            sigmoid_f := 2019;
        ELSIF x = 8700 THEN
            sigmoid_f := 2019;
        ELSIF x = 8701 THEN
            sigmoid_f := 2019;
        ELSIF x = 8702 THEN
            sigmoid_f := 2019;
        ELSIF x = 8703 THEN
            sigmoid_f := 2019;
        ELSIF x = 8704 THEN
            sigmoid_f := 2019;
        ELSIF x = 8705 THEN
            sigmoid_f := 2019;
        ELSIF x = 8706 THEN
            sigmoid_f := 2019;
        ELSIF x = 8707 THEN
            sigmoid_f := 2019;
        ELSIF x = 8708 THEN
            sigmoid_f := 2019;
        ELSIF x = 8709 THEN
            sigmoid_f := 2019;
        ELSIF x = 8710 THEN
            sigmoid_f := 2019;
        ELSIF x = 8711 THEN
            sigmoid_f := 2019;
        ELSIF x = 8712 THEN
            sigmoid_f := 2019;
        ELSIF x = 8713 THEN
            sigmoid_f := 2019;
        ELSIF x = 8714 THEN
            sigmoid_f := 2019;
        ELSIF x = 8715 THEN
            sigmoid_f := 2019;
        ELSIF x = 8716 THEN
            sigmoid_f := 2019;
        ELSIF x = 8717 THEN
            sigmoid_f := 2019;
        ELSIF x = 8718 THEN
            sigmoid_f := 2019;
        ELSIF x = 8719 THEN
            sigmoid_f := 2019;
        ELSIF x = 8720 THEN
            sigmoid_f := 2019;
        ELSIF x = 8721 THEN
            sigmoid_f := 2019;
        ELSIF x = 8722 THEN
            sigmoid_f := 2019;
        ELSIF x = 8723 THEN
            sigmoid_f := 2019;
        ELSIF x = 8724 THEN
            sigmoid_f := 2019;
        ELSIF x = 8725 THEN
            sigmoid_f := 2019;
        ELSIF x = 8726 THEN
            sigmoid_f := 2019;
        ELSIF x = 8727 THEN
            sigmoid_f := 2019;
        ELSIF x = 8728 THEN
            sigmoid_f := 2019;
        ELSIF x = 8729 THEN
            sigmoid_f := 2019;
        ELSIF x = 8730 THEN
            sigmoid_f := 2019;
        ELSIF x = 8731 THEN
            sigmoid_f := 2019;
        ELSIF x = 8732 THEN
            sigmoid_f := 2019;
        ELSIF x = 8733 THEN
            sigmoid_f := 2019;
        ELSIF x = 8734 THEN
            sigmoid_f := 2019;
        ELSIF x = 8735 THEN
            sigmoid_f := 2019;
        ELSIF x = 8736 THEN
            sigmoid_f := 2019;
        ELSIF x = 8737 THEN
            sigmoid_f := 2019;
        ELSIF x = 8738 THEN
            sigmoid_f := 2019;
        ELSIF x = 8739 THEN
            sigmoid_f := 2019;
        ELSIF x = 8740 THEN
            sigmoid_f := 2019;
        ELSIF x = 8741 THEN
            sigmoid_f := 2019;
        ELSIF x = 8742 THEN
            sigmoid_f := 2019;
        ELSIF x = 8743 THEN
            sigmoid_f := 2019;
        ELSIF x = 8744 THEN
            sigmoid_f := 2019;
        ELSIF x = 8745 THEN
            sigmoid_f := 2019;
        ELSIF x = 8746 THEN
            sigmoid_f := 2019;
        ELSIF x = 8747 THEN
            sigmoid_f := 2019;
        ELSIF x = 8748 THEN
            sigmoid_f := 2019;
        ELSIF x = 8749 THEN
            sigmoid_f := 2019;
        ELSIF x = 8750 THEN
            sigmoid_f := 2019;
        ELSIF x = 8751 THEN
            sigmoid_f := 2019;
        ELSIF x = 8752 THEN
            sigmoid_f := 2019;
        ELSIF x = 8753 THEN
            sigmoid_f := 2019;
        ELSIF x = 8754 THEN
            sigmoid_f := 2019;
        ELSIF x = 8755 THEN
            sigmoid_f := 2019;
        ELSIF x = 8756 THEN
            sigmoid_f := 2019;
        ELSIF x = 8757 THEN
            sigmoid_f := 2019;
        ELSIF x = 8758 THEN
            sigmoid_f := 2019;
        ELSIF x = 8759 THEN
            sigmoid_f := 2019;
        ELSIF x = 8760 THEN
            sigmoid_f := 2019;
        ELSIF x = 8761 THEN
            sigmoid_f := 2019;
        ELSIF x = 8762 THEN
            sigmoid_f := 2019;
        ELSIF x = 8763 THEN
            sigmoid_f := 2019;
        ELSIF x = 8764 THEN
            sigmoid_f := 2019;
        ELSIF x = 8765 THEN
            sigmoid_f := 2019;
        ELSIF x = 8766 THEN
            sigmoid_f := 2020;
        ELSIF x = 8767 THEN
            sigmoid_f := 2020;
        ELSIF x = 8768 THEN
            sigmoid_f := 2020;
        ELSIF x = 8769 THEN
            sigmoid_f := 2020;
        ELSIF x = 8770 THEN
            sigmoid_f := 2020;
        ELSIF x = 8771 THEN
            sigmoid_f := 2020;
        ELSIF x = 8772 THEN
            sigmoid_f := 2020;
        ELSIF x = 8773 THEN
            sigmoid_f := 2020;
        ELSIF x = 8774 THEN
            sigmoid_f := 2020;
        ELSIF x = 8775 THEN
            sigmoid_f := 2020;
        ELSIF x = 8776 THEN
            sigmoid_f := 2020;
        ELSIF x = 8777 THEN
            sigmoid_f := 2020;
        ELSIF x = 8778 THEN
            sigmoid_f := 2020;
        ELSIF x = 8779 THEN
            sigmoid_f := 2020;
        ELSIF x = 8780 THEN
            sigmoid_f := 2020;
        ELSIF x = 8781 THEN
            sigmoid_f := 2020;
        ELSIF x = 8782 THEN
            sigmoid_f := 2020;
        ELSIF x = 8783 THEN
            sigmoid_f := 2020;
        ELSIF x = 8784 THEN
            sigmoid_f := 2020;
        ELSIF x = 8785 THEN
            sigmoid_f := 2020;
        ELSIF x = 8786 THEN
            sigmoid_f := 2020;
        ELSIF x = 8787 THEN
            sigmoid_f := 2020;
        ELSIF x = 8788 THEN
            sigmoid_f := 2020;
        ELSIF x = 8789 THEN
            sigmoid_f := 2020;
        ELSIF x = 8790 THEN
            sigmoid_f := 2020;
        ELSIF x = 8791 THEN
            sigmoid_f := 2020;
        ELSIF x = 8792 THEN
            sigmoid_f := 2020;
        ELSIF x = 8793 THEN
            sigmoid_f := 2020;
        ELSIF x = 8794 THEN
            sigmoid_f := 2020;
        ELSIF x = 8795 THEN
            sigmoid_f := 2020;
        ELSIF x = 8796 THEN
            sigmoid_f := 2020;
        ELSIF x = 8797 THEN
            sigmoid_f := 2020;
        ELSIF x = 8798 THEN
            sigmoid_f := 2020;
        ELSIF x = 8799 THEN
            sigmoid_f := 2020;
        ELSIF x = 8800 THEN
            sigmoid_f := 2020;
        ELSIF x = 8801 THEN
            sigmoid_f := 2020;
        ELSIF x = 8802 THEN
            sigmoid_f := 2020;
        ELSIF x = 8803 THEN
            sigmoid_f := 2020;
        ELSIF x = 8804 THEN
            sigmoid_f := 2020;
        ELSIF x = 8805 THEN
            sigmoid_f := 2020;
        ELSIF x = 8806 THEN
            sigmoid_f := 2020;
        ELSIF x = 8807 THEN
            sigmoid_f := 2020;
        ELSIF x = 8808 THEN
            sigmoid_f := 2020;
        ELSIF x = 8809 THEN
            sigmoid_f := 2020;
        ELSIF x = 8810 THEN
            sigmoid_f := 2020;
        ELSIF x = 8811 THEN
            sigmoid_f := 2020;
        ELSIF x = 8812 THEN
            sigmoid_f := 2020;
        ELSIF x = 8813 THEN
            sigmoid_f := 2020;
        ELSIF x = 8814 THEN
            sigmoid_f := 2020;
        ELSIF x = 8815 THEN
            sigmoid_f := 2020;
        ELSIF x = 8816 THEN
            sigmoid_f := 2020;
        ELSIF x = 8817 THEN
            sigmoid_f := 2020;
        ELSIF x = 8818 THEN
            sigmoid_f := 2020;
        ELSIF x = 8819 THEN
            sigmoid_f := 2020;
        ELSIF x = 8820 THEN
            sigmoid_f := 2020;
        ELSIF x = 8821 THEN
            sigmoid_f := 2020;
        ELSIF x = 8822 THEN
            sigmoid_f := 2020;
        ELSIF x = 8823 THEN
            sigmoid_f := 2020;
        ELSIF x = 8824 THEN
            sigmoid_f := 2020;
        ELSIF x = 8825 THEN
            sigmoid_f := 2020;
        ELSIF x = 8826 THEN
            sigmoid_f := 2020;
        ELSIF x = 8827 THEN
            sigmoid_f := 2020;
        ELSIF x = 8828 THEN
            sigmoid_f := 2020;
        ELSIF x = 8829 THEN
            sigmoid_f := 2020;
        ELSIF x = 8830 THEN
            sigmoid_f := 2020;
        ELSIF x = 8831 THEN
            sigmoid_f := 2020;
        ELSIF x = 8832 THEN
            sigmoid_f := 2020;
        ELSIF x = 8833 THEN
            sigmoid_f := 2020;
        ELSIF x = 8834 THEN
            sigmoid_f := 2020;
        ELSIF x = 8835 THEN
            sigmoid_f := 2020;
        ELSIF x = 8836 THEN
            sigmoid_f := 2020;
        ELSIF x = 8837 THEN
            sigmoid_f := 2020;
        ELSIF x = 8838 THEN
            sigmoid_f := 2020;
        ELSIF x = 8839 THEN
            sigmoid_f := 2020;
        ELSIF x = 8840 THEN
            sigmoid_f := 2020;
        ELSIF x = 8841 THEN
            sigmoid_f := 2020;
        ELSIF x = 8842 THEN
            sigmoid_f := 2020;
        ELSIF x = 8843 THEN
            sigmoid_f := 2020;
        ELSIF x = 8844 THEN
            sigmoid_f := 2020;
        ELSIF x = 8845 THEN
            sigmoid_f := 2020;
        ELSIF x = 8846 THEN
            sigmoid_f := 2020;
        ELSIF x = 8847 THEN
            sigmoid_f := 2020;
        ELSIF x = 8848 THEN
            sigmoid_f := 2021;
        ELSIF x = 8849 THEN
            sigmoid_f := 2021;
        ELSIF x = 8850 THEN
            sigmoid_f := 2021;
        ELSIF x = 8851 THEN
            sigmoid_f := 2021;
        ELSIF x = 8852 THEN
            sigmoid_f := 2021;
        ELSIF x = 8853 THEN
            sigmoid_f := 2021;
        ELSIF x = 8854 THEN
            sigmoid_f := 2021;
        ELSIF x = 8855 THEN
            sigmoid_f := 2021;
        ELSIF x = 8856 THEN
            sigmoid_f := 2021;
        ELSIF x = 8857 THEN
            sigmoid_f := 2021;
        ELSIF x = 8858 THEN
            sigmoid_f := 2021;
        ELSIF x = 8859 THEN
            sigmoid_f := 2021;
        ELSIF x = 8860 THEN
            sigmoid_f := 2021;
        ELSIF x = 8861 THEN
            sigmoid_f := 2021;
        ELSIF x = 8862 THEN
            sigmoid_f := 2021;
        ELSIF x = 8863 THEN
            sigmoid_f := 2021;
        ELSIF x = 8864 THEN
            sigmoid_f := 2021;
        ELSIF x = 8865 THEN
            sigmoid_f := 2021;
        ELSIF x = 8866 THEN
            sigmoid_f := 2021;
        ELSIF x = 8867 THEN
            sigmoid_f := 2021;
        ELSIF x = 8868 THEN
            sigmoid_f := 2021;
        ELSIF x = 8869 THEN
            sigmoid_f := 2021;
        ELSIF x = 8870 THEN
            sigmoid_f := 2021;
        ELSIF x = 8871 THEN
            sigmoid_f := 2021;
        ELSIF x = 8872 THEN
            sigmoid_f := 2021;
        ELSIF x = 8873 THEN
            sigmoid_f := 2021;
        ELSIF x = 8874 THEN
            sigmoid_f := 2021;
        ELSIF x = 8875 THEN
            sigmoid_f := 2021;
        ELSIF x = 8876 THEN
            sigmoid_f := 2021;
        ELSIF x = 8877 THEN
            sigmoid_f := 2021;
        ELSIF x = 8878 THEN
            sigmoid_f := 2021;
        ELSIF x = 8879 THEN
            sigmoid_f := 2021;
        ELSIF x = 8880 THEN
            sigmoid_f := 2021;
        ELSIF x = 8881 THEN
            sigmoid_f := 2021;
        ELSIF x = 8882 THEN
            sigmoid_f := 2021;
        ELSIF x = 8883 THEN
            sigmoid_f := 2021;
        ELSIF x = 8884 THEN
            sigmoid_f := 2021;
        ELSIF x = 8885 THEN
            sigmoid_f := 2021;
        ELSIF x = 8886 THEN
            sigmoid_f := 2021;
        ELSIF x = 8887 THEN
            sigmoid_f := 2021;
        ELSIF x = 8888 THEN
            sigmoid_f := 2021;
        ELSIF x = 8889 THEN
            sigmoid_f := 2021;
        ELSIF x = 8890 THEN
            sigmoid_f := 2021;
        ELSIF x = 8891 THEN
            sigmoid_f := 2021;
        ELSIF x = 8892 THEN
            sigmoid_f := 2021;
        ELSIF x = 8893 THEN
            sigmoid_f := 2021;
        ELSIF x = 8894 THEN
            sigmoid_f := 2021;
        ELSIF x = 8895 THEN
            sigmoid_f := 2021;
        ELSIF x = 8896 THEN
            sigmoid_f := 2021;
        ELSIF x = 8897 THEN
            sigmoid_f := 2021;
        ELSIF x = 8898 THEN
            sigmoid_f := 2021;
        ELSIF x = 8899 THEN
            sigmoid_f := 2021;
        ELSIF x = 8900 THEN
            sigmoid_f := 2021;
        ELSIF x = 8901 THEN
            sigmoid_f := 2021;
        ELSIF x = 8902 THEN
            sigmoid_f := 2021;
        ELSIF x = 8903 THEN
            sigmoid_f := 2021;
        ELSIF x = 8904 THEN
            sigmoid_f := 2021;
        ELSIF x = 8905 THEN
            sigmoid_f := 2021;
        ELSIF x = 8906 THEN
            sigmoid_f := 2021;
        ELSIF x = 8907 THEN
            sigmoid_f := 2021;
        ELSIF x = 8908 THEN
            sigmoid_f := 2021;
        ELSIF x = 8909 THEN
            sigmoid_f := 2021;
        ELSIF x = 8910 THEN
            sigmoid_f := 2021;
        ELSIF x = 8911 THEN
            sigmoid_f := 2021;
        ELSIF x = 8912 THEN
            sigmoid_f := 2021;
        ELSIF x = 8913 THEN
            sigmoid_f := 2021;
        ELSIF x = 8914 THEN
            sigmoid_f := 2021;
        ELSIF x = 8915 THEN
            sigmoid_f := 2021;
        ELSIF x = 8916 THEN
            sigmoid_f := 2021;
        ELSIF x = 8917 THEN
            sigmoid_f := 2021;
        ELSIF x = 8918 THEN
            sigmoid_f := 2021;
        ELSIF x = 8919 THEN
            sigmoid_f := 2021;
        ELSIF x = 8920 THEN
            sigmoid_f := 2021;
        ELSIF x = 8921 THEN
            sigmoid_f := 2021;
        ELSIF x = 8922 THEN
            sigmoid_f := 2021;
        ELSIF x = 8923 THEN
            sigmoid_f := 2021;
        ELSIF x = 8924 THEN
            sigmoid_f := 2021;
        ELSIF x = 8925 THEN
            sigmoid_f := 2021;
        ELSIF x = 8926 THEN
            sigmoid_f := 2021;
        ELSIF x = 8927 THEN
            sigmoid_f := 2021;
        ELSIF x = 8928 THEN
            sigmoid_f := 2021;
        ELSIF x = 8929 THEN
            sigmoid_f := 2021;
        ELSIF x = 8930 THEN
            sigmoid_f := 2022;
        ELSIF x = 8931 THEN
            sigmoid_f := 2022;
        ELSIF x = 8932 THEN
            sigmoid_f := 2022;
        ELSIF x = 8933 THEN
            sigmoid_f := 2022;
        ELSIF x = 8934 THEN
            sigmoid_f := 2022;
        ELSIF x = 8935 THEN
            sigmoid_f := 2022;
        ELSIF x = 8936 THEN
            sigmoid_f := 2022;
        ELSIF x = 8937 THEN
            sigmoid_f := 2022;
        ELSIF x = 8938 THEN
            sigmoid_f := 2022;
        ELSIF x = 8939 THEN
            sigmoid_f := 2022;
        ELSIF x = 8940 THEN
            sigmoid_f := 2022;
        ELSIF x = 8941 THEN
            sigmoid_f := 2022;
        ELSIF x = 8942 THEN
            sigmoid_f := 2022;
        ELSIF x = 8943 THEN
            sigmoid_f := 2022;
        ELSIF x = 8944 THEN
            sigmoid_f := 2022;
        ELSIF x = 8945 THEN
            sigmoid_f := 2022;
        ELSIF x = 8946 THEN
            sigmoid_f := 2022;
        ELSIF x = 8947 THEN
            sigmoid_f := 2022;
        ELSIF x = 8948 THEN
            sigmoid_f := 2022;
        ELSIF x = 8949 THEN
            sigmoid_f := 2022;
        ELSIF x = 8950 THEN
            sigmoid_f := 2022;
        ELSIF x = 8951 THEN
            sigmoid_f := 2022;
        ELSIF x = 8952 THEN
            sigmoid_f := 2022;
        ELSIF x = 8953 THEN
            sigmoid_f := 2022;
        ELSIF x = 8954 THEN
            sigmoid_f := 2022;
        ELSIF x = 8955 THEN
            sigmoid_f := 2022;
        ELSIF x = 8956 THEN
            sigmoid_f := 2022;
        ELSIF x = 8957 THEN
            sigmoid_f := 2022;
        ELSIF x = 8958 THEN
            sigmoid_f := 2022;
        ELSIF x = 8959 THEN
            sigmoid_f := 2022;
        ELSIF x = 8960 THEN
            sigmoid_f := 2022;
        ELSIF x = 8961 THEN
            sigmoid_f := 2022;
        ELSIF x = 8962 THEN
            sigmoid_f := 2022;
        ELSIF x = 8963 THEN
            sigmoid_f := 2022;
        ELSIF x = 8964 THEN
            sigmoid_f := 2022;
        ELSIF x = 8965 THEN
            sigmoid_f := 2022;
        ELSIF x = 8966 THEN
            sigmoid_f := 2022;
        ELSIF x = 8967 THEN
            sigmoid_f := 2022;
        ELSIF x = 8968 THEN
            sigmoid_f := 2022;
        ELSIF x = 8969 THEN
            sigmoid_f := 2022;
        ELSIF x = 8970 THEN
            sigmoid_f := 2022;
        ELSIF x = 8971 THEN
            sigmoid_f := 2022;
        ELSIF x = 8972 THEN
            sigmoid_f := 2022;
        ELSIF x = 8973 THEN
            sigmoid_f := 2022;
        ELSIF x = 8974 THEN
            sigmoid_f := 2022;
        ELSIF x = 8975 THEN
            sigmoid_f := 2022;
        ELSIF x = 8976 THEN
            sigmoid_f := 2022;
        ELSIF x = 8977 THEN
            sigmoid_f := 2022;
        ELSIF x = 8978 THEN
            sigmoid_f := 2022;
        ELSIF x = 8979 THEN
            sigmoid_f := 2022;
        ELSIF x = 8980 THEN
            sigmoid_f := 2022;
        ELSIF x = 8981 THEN
            sigmoid_f := 2022;
        ELSIF x = 8982 THEN
            sigmoid_f := 2022;
        ELSIF x = 8983 THEN
            sigmoid_f := 2022;
        ELSIF x = 8984 THEN
            sigmoid_f := 2022;
        ELSIF x = 8985 THEN
            sigmoid_f := 2022;
        ELSIF x = 8986 THEN
            sigmoid_f := 2022;
        ELSIF x = 8987 THEN
            sigmoid_f := 2022;
        ELSIF x = 8988 THEN
            sigmoid_f := 2022;
        ELSIF x = 8989 THEN
            sigmoid_f := 2022;
        ELSIF x = 8990 THEN
            sigmoid_f := 2022;
        ELSIF x = 8991 THEN
            sigmoid_f := 2022;
        ELSIF x = 8992 THEN
            sigmoid_f := 2022;
        ELSIF x = 8993 THEN
            sigmoid_f := 2022;
        ELSIF x = 8994 THEN
            sigmoid_f := 2022;
        ELSIF x = 8995 THEN
            sigmoid_f := 2022;
        ELSIF x = 8996 THEN
            sigmoid_f := 2022;
        ELSIF x = 8997 THEN
            sigmoid_f := 2022;
        ELSIF x = 8998 THEN
            sigmoid_f := 2022;
        ELSIF x = 8999 THEN
            sigmoid_f := 2022;
        ELSIF x = 9000 THEN
            sigmoid_f := 2022;
        ELSIF x = 9001 THEN
            sigmoid_f := 2022;
        ELSIF x = 9002 THEN
            sigmoid_f := 2022;
        ELSIF x = 9003 THEN
            sigmoid_f := 2022;
        ELSIF x = 9004 THEN
            sigmoid_f := 2022;
        ELSIF x = 9005 THEN
            sigmoid_f := 2022;
        ELSIF x = 9006 THEN
            sigmoid_f := 2022;
        ELSIF x = 9007 THEN
            sigmoid_f := 2022;
        ELSIF x = 9008 THEN
            sigmoid_f := 2022;
        ELSIF x = 9009 THEN
            sigmoid_f := 2022;
        ELSIF x = 9010 THEN
            sigmoid_f := 2022;
        ELSIF x = 9011 THEN
            sigmoid_f := 2022;
        ELSIF x = 9012 THEN
            sigmoid_f := 2023;
        ELSIF x = 9013 THEN
            sigmoid_f := 2023;
        ELSIF x = 9014 THEN
            sigmoid_f := 2023;
        ELSIF x = 9015 THEN
            sigmoid_f := 2023;
        ELSIF x = 9016 THEN
            sigmoid_f := 2023;
        ELSIF x = 9017 THEN
            sigmoid_f := 2023;
        ELSIF x = 9018 THEN
            sigmoid_f := 2023;
        ELSIF x = 9019 THEN
            sigmoid_f := 2023;
        ELSIF x = 9020 THEN
            sigmoid_f := 2023;
        ELSIF x = 9021 THEN
            sigmoid_f := 2023;
        ELSIF x = 9022 THEN
            sigmoid_f := 2023;
        ELSIF x = 9023 THEN
            sigmoid_f := 2023;
        ELSIF x = 9024 THEN
            sigmoid_f := 2023;
        ELSIF x = 9025 THEN
            sigmoid_f := 2023;
        ELSIF x = 9026 THEN
            sigmoid_f := 2023;
        ELSIF x = 9027 THEN
            sigmoid_f := 2023;
        ELSIF x = 9028 THEN
            sigmoid_f := 2023;
        ELSIF x = 9029 THEN
            sigmoid_f := 2023;
        ELSIF x = 9030 THEN
            sigmoid_f := 2023;
        ELSIF x = 9031 THEN
            sigmoid_f := 2023;
        ELSIF x = 9032 THEN
            sigmoid_f := 2023;
        ELSIF x = 9033 THEN
            sigmoid_f := 2023;
        ELSIF x = 9034 THEN
            sigmoid_f := 2023;
        ELSIF x = 9035 THEN
            sigmoid_f := 2023;
        ELSIF x = 9036 THEN
            sigmoid_f := 2023;
        ELSIF x = 9037 THEN
            sigmoid_f := 2023;
        ELSIF x = 9038 THEN
            sigmoid_f := 2023;
        ELSIF x = 9039 THEN
            sigmoid_f := 2023;
        ELSIF x = 9040 THEN
            sigmoid_f := 2023;
        ELSIF x = 9041 THEN
            sigmoid_f := 2023;
        ELSIF x = 9042 THEN
            sigmoid_f := 2023;
        ELSIF x = 9043 THEN
            sigmoid_f := 2023;
        ELSIF x = 9044 THEN
            sigmoid_f := 2023;
        ELSIF x = 9045 THEN
            sigmoid_f := 2023;
        ELSIF x = 9046 THEN
            sigmoid_f := 2023;
        ELSIF x = 9047 THEN
            sigmoid_f := 2023;
        ELSIF x = 9048 THEN
            sigmoid_f := 2023;
        ELSIF x = 9049 THEN
            sigmoid_f := 2023;
        ELSIF x = 9050 THEN
            sigmoid_f := 2023;
        ELSIF x = 9051 THEN
            sigmoid_f := 2023;
        ELSIF x = 9052 THEN
            sigmoid_f := 2023;
        ELSIF x = 9053 THEN
            sigmoid_f := 2023;
        ELSIF x = 9054 THEN
            sigmoid_f := 2023;
        ELSIF x = 9055 THEN
            sigmoid_f := 2023;
        ELSIF x = 9056 THEN
            sigmoid_f := 2023;
        ELSIF x = 9057 THEN
            sigmoid_f := 2023;
        ELSIF x = 9058 THEN
            sigmoid_f := 2023;
        ELSIF x = 9059 THEN
            sigmoid_f := 2023;
        ELSIF x = 9060 THEN
            sigmoid_f := 2023;
        ELSIF x = 9061 THEN
            sigmoid_f := 2023;
        ELSIF x = 9062 THEN
            sigmoid_f := 2023;
        ELSIF x = 9063 THEN
            sigmoid_f := 2023;
        ELSIF x = 9064 THEN
            sigmoid_f := 2023;
        ELSIF x = 9065 THEN
            sigmoid_f := 2023;
        ELSIF x = 9066 THEN
            sigmoid_f := 2023;
        ELSIF x = 9067 THEN
            sigmoid_f := 2023;
        ELSIF x = 9068 THEN
            sigmoid_f := 2023;
        ELSIF x = 9069 THEN
            sigmoid_f := 2023;
        ELSIF x = 9070 THEN
            sigmoid_f := 2023;
        ELSIF x = 9071 THEN
            sigmoid_f := 2023;
        ELSIF x = 9072 THEN
            sigmoid_f := 2023;
        ELSIF x = 9073 THEN
            sigmoid_f := 2023;
        ELSIF x = 9074 THEN
            sigmoid_f := 2023;
        ELSIF x = 9075 THEN
            sigmoid_f := 2023;
        ELSIF x = 9076 THEN
            sigmoid_f := 2023;
        ELSIF x = 9077 THEN
            sigmoid_f := 2023;
        ELSIF x = 9078 THEN
            sigmoid_f := 2023;
        ELSIF x = 9079 THEN
            sigmoid_f := 2023;
        ELSIF x = 9080 THEN
            sigmoid_f := 2023;
        ELSIF x = 9081 THEN
            sigmoid_f := 2023;
        ELSIF x = 9082 THEN
            sigmoid_f := 2023;
        ELSIF x = 9083 THEN
            sigmoid_f := 2023;
        ELSIF x = 9084 THEN
            sigmoid_f := 2023;
        ELSIF x = 9085 THEN
            sigmoid_f := 2023;
        ELSIF x = 9086 THEN
            sigmoid_f := 2023;
        ELSIF x = 9087 THEN
            sigmoid_f := 2023;
        ELSIF x = 9088 THEN
            sigmoid_f := 2023;
        ELSIF x = 9089 THEN
            sigmoid_f := 2023;
        ELSIF x = 9090 THEN
            sigmoid_f := 2023;
        ELSIF x = 9091 THEN
            sigmoid_f := 2023;
        ELSIF x = 9092 THEN
            sigmoid_f := 2023;
        ELSIF x = 9093 THEN
            sigmoid_f := 2023;
        ELSIF x = 9094 THEN
            sigmoid_f := 2024;
        ELSIF x = 9095 THEN
            sigmoid_f := 2024;
        ELSIF x = 9096 THEN
            sigmoid_f := 2024;
        ELSIF x = 9097 THEN
            sigmoid_f := 2024;
        ELSIF x = 9098 THEN
            sigmoid_f := 2024;
        ELSIF x = 9099 THEN
            sigmoid_f := 2024;
        ELSIF x = 9100 THEN
            sigmoid_f := 2024;
        ELSIF x = 9101 THEN
            sigmoid_f := 2024;
        ELSIF x = 9102 THEN
            sigmoid_f := 2024;
        ELSIF x = 9103 THEN
            sigmoid_f := 2024;
        ELSIF x = 9104 THEN
            sigmoid_f := 2024;
        ELSIF x = 9105 THEN
            sigmoid_f := 2024;
        ELSIF x = 9106 THEN
            sigmoid_f := 2024;
        ELSIF x = 9107 THEN
            sigmoid_f := 2024;
        ELSIF x = 9108 THEN
            sigmoid_f := 2024;
        ELSIF x = 9109 THEN
            sigmoid_f := 2024;
        ELSIF x = 9110 THEN
            sigmoid_f := 2024;
        ELSIF x = 9111 THEN
            sigmoid_f := 2024;
        ELSIF x = 9112 THEN
            sigmoid_f := 2024;
        ELSIF x = 9113 THEN
            sigmoid_f := 2024;
        ELSIF x = 9114 THEN
            sigmoid_f := 2024;
        ELSIF x = 9115 THEN
            sigmoid_f := 2024;
        ELSIF x = 9116 THEN
            sigmoid_f := 2024;
        ELSIF x = 9117 THEN
            sigmoid_f := 2024;
        ELSIF x = 9118 THEN
            sigmoid_f := 2024;
        ELSIF x = 9119 THEN
            sigmoid_f := 2024;
        ELSIF x = 9120 THEN
            sigmoid_f := 2024;
        ELSIF x = 9121 THEN
            sigmoid_f := 2024;
        ELSIF x = 9122 THEN
            sigmoid_f := 2024;
        ELSIF x = 9123 THEN
            sigmoid_f := 2024;
        ELSIF x = 9124 THEN
            sigmoid_f := 2024;
        ELSIF x = 9125 THEN
            sigmoid_f := 2024;
        ELSIF x = 9126 THEN
            sigmoid_f := 2024;
        ELSIF x = 9127 THEN
            sigmoid_f := 2024;
        ELSIF x = 9128 THEN
            sigmoid_f := 2024;
        ELSIF x = 9129 THEN
            sigmoid_f := 2024;
        ELSIF x = 9130 THEN
            sigmoid_f := 2024;
        ELSIF x = 9131 THEN
            sigmoid_f := 2024;
        ELSIF x = 9132 THEN
            sigmoid_f := 2024;
        ELSIF x = 9133 THEN
            sigmoid_f := 2024;
        ELSIF x = 9134 THEN
            sigmoid_f := 2024;
        ELSIF x = 9135 THEN
            sigmoid_f := 2024;
        ELSIF x = 9136 THEN
            sigmoid_f := 2024;
        ELSIF x = 9137 THEN
            sigmoid_f := 2024;
        ELSIF x = 9138 THEN
            sigmoid_f := 2024;
        ELSIF x = 9139 THEN
            sigmoid_f := 2024;
        ELSIF x = 9140 THEN
            sigmoid_f := 2024;
        ELSIF x = 9141 THEN
            sigmoid_f := 2024;
        ELSIF x = 9142 THEN
            sigmoid_f := 2024;
        ELSIF x = 9143 THEN
            sigmoid_f := 2024;
        ELSIF x = 9144 THEN
            sigmoid_f := 2024;
        ELSIF x = 9145 THEN
            sigmoid_f := 2024;
        ELSIF x = 9146 THEN
            sigmoid_f := 2024;
        ELSIF x = 9147 THEN
            sigmoid_f := 2024;
        ELSIF x = 9148 THEN
            sigmoid_f := 2024;
        ELSIF x = 9149 THEN
            sigmoid_f := 2024;
        ELSIF x = 9150 THEN
            sigmoid_f := 2024;
        ELSIF x = 9151 THEN
            sigmoid_f := 2024;
        ELSIF x = 9152 THEN
            sigmoid_f := 2024;
        ELSIF x = 9153 THEN
            sigmoid_f := 2024;
        ELSIF x = 9154 THEN
            sigmoid_f := 2024;
        ELSIF x = 9155 THEN
            sigmoid_f := 2024;
        ELSIF x = 9156 THEN
            sigmoid_f := 2024;
        ELSIF x = 9157 THEN
            sigmoid_f := 2024;
        ELSIF x = 9158 THEN
            sigmoid_f := 2024;
        ELSIF x = 9159 THEN
            sigmoid_f := 2024;
        ELSIF x = 9160 THEN
            sigmoid_f := 2024;
        ELSIF x = 9161 THEN
            sigmoid_f := 2024;
        ELSIF x = 9162 THEN
            sigmoid_f := 2024;
        ELSIF x = 9163 THEN
            sigmoid_f := 2024;
        ELSIF x = 9164 THEN
            sigmoid_f := 2024;
        ELSIF x = 9165 THEN
            sigmoid_f := 2024;
        ELSIF x = 9166 THEN
            sigmoid_f := 2024;
        ELSIF x = 9167 THEN
            sigmoid_f := 2024;
        ELSIF x = 9168 THEN
            sigmoid_f := 2024;
        ELSIF x = 9169 THEN
            sigmoid_f := 2024;
        ELSIF x = 9170 THEN
            sigmoid_f := 2024;
        ELSIF x = 9171 THEN
            sigmoid_f := 2024;
        ELSIF x = 9172 THEN
            sigmoid_f := 2024;
        ELSIF x = 9173 THEN
            sigmoid_f := 2024;
        ELSIF x = 9174 THEN
            sigmoid_f := 2024;
        ELSIF x = 9175 THEN
            sigmoid_f := 2024;
        ELSIF x = 9176 THEN
            sigmoid_f := 2025;
        ELSIF x = 9177 THEN
            sigmoid_f := 2025;
        ELSIF x = 9178 THEN
            sigmoid_f := 2025;
        ELSIF x = 9179 THEN
            sigmoid_f := 2025;
        ELSIF x = 9180 THEN
            sigmoid_f := 2025;
        ELSIF x = 9181 THEN
            sigmoid_f := 2025;
        ELSIF x = 9182 THEN
            sigmoid_f := 2025;
        ELSIF x = 9183 THEN
            sigmoid_f := 2025;
        ELSIF x = 9184 THEN
            sigmoid_f := 2025;
        ELSIF x = 9185 THEN
            sigmoid_f := 2025;
        ELSIF x = 9186 THEN
            sigmoid_f := 2025;
        ELSIF x = 9187 THEN
            sigmoid_f := 2025;
        ELSIF x = 9188 THEN
            sigmoid_f := 2025;
        ELSIF x = 9189 THEN
            sigmoid_f := 2025;
        ELSIF x = 9190 THEN
            sigmoid_f := 2025;
        ELSIF x = 9191 THEN
            sigmoid_f := 2025;
        ELSIF x = 9192 THEN
            sigmoid_f := 2025;
        ELSIF x = 9193 THEN
            sigmoid_f := 2025;
        ELSIF x = 9194 THEN
            sigmoid_f := 2025;
        ELSIF x = 9195 THEN
            sigmoid_f := 2025;
        ELSIF x = 9196 THEN
            sigmoid_f := 2025;
        ELSIF x = 9197 THEN
            sigmoid_f := 2025;
        ELSIF x = 9198 THEN
            sigmoid_f := 2025;
        ELSIF x = 9199 THEN
            sigmoid_f := 2025;
        ELSIF x = 9200 THEN
            sigmoid_f := 2025;
        ELSIF x = 9201 THEN
            sigmoid_f := 2025;
        ELSIF x = 9202 THEN
            sigmoid_f := 2025;
        ELSIF x = 9203 THEN
            sigmoid_f := 2025;
        ELSIF x = 9204 THEN
            sigmoid_f := 2025;
        ELSIF x = 9205 THEN
            sigmoid_f := 2025;
        ELSIF x = 9206 THEN
            sigmoid_f := 2025;
        ELSIF x = 9207 THEN
            sigmoid_f := 2025;
        ELSIF x = 9208 THEN
            sigmoid_f := 2025;
        ELSIF x = 9209 THEN
            sigmoid_f := 2025;
        ELSIF x = 9210 THEN
            sigmoid_f := 2025;
        ELSIF x = 9211 THEN
            sigmoid_f := 2025;
        ELSIF x = 9212 THEN
            sigmoid_f := 2025;
        ELSIF x = 9213 THEN
            sigmoid_f := 2025;
        ELSIF x = 9214 THEN
            sigmoid_f := 2025;
        ELSIF x = 9215 THEN
            sigmoid_f := 2025;
        ELSIF x = 9216 THEN
            sigmoid_f := 2025;
        ELSIF x = 9217 THEN
            sigmoid_f := 2025;
        ELSIF x = 9218 THEN
            sigmoid_f := 2025;
        ELSIF x = 9219 THEN
            sigmoid_f := 2025;
        ELSIF x = 9220 THEN
            sigmoid_f := 2025;
        ELSIF x = 9221 THEN
            sigmoid_f := 2025;
        ELSIF x = 9222 THEN
            sigmoid_f := 2025;
        ELSIF x = 9223 THEN
            sigmoid_f := 2025;
        ELSIF x = 9224 THEN
            sigmoid_f := 2025;
        ELSIF x = 9225 THEN
            sigmoid_f := 2025;
        ELSIF x = 9226 THEN
            sigmoid_f := 2025;
        ELSIF x = 9227 THEN
            sigmoid_f := 2025;
        ELSIF x = 9228 THEN
            sigmoid_f := 2025;
        ELSIF x = 9229 THEN
            sigmoid_f := 2025;
        ELSIF x = 9230 THEN
            sigmoid_f := 2025;
        ELSIF x = 9231 THEN
            sigmoid_f := 2025;
        ELSIF x = 9232 THEN
            sigmoid_f := 2025;
        ELSIF x = 9233 THEN
            sigmoid_f := 2025;
        ELSIF x = 9234 THEN
            sigmoid_f := 2025;
        ELSIF x = 9235 THEN
            sigmoid_f := 2025;
        ELSIF x = 9236 THEN
            sigmoid_f := 2025;
        ELSIF x = 9237 THEN
            sigmoid_f := 2025;
        ELSIF x = 9238 THEN
            sigmoid_f := 2025;
        ELSIF x = 9239 THEN
            sigmoid_f := 2025;
        ELSIF x = 9240 THEN
            sigmoid_f := 2025;
        ELSIF x = 9241 THEN
            sigmoid_f := 2025;
        ELSIF x = 9242 THEN
            sigmoid_f := 2025;
        ELSIF x = 9243 THEN
            sigmoid_f := 2025;
        ELSIF x = 9244 THEN
            sigmoid_f := 2025;
        ELSIF x = 9245 THEN
            sigmoid_f := 2025;
        ELSIF x = 9246 THEN
            sigmoid_f := 2025;
        ELSIF x = 9247 THEN
            sigmoid_f := 2025;
        ELSIF x = 9248 THEN
            sigmoid_f := 2025;
        ELSIF x = 9249 THEN
            sigmoid_f := 2025;
        ELSIF x = 9250 THEN
            sigmoid_f := 2025;
        ELSIF x = 9251 THEN
            sigmoid_f := 2025;
        ELSIF x = 9252 THEN
            sigmoid_f := 2025;
        ELSIF x = 9253 THEN
            sigmoid_f := 2025;
        ELSIF x = 9254 THEN
            sigmoid_f := 2025;
        ELSIF x = 9255 THEN
            sigmoid_f := 2025;
        ELSIF x = 9256 THEN
            sigmoid_f := 2025;
        ELSIF x = 9257 THEN
            sigmoid_f := 2025;
        ELSIF x = 9258 THEN
            sigmoid_f := 2025;
        ELSIF x = 9259 THEN
            sigmoid_f := 2025;
        ELSIF x = 9260 THEN
            sigmoid_f := 2025;
        ELSIF x = 9261 THEN
            sigmoid_f := 2025;
        ELSIF x = 9262 THEN
            sigmoid_f := 2025;
        ELSIF x = 9263 THEN
            sigmoid_f := 2025;
        ELSIF x = 9264 THEN
            sigmoid_f := 2025;
        ELSIF x = 9265 THEN
            sigmoid_f := 2026;
        ELSIF x = 9266 THEN
            sigmoid_f := 2026;
        ELSIF x = 9267 THEN
            sigmoid_f := 2026;
        ELSIF x = 9268 THEN
            sigmoid_f := 2026;
        ELSIF x = 9269 THEN
            sigmoid_f := 2026;
        ELSIF x = 9270 THEN
            sigmoid_f := 2026;
        ELSIF x = 9271 THEN
            sigmoid_f := 2026;
        ELSIF x = 9272 THEN
            sigmoid_f := 2026;
        ELSIF x = 9273 THEN
            sigmoid_f := 2026;
        ELSIF x = 9274 THEN
            sigmoid_f := 2026;
        ELSIF x = 9275 THEN
            sigmoid_f := 2026;
        ELSIF x = 9276 THEN
            sigmoid_f := 2026;
        ELSIF x = 9277 THEN
            sigmoid_f := 2026;
        ELSIF x = 9278 THEN
            sigmoid_f := 2026;
        ELSIF x = 9279 THEN
            sigmoid_f := 2026;
        ELSIF x = 9280 THEN
            sigmoid_f := 2026;
        ELSIF x = 9281 THEN
            sigmoid_f := 2026;
        ELSIF x = 9282 THEN
            sigmoid_f := 2026;
        ELSIF x = 9283 THEN
            sigmoid_f := 2026;
        ELSIF x = 9284 THEN
            sigmoid_f := 2026;
        ELSIF x = 9285 THEN
            sigmoid_f := 2026;
        ELSIF x = 9286 THEN
            sigmoid_f := 2026;
        ELSIF x = 9287 THEN
            sigmoid_f := 2026;
        ELSIF x = 9288 THEN
            sigmoid_f := 2026;
        ELSIF x = 9289 THEN
            sigmoid_f := 2026;
        ELSIF x = 9290 THEN
            sigmoid_f := 2026;
        ELSIF x = 9291 THEN
            sigmoid_f := 2026;
        ELSIF x = 9292 THEN
            sigmoid_f := 2026;
        ELSIF x = 9293 THEN
            sigmoid_f := 2026;
        ELSIF x = 9294 THEN
            sigmoid_f := 2026;
        ELSIF x = 9295 THEN
            sigmoid_f := 2026;
        ELSIF x = 9296 THEN
            sigmoid_f := 2026;
        ELSIF x = 9297 THEN
            sigmoid_f := 2026;
        ELSIF x = 9298 THEN
            sigmoid_f := 2026;
        ELSIF x = 9299 THEN
            sigmoid_f := 2026;
        ELSIF x = 9300 THEN
            sigmoid_f := 2026;
        ELSIF x = 9301 THEN
            sigmoid_f := 2026;
        ELSIF x = 9302 THEN
            sigmoid_f := 2026;
        ELSIF x = 9303 THEN
            sigmoid_f := 2026;
        ELSIF x = 9304 THEN
            sigmoid_f := 2026;
        ELSIF x = 9305 THEN
            sigmoid_f := 2026;
        ELSIF x = 9306 THEN
            sigmoid_f := 2026;
        ELSIF x = 9307 THEN
            sigmoid_f := 2026;
        ELSIF x = 9308 THEN
            sigmoid_f := 2026;
        ELSIF x = 9309 THEN
            sigmoid_f := 2026;
        ELSIF x = 9310 THEN
            sigmoid_f := 2026;
        ELSIF x = 9311 THEN
            sigmoid_f := 2026;
        ELSIF x = 9312 THEN
            sigmoid_f := 2026;
        ELSIF x = 9313 THEN
            sigmoid_f := 2026;
        ELSIF x = 9314 THEN
            sigmoid_f := 2026;
        ELSIF x = 9315 THEN
            sigmoid_f := 2026;
        ELSIF x = 9316 THEN
            sigmoid_f := 2026;
        ELSIF x = 9317 THEN
            sigmoid_f := 2026;
        ELSIF x = 9318 THEN
            sigmoid_f := 2026;
        ELSIF x = 9319 THEN
            sigmoid_f := 2026;
        ELSIF x = 9320 THEN
            sigmoid_f := 2026;
        ELSIF x = 9321 THEN
            sigmoid_f := 2026;
        ELSIF x = 9322 THEN
            sigmoid_f := 2026;
        ELSIF x = 9323 THEN
            sigmoid_f := 2026;
        ELSIF x = 9324 THEN
            sigmoid_f := 2026;
        ELSIF x = 9325 THEN
            sigmoid_f := 2026;
        ELSIF x = 9326 THEN
            sigmoid_f := 2026;
        ELSIF x = 9327 THEN
            sigmoid_f := 2026;
        ELSIF x = 9328 THEN
            sigmoid_f := 2026;
        ELSIF x = 9329 THEN
            sigmoid_f := 2026;
        ELSIF x = 9330 THEN
            sigmoid_f := 2026;
        ELSIF x = 9331 THEN
            sigmoid_f := 2026;
        ELSIF x = 9332 THEN
            sigmoid_f := 2026;
        ELSIF x = 9333 THEN
            sigmoid_f := 2026;
        ELSIF x = 9334 THEN
            sigmoid_f := 2026;
        ELSIF x = 9335 THEN
            sigmoid_f := 2026;
        ELSIF x = 9336 THEN
            sigmoid_f := 2026;
        ELSIF x = 9337 THEN
            sigmoid_f := 2026;
        ELSIF x = 9338 THEN
            sigmoid_f := 2026;
        ELSIF x = 9339 THEN
            sigmoid_f := 2026;
        ELSIF x = 9340 THEN
            sigmoid_f := 2026;
        ELSIF x = 9341 THEN
            sigmoid_f := 2026;
        ELSIF x = 9342 THEN
            sigmoid_f := 2026;
        ELSIF x = 9343 THEN
            sigmoid_f := 2026;
        ELSIF x = 9344 THEN
            sigmoid_f := 2026;
        ELSIF x = 9345 THEN
            sigmoid_f := 2026;
        ELSIF x = 9346 THEN
            sigmoid_f := 2026;
        ELSIF x = 9347 THEN
            sigmoid_f := 2026;
        ELSIF x = 9348 THEN
            sigmoid_f := 2026;
        ELSIF x = 9349 THEN
            sigmoid_f := 2026;
        ELSIF x = 9350 THEN
            sigmoid_f := 2026;
        ELSIF x = 9351 THEN
            sigmoid_f := 2026;
        ELSIF x = 9352 THEN
            sigmoid_f := 2026;
        ELSIF x = 9353 THEN
            sigmoid_f := 2026;
        ELSIF x = 9354 THEN
            sigmoid_f := 2026;
        ELSIF x = 9355 THEN
            sigmoid_f := 2026;
        ELSIF x = 9356 THEN
            sigmoid_f := 2026;
        ELSIF x = 9357 THEN
            sigmoid_f := 2026;
        ELSIF x = 9358 THEN
            sigmoid_f := 2026;
        ELSIF x = 9359 THEN
            sigmoid_f := 2026;
        ELSIF x = 9360 THEN
            sigmoid_f := 2026;
        ELSIF x = 9361 THEN
            sigmoid_f := 2026;
        ELSIF x = 9362 THEN
            sigmoid_f := 2026;
        ELSIF x = 9363 THEN
            sigmoid_f := 2027;
        ELSIF x = 9364 THEN
            sigmoid_f := 2027;
        ELSIF x = 9365 THEN
            sigmoid_f := 2027;
        ELSIF x = 9366 THEN
            sigmoid_f := 2027;
        ELSIF x = 9367 THEN
            sigmoid_f := 2027;
        ELSIF x = 9368 THEN
            sigmoid_f := 2027;
        ELSIF x = 9369 THEN
            sigmoid_f := 2027;
        ELSIF x = 9370 THEN
            sigmoid_f := 2027;
        ELSIF x = 9371 THEN
            sigmoid_f := 2027;
        ELSIF x = 9372 THEN
            sigmoid_f := 2027;
        ELSIF x = 9373 THEN
            sigmoid_f := 2027;
        ELSIF x = 9374 THEN
            sigmoid_f := 2027;
        ELSIF x = 9375 THEN
            sigmoid_f := 2027;
        ELSIF x = 9376 THEN
            sigmoid_f := 2027;
        ELSIF x = 9377 THEN
            sigmoid_f := 2027;
        ELSIF x = 9378 THEN
            sigmoid_f := 2027;
        ELSIF x = 9379 THEN
            sigmoid_f := 2027;
        ELSIF x = 9380 THEN
            sigmoid_f := 2027;
        ELSIF x = 9381 THEN
            sigmoid_f := 2027;
        ELSIF x = 9382 THEN
            sigmoid_f := 2027;
        ELSIF x = 9383 THEN
            sigmoid_f := 2027;
        ELSIF x = 9384 THEN
            sigmoid_f := 2027;
        ELSIF x = 9385 THEN
            sigmoid_f := 2027;
        ELSIF x = 9386 THEN
            sigmoid_f := 2027;
        ELSIF x = 9387 THEN
            sigmoid_f := 2027;
        ELSIF x = 9388 THEN
            sigmoid_f := 2027;
        ELSIF x = 9389 THEN
            sigmoid_f := 2027;
        ELSIF x = 9390 THEN
            sigmoid_f := 2027;
        ELSIF x = 9391 THEN
            sigmoid_f := 2027;
        ELSIF x = 9392 THEN
            sigmoid_f := 2027;
        ELSIF x = 9393 THEN
            sigmoid_f := 2027;
        ELSIF x = 9394 THEN
            sigmoid_f := 2027;
        ELSIF x = 9395 THEN
            sigmoid_f := 2027;
        ELSIF x = 9396 THEN
            sigmoid_f := 2027;
        ELSIF x = 9397 THEN
            sigmoid_f := 2027;
        ELSIF x = 9398 THEN
            sigmoid_f := 2027;
        ELSIF x = 9399 THEN
            sigmoid_f := 2027;
        ELSIF x = 9400 THEN
            sigmoid_f := 2027;
        ELSIF x = 9401 THEN
            sigmoid_f := 2027;
        ELSIF x = 9402 THEN
            sigmoid_f := 2027;
        ELSIF x = 9403 THEN
            sigmoid_f := 2027;
        ELSIF x = 9404 THEN
            sigmoid_f := 2027;
        ELSIF x = 9405 THEN
            sigmoid_f := 2027;
        ELSIF x = 9406 THEN
            sigmoid_f := 2027;
        ELSIF x = 9407 THEN
            sigmoid_f := 2027;
        ELSIF x = 9408 THEN
            sigmoid_f := 2027;
        ELSIF x = 9409 THEN
            sigmoid_f := 2027;
        ELSIF x = 9410 THEN
            sigmoid_f := 2027;
        ELSIF x = 9411 THEN
            sigmoid_f := 2027;
        ELSIF x = 9412 THEN
            sigmoid_f := 2027;
        ELSIF x = 9413 THEN
            sigmoid_f := 2027;
        ELSIF x = 9414 THEN
            sigmoid_f := 2027;
        ELSIF x = 9415 THEN
            sigmoid_f := 2027;
        ELSIF x = 9416 THEN
            sigmoid_f := 2027;
        ELSIF x = 9417 THEN
            sigmoid_f := 2027;
        ELSIF x = 9418 THEN
            sigmoid_f := 2027;
        ELSIF x = 9419 THEN
            sigmoid_f := 2027;
        ELSIF x = 9420 THEN
            sigmoid_f := 2027;
        ELSIF x = 9421 THEN
            sigmoid_f := 2027;
        ELSIF x = 9422 THEN
            sigmoid_f := 2027;
        ELSIF x = 9423 THEN
            sigmoid_f := 2027;
        ELSIF x = 9424 THEN
            sigmoid_f := 2027;
        ELSIF x = 9425 THEN
            sigmoid_f := 2027;
        ELSIF x = 9426 THEN
            sigmoid_f := 2027;
        ELSIF x = 9427 THEN
            sigmoid_f := 2027;
        ELSIF x = 9428 THEN
            sigmoid_f := 2027;
        ELSIF x = 9429 THEN
            sigmoid_f := 2027;
        ELSIF x = 9430 THEN
            sigmoid_f := 2027;
        ELSIF x = 9431 THEN
            sigmoid_f := 2027;
        ELSIF x = 9432 THEN
            sigmoid_f := 2027;
        ELSIF x = 9433 THEN
            sigmoid_f := 2027;
        ELSIF x = 9434 THEN
            sigmoid_f := 2027;
        ELSIF x = 9435 THEN
            sigmoid_f := 2027;
        ELSIF x = 9436 THEN
            sigmoid_f := 2027;
        ELSIF x = 9437 THEN
            sigmoid_f := 2027;
        ELSIF x = 9438 THEN
            sigmoid_f := 2027;
        ELSIF x = 9439 THEN
            sigmoid_f := 2027;
        ELSIF x = 9440 THEN
            sigmoid_f := 2027;
        ELSIF x = 9441 THEN
            sigmoid_f := 2027;
        ELSIF x = 9442 THEN
            sigmoid_f := 2027;
        ELSIF x = 9443 THEN
            sigmoid_f := 2027;
        ELSIF x = 9444 THEN
            sigmoid_f := 2027;
        ELSIF x = 9445 THEN
            sigmoid_f := 2027;
        ELSIF x = 9446 THEN
            sigmoid_f := 2027;
        ELSIF x = 9447 THEN
            sigmoid_f := 2027;
        ELSIF x = 9448 THEN
            sigmoid_f := 2027;
        ELSIF x = 9449 THEN
            sigmoid_f := 2027;
        ELSIF x = 9450 THEN
            sigmoid_f := 2027;
        ELSIF x = 9451 THEN
            sigmoid_f := 2027;
        ELSIF x = 9452 THEN
            sigmoid_f := 2027;
        ELSIF x = 9453 THEN
            sigmoid_f := 2027;
        ELSIF x = 9454 THEN
            sigmoid_f := 2027;
        ELSIF x = 9455 THEN
            sigmoid_f := 2027;
        ELSIF x = 9456 THEN
            sigmoid_f := 2027;
        ELSIF x = 9457 THEN
            sigmoid_f := 2027;
        ELSIF x = 9458 THEN
            sigmoid_f := 2027;
        ELSIF x = 9459 THEN
            sigmoid_f := 2027;
        ELSIF x = 9460 THEN
            sigmoid_f := 2028;
        ELSIF x = 9461 THEN
            sigmoid_f := 2028;
        ELSIF x = 9462 THEN
            sigmoid_f := 2028;
        ELSIF x = 9463 THEN
            sigmoid_f := 2028;
        ELSIF x = 9464 THEN
            sigmoid_f := 2028;
        ELSIF x = 9465 THEN
            sigmoid_f := 2028;
        ELSIF x = 9466 THEN
            sigmoid_f := 2028;
        ELSIF x = 9467 THEN
            sigmoid_f := 2028;
        ELSIF x = 9468 THEN
            sigmoid_f := 2028;
        ELSIF x = 9469 THEN
            sigmoid_f := 2028;
        ELSIF x = 9470 THEN
            sigmoid_f := 2028;
        ELSIF x = 9471 THEN
            sigmoid_f := 2028;
        ELSIF x = 9472 THEN
            sigmoid_f := 2028;
        ELSIF x = 9473 THEN
            sigmoid_f := 2028;
        ELSIF x = 9474 THEN
            sigmoid_f := 2028;
        ELSIF x = 9475 THEN
            sigmoid_f := 2028;
        ELSIF x = 9476 THEN
            sigmoid_f := 2028;
        ELSIF x = 9477 THEN
            sigmoid_f := 2028;
        ELSIF x = 9478 THEN
            sigmoid_f := 2028;
        ELSIF x = 9479 THEN
            sigmoid_f := 2028;
        ELSIF x = 9480 THEN
            sigmoid_f := 2028;
        ELSIF x = 9481 THEN
            sigmoid_f := 2028;
        ELSIF x = 9482 THEN
            sigmoid_f := 2028;
        ELSIF x = 9483 THEN
            sigmoid_f := 2028;
        ELSIF x = 9484 THEN
            sigmoid_f := 2028;
        ELSIF x = 9485 THEN
            sigmoid_f := 2028;
        ELSIF x = 9486 THEN
            sigmoid_f := 2028;
        ELSIF x = 9487 THEN
            sigmoid_f := 2028;
        ELSIF x = 9488 THEN
            sigmoid_f := 2028;
        ELSIF x = 9489 THEN
            sigmoid_f := 2028;
        ELSIF x = 9490 THEN
            sigmoid_f := 2028;
        ELSIF x = 9491 THEN
            sigmoid_f := 2028;
        ELSIF x = 9492 THEN
            sigmoid_f := 2028;
        ELSIF x = 9493 THEN
            sigmoid_f := 2028;
        ELSIF x = 9494 THEN
            sigmoid_f := 2028;
        ELSIF x = 9495 THEN
            sigmoid_f := 2028;
        ELSIF x = 9496 THEN
            sigmoid_f := 2028;
        ELSIF x = 9497 THEN
            sigmoid_f := 2028;
        ELSIF x = 9498 THEN
            sigmoid_f := 2028;
        ELSIF x = 9499 THEN
            sigmoid_f := 2028;
        ELSIF x = 9500 THEN
            sigmoid_f := 2028;
        ELSIF x = 9501 THEN
            sigmoid_f := 2028;
        ELSIF x = 9502 THEN
            sigmoid_f := 2028;
        ELSIF x = 9503 THEN
            sigmoid_f := 2028;
        ELSIF x = 9504 THEN
            sigmoid_f := 2028;
        ELSIF x = 9505 THEN
            sigmoid_f := 2028;
        ELSIF x = 9506 THEN
            sigmoid_f := 2028;
        ELSIF x = 9507 THEN
            sigmoid_f := 2028;
        ELSIF x = 9508 THEN
            sigmoid_f := 2028;
        ELSIF x = 9509 THEN
            sigmoid_f := 2028;
        ELSIF x = 9510 THEN
            sigmoid_f := 2028;
        ELSIF x = 9511 THEN
            sigmoid_f := 2028;
        ELSIF x = 9512 THEN
            sigmoid_f := 2028;
        ELSIF x = 9513 THEN
            sigmoid_f := 2028;
        ELSIF x = 9514 THEN
            sigmoid_f := 2028;
        ELSIF x = 9515 THEN
            sigmoid_f := 2028;
        ELSIF x = 9516 THEN
            sigmoid_f := 2028;
        ELSIF x = 9517 THEN
            sigmoid_f := 2028;
        ELSIF x = 9518 THEN
            sigmoid_f := 2028;
        ELSIF x = 9519 THEN
            sigmoid_f := 2028;
        ELSIF x = 9520 THEN
            sigmoid_f := 2028;
        ELSIF x = 9521 THEN
            sigmoid_f := 2028;
        ELSIF x = 9522 THEN
            sigmoid_f := 2028;
        ELSIF x = 9523 THEN
            sigmoid_f := 2028;
        ELSIF x = 9524 THEN
            sigmoid_f := 2028;
        ELSIF x = 9525 THEN
            sigmoid_f := 2028;
        ELSIF x = 9526 THEN
            sigmoid_f := 2028;
        ELSIF x = 9527 THEN
            sigmoid_f := 2028;
        ELSIF x = 9528 THEN
            sigmoid_f := 2028;
        ELSIF x = 9529 THEN
            sigmoid_f := 2028;
        ELSIF x = 9530 THEN
            sigmoid_f := 2028;
        ELSIF x = 9531 THEN
            sigmoid_f := 2028;
        ELSIF x = 9532 THEN
            sigmoid_f := 2028;
        ELSIF x = 9533 THEN
            sigmoid_f := 2028;
        ELSIF x = 9534 THEN
            sigmoid_f := 2028;
        ELSIF x = 9535 THEN
            sigmoid_f := 2028;
        ELSIF x = 9536 THEN
            sigmoid_f := 2028;
        ELSIF x = 9537 THEN
            sigmoid_f := 2028;
        ELSIF x = 9538 THEN
            sigmoid_f := 2028;
        ELSIF x = 9539 THEN
            sigmoid_f := 2028;
        ELSIF x = 9540 THEN
            sigmoid_f := 2028;
        ELSIF x = 9541 THEN
            sigmoid_f := 2028;
        ELSIF x = 9542 THEN
            sigmoid_f := 2028;
        ELSIF x = 9543 THEN
            sigmoid_f := 2028;
        ELSIF x = 9544 THEN
            sigmoid_f := 2028;
        ELSIF x = 9545 THEN
            sigmoid_f := 2028;
        ELSIF x = 9546 THEN
            sigmoid_f := 2028;
        ELSIF x = 9547 THEN
            sigmoid_f := 2028;
        ELSIF x = 9548 THEN
            sigmoid_f := 2028;
        ELSIF x = 9549 THEN
            sigmoid_f := 2028;
        ELSIF x = 9550 THEN
            sigmoid_f := 2028;
        ELSIF x = 9551 THEN
            sigmoid_f := 2028;
        ELSIF x = 9552 THEN
            sigmoid_f := 2028;
        ELSIF x = 9553 THEN
            sigmoid_f := 2028;
        ELSIF x = 9554 THEN
            sigmoid_f := 2028;
        ELSIF x = 9555 THEN
            sigmoid_f := 2028;
        ELSIF x = 9556 THEN
            sigmoid_f := 2028;
        ELSIF x = 9557 THEN
            sigmoid_f := 2028;
        ELSIF x = 9558 THEN
            sigmoid_f := 2029;
        ELSIF x = 9559 THEN
            sigmoid_f := 2029;
        ELSIF x = 9560 THEN
            sigmoid_f := 2029;
        ELSIF x = 9561 THEN
            sigmoid_f := 2029;
        ELSIF x = 9562 THEN
            sigmoid_f := 2029;
        ELSIF x = 9563 THEN
            sigmoid_f := 2029;
        ELSIF x = 9564 THEN
            sigmoid_f := 2029;
        ELSIF x = 9565 THEN
            sigmoid_f := 2029;
        ELSIF x = 9566 THEN
            sigmoid_f := 2029;
        ELSIF x = 9567 THEN
            sigmoid_f := 2029;
        ELSIF x = 9568 THEN
            sigmoid_f := 2029;
        ELSIF x = 9569 THEN
            sigmoid_f := 2029;
        ELSIF x = 9570 THEN
            sigmoid_f := 2029;
        ELSIF x = 9571 THEN
            sigmoid_f := 2029;
        ELSIF x = 9572 THEN
            sigmoid_f := 2029;
        ELSIF x = 9573 THEN
            sigmoid_f := 2029;
        ELSIF x = 9574 THEN
            sigmoid_f := 2029;
        ELSIF x = 9575 THEN
            sigmoid_f := 2029;
        ELSIF x = 9576 THEN
            sigmoid_f := 2029;
        ELSIF x = 9577 THEN
            sigmoid_f := 2029;
        ELSIF x = 9578 THEN
            sigmoid_f := 2029;
        ELSIF x = 9579 THEN
            sigmoid_f := 2029;
        ELSIF x = 9580 THEN
            sigmoid_f := 2029;
        ELSIF x = 9581 THEN
            sigmoid_f := 2029;
        ELSIF x = 9582 THEN
            sigmoid_f := 2029;
        ELSIF x = 9583 THEN
            sigmoid_f := 2029;
        ELSIF x = 9584 THEN
            sigmoid_f := 2029;
        ELSIF x = 9585 THEN
            sigmoid_f := 2029;
        ELSIF x = 9586 THEN
            sigmoid_f := 2029;
        ELSIF x = 9587 THEN
            sigmoid_f := 2029;
        ELSIF x = 9588 THEN
            sigmoid_f := 2029;
        ELSIF x = 9589 THEN
            sigmoid_f := 2029;
        ELSIF x = 9590 THEN
            sigmoid_f := 2029;
        ELSIF x = 9591 THEN
            sigmoid_f := 2029;
        ELSIF x = 9592 THEN
            sigmoid_f := 2029;
        ELSIF x = 9593 THEN
            sigmoid_f := 2029;
        ELSIF x = 9594 THEN
            sigmoid_f := 2029;
        ELSIF x = 9595 THEN
            sigmoid_f := 2029;
        ELSIF x = 9596 THEN
            sigmoid_f := 2029;
        ELSIF x = 9597 THEN
            sigmoid_f := 2029;
        ELSIF x = 9598 THEN
            sigmoid_f := 2029;
        ELSIF x = 9599 THEN
            sigmoid_f := 2029;
        ELSIF x = 9600 THEN
            sigmoid_f := 2029;
        ELSIF x = 9601 THEN
            sigmoid_f := 2029;
        ELSIF x = 9602 THEN
            sigmoid_f := 2029;
        ELSIF x = 9603 THEN
            sigmoid_f := 2029;
        ELSIF x = 9604 THEN
            sigmoid_f := 2029;
        ELSIF x = 9605 THEN
            sigmoid_f := 2029;
        ELSIF x = 9606 THEN
            sigmoid_f := 2029;
        ELSIF x = 9607 THEN
            sigmoid_f := 2029;
        ELSIF x = 9608 THEN
            sigmoid_f := 2029;
        ELSIF x = 9609 THEN
            sigmoid_f := 2029;
        ELSIF x = 9610 THEN
            sigmoid_f := 2029;
        ELSIF x = 9611 THEN
            sigmoid_f := 2029;
        ELSIF x = 9612 THEN
            sigmoid_f := 2029;
        ELSIF x = 9613 THEN
            sigmoid_f := 2029;
        ELSIF x = 9614 THEN
            sigmoid_f := 2029;
        ELSIF x = 9615 THEN
            sigmoid_f := 2029;
        ELSIF x = 9616 THEN
            sigmoid_f := 2029;
        ELSIF x = 9617 THEN
            sigmoid_f := 2029;
        ELSIF x = 9618 THEN
            sigmoid_f := 2029;
        ELSIF x = 9619 THEN
            sigmoid_f := 2029;
        ELSIF x = 9620 THEN
            sigmoid_f := 2029;
        ELSIF x = 9621 THEN
            sigmoid_f := 2029;
        ELSIF x = 9622 THEN
            sigmoid_f := 2029;
        ELSIF x = 9623 THEN
            sigmoid_f := 2029;
        ELSIF x = 9624 THEN
            sigmoid_f := 2029;
        ELSIF x = 9625 THEN
            sigmoid_f := 2029;
        ELSIF x = 9626 THEN
            sigmoid_f := 2029;
        ELSIF x = 9627 THEN
            sigmoid_f := 2029;
        ELSIF x = 9628 THEN
            sigmoid_f := 2029;
        ELSIF x = 9629 THEN
            sigmoid_f := 2029;
        ELSIF x = 9630 THEN
            sigmoid_f := 2029;
        ELSIF x = 9631 THEN
            sigmoid_f := 2029;
        ELSIF x = 9632 THEN
            sigmoid_f := 2029;
        ELSIF x = 9633 THEN
            sigmoid_f := 2029;
        ELSIF x = 9634 THEN
            sigmoid_f := 2029;
        ELSIF x = 9635 THEN
            sigmoid_f := 2029;
        ELSIF x = 9636 THEN
            sigmoid_f := 2029;
        ELSIF x = 9637 THEN
            sigmoid_f := 2029;
        ELSIF x = 9638 THEN
            sigmoid_f := 2029;
        ELSIF x = 9639 THEN
            sigmoid_f := 2029;
        ELSIF x = 9640 THEN
            sigmoid_f := 2029;
        ELSIF x = 9641 THEN
            sigmoid_f := 2029;
        ELSIF x = 9642 THEN
            sigmoid_f := 2029;
        ELSIF x = 9643 THEN
            sigmoid_f := 2029;
        ELSIF x = 9644 THEN
            sigmoid_f := 2029;
        ELSIF x = 9645 THEN
            sigmoid_f := 2029;
        ELSIF x = 9646 THEN
            sigmoid_f := 2029;
        ELSIF x = 9647 THEN
            sigmoid_f := 2029;
        ELSIF x = 9648 THEN
            sigmoid_f := 2029;
        ELSIF x = 9649 THEN
            sigmoid_f := 2029;
        ELSIF x = 9650 THEN
            sigmoid_f := 2029;
        ELSIF x = 9651 THEN
            sigmoid_f := 2029;
        ELSIF x = 9652 THEN
            sigmoid_f := 2029;
        ELSIF x = 9653 THEN
            sigmoid_f := 2029;
        ELSIF x = 9654 THEN
            sigmoid_f := 2029;
        ELSIF x = 9655 THEN
            sigmoid_f := 2030;
        ELSIF x = 9656 THEN
            sigmoid_f := 2030;
        ELSIF x = 9657 THEN
            sigmoid_f := 2030;
        ELSIF x = 9658 THEN
            sigmoid_f := 2030;
        ELSIF x = 9659 THEN
            sigmoid_f := 2030;
        ELSIF x = 9660 THEN
            sigmoid_f := 2030;
        ELSIF x = 9661 THEN
            sigmoid_f := 2030;
        ELSIF x = 9662 THEN
            sigmoid_f := 2030;
        ELSIF x = 9663 THEN
            sigmoid_f := 2030;
        ELSIF x = 9664 THEN
            sigmoid_f := 2030;
        ELSIF x = 9665 THEN
            sigmoid_f := 2030;
        ELSIF x = 9666 THEN
            sigmoid_f := 2030;
        ELSIF x = 9667 THEN
            sigmoid_f := 2030;
        ELSIF x = 9668 THEN
            sigmoid_f := 2030;
        ELSIF x = 9669 THEN
            sigmoid_f := 2030;
        ELSIF x = 9670 THEN
            sigmoid_f := 2030;
        ELSIF x = 9671 THEN
            sigmoid_f := 2030;
        ELSIF x = 9672 THEN
            sigmoid_f := 2030;
        ELSIF x = 9673 THEN
            sigmoid_f := 2030;
        ELSIF x = 9674 THEN
            sigmoid_f := 2030;
        ELSIF x = 9675 THEN
            sigmoid_f := 2030;
        ELSIF x = 9676 THEN
            sigmoid_f := 2030;
        ELSIF x = 9677 THEN
            sigmoid_f := 2030;
        ELSIF x = 9678 THEN
            sigmoid_f := 2030;
        ELSIF x = 9679 THEN
            sigmoid_f := 2030;
        ELSIF x = 9680 THEN
            sigmoid_f := 2030;
        ELSIF x = 9681 THEN
            sigmoid_f := 2030;
        ELSIF x = 9682 THEN
            sigmoid_f := 2030;
        ELSIF x = 9683 THEN
            sigmoid_f := 2030;
        ELSIF x = 9684 THEN
            sigmoid_f := 2030;
        ELSIF x = 9685 THEN
            sigmoid_f := 2030;
        ELSIF x = 9686 THEN
            sigmoid_f := 2030;
        ELSIF x = 9687 THEN
            sigmoid_f := 2030;
        ELSIF x = 9688 THEN
            sigmoid_f := 2030;
        ELSIF x = 9689 THEN
            sigmoid_f := 2030;
        ELSIF x = 9690 THEN
            sigmoid_f := 2030;
        ELSIF x = 9691 THEN
            sigmoid_f := 2030;
        ELSIF x = 9692 THEN
            sigmoid_f := 2030;
        ELSIF x = 9693 THEN
            sigmoid_f := 2030;
        ELSIF x = 9694 THEN
            sigmoid_f := 2030;
        ELSIF x = 9695 THEN
            sigmoid_f := 2030;
        ELSIF x = 9696 THEN
            sigmoid_f := 2030;
        ELSIF x = 9697 THEN
            sigmoid_f := 2030;
        ELSIF x = 9698 THEN
            sigmoid_f := 2030;
        ELSIF x = 9699 THEN
            sigmoid_f := 2030;
        ELSIF x = 9700 THEN
            sigmoid_f := 2030;
        ELSIF x = 9701 THEN
            sigmoid_f := 2030;
        ELSIF x = 9702 THEN
            sigmoid_f := 2030;
        ELSIF x = 9703 THEN
            sigmoid_f := 2030;
        ELSIF x = 9704 THEN
            sigmoid_f := 2030;
        ELSIF x = 9705 THEN
            sigmoid_f := 2030;
        ELSIF x = 9706 THEN
            sigmoid_f := 2030;
        ELSIF x = 9707 THEN
            sigmoid_f := 2030;
        ELSIF x = 9708 THEN
            sigmoid_f := 2030;
        ELSIF x = 9709 THEN
            sigmoid_f := 2030;
        ELSIF x = 9710 THEN
            sigmoid_f := 2030;
        ELSIF x = 9711 THEN
            sigmoid_f := 2030;
        ELSIF x = 9712 THEN
            sigmoid_f := 2030;
        ELSIF x = 9713 THEN
            sigmoid_f := 2030;
        ELSIF x = 9714 THEN
            sigmoid_f := 2030;
        ELSIF x = 9715 THEN
            sigmoid_f := 2030;
        ELSIF x = 9716 THEN
            sigmoid_f := 2030;
        ELSIF x = 9717 THEN
            sigmoid_f := 2030;
        ELSIF x = 9718 THEN
            sigmoid_f := 2030;
        ELSIF x = 9719 THEN
            sigmoid_f := 2030;
        ELSIF x = 9720 THEN
            sigmoid_f := 2030;
        ELSIF x = 9721 THEN
            sigmoid_f := 2030;
        ELSIF x = 9722 THEN
            sigmoid_f := 2030;
        ELSIF x = 9723 THEN
            sigmoid_f := 2030;
        ELSIF x = 9724 THEN
            sigmoid_f := 2030;
        ELSIF x = 9725 THEN
            sigmoid_f := 2030;
        ELSIF x = 9726 THEN
            sigmoid_f := 2030;
        ELSIF x = 9727 THEN
            sigmoid_f := 2030;
        ELSIF x = 9728 THEN
            sigmoid_f := 2030;
        ELSIF x = 9729 THEN
            sigmoid_f := 2030;
        ELSIF x = 9730 THEN
            sigmoid_f := 2030;
        ELSIF x = 9731 THEN
            sigmoid_f := 2030;
        ELSIF x = 9732 THEN
            sigmoid_f := 2030;
        ELSIF x = 9733 THEN
            sigmoid_f := 2030;
        ELSIF x = 9734 THEN
            sigmoid_f := 2030;
        ELSIF x = 9735 THEN
            sigmoid_f := 2030;
        ELSIF x = 9736 THEN
            sigmoid_f := 2030;
        ELSIF x = 9737 THEN
            sigmoid_f := 2030;
        ELSIF x = 9738 THEN
            sigmoid_f := 2030;
        ELSIF x = 9739 THEN
            sigmoid_f := 2030;
        ELSIF x = 9740 THEN
            sigmoid_f := 2030;
        ELSIF x = 9741 THEN
            sigmoid_f := 2030;
        ELSIF x = 9742 THEN
            sigmoid_f := 2030;
        ELSIF x = 9743 THEN
            sigmoid_f := 2030;
        ELSIF x = 9744 THEN
            sigmoid_f := 2030;
        ELSIF x = 9745 THEN
            sigmoid_f := 2030;
        ELSIF x = 9746 THEN
            sigmoid_f := 2030;
        ELSIF x = 9747 THEN
            sigmoid_f := 2030;
        ELSIF x = 9748 THEN
            sigmoid_f := 2030;
        ELSIF x = 9749 THEN
            sigmoid_f := 2030;
        ELSIF x = 9750 THEN
            sigmoid_f := 2030;
        ELSIF x = 9751 THEN
            sigmoid_f := 2030;
        ELSIF x = 9752 THEN
            sigmoid_f := 2030;
        ELSIF x = 9753 THEN
            sigmoid_f := 2030;
        ELSIF x = 9754 THEN
            sigmoid_f := 2030;
        ELSIF x = 9755 THEN
            sigmoid_f := 2030;
        ELSIF x = 9756 THEN
            sigmoid_f := 2030;
        ELSIF x = 9757 THEN
            sigmoid_f := 2030;
        ELSIF x = 9758 THEN
            sigmoid_f := 2030;
        ELSIF x = 9759 THEN
            sigmoid_f := 2030;
        ELSIF x = 9760 THEN
            sigmoid_f := 2030;
        ELSIF x = 9761 THEN
            sigmoid_f := 2030;
        ELSIF x = 9762 THEN
            sigmoid_f := 2030;
        ELSIF x = 9763 THEN
            sigmoid_f := 2030;
        ELSIF x = 9764 THEN
            sigmoid_f := 2030;
        ELSIF x = 9765 THEN
            sigmoid_f := 2030;
        ELSIF x = 9766 THEN
            sigmoid_f := 2030;
        ELSIF x = 9767 THEN
            sigmoid_f := 2030;
        ELSIF x = 9768 THEN
            sigmoid_f := 2031;
        ELSIF x = 9769 THEN
            sigmoid_f := 2031;
        ELSIF x = 9770 THEN
            sigmoid_f := 2031;
        ELSIF x = 9771 THEN
            sigmoid_f := 2031;
        ELSIF x = 9772 THEN
            sigmoid_f := 2031;
        ELSIF x = 9773 THEN
            sigmoid_f := 2031;
        ELSIF x = 9774 THEN
            sigmoid_f := 2031;
        ELSIF x = 9775 THEN
            sigmoid_f := 2031;
        ELSIF x = 9776 THEN
            sigmoid_f := 2031;
        ELSIF x = 9777 THEN
            sigmoid_f := 2031;
        ELSIF x = 9778 THEN
            sigmoid_f := 2031;
        ELSIF x = 9779 THEN
            sigmoid_f := 2031;
        ELSIF x = 9780 THEN
            sigmoid_f := 2031;
        ELSIF x = 9781 THEN
            sigmoid_f := 2031;
        ELSIF x = 9782 THEN
            sigmoid_f := 2031;
        ELSIF x = 9783 THEN
            sigmoid_f := 2031;
        ELSIF x = 9784 THEN
            sigmoid_f := 2031;
        ELSIF x = 9785 THEN
            sigmoid_f := 2031;
        ELSIF x = 9786 THEN
            sigmoid_f := 2031;
        ELSIF x = 9787 THEN
            sigmoid_f := 2031;
        ELSIF x = 9788 THEN
            sigmoid_f := 2031;
        ELSIF x = 9789 THEN
            sigmoid_f := 2031;
        ELSIF x = 9790 THEN
            sigmoid_f := 2031;
        ELSIF x = 9791 THEN
            sigmoid_f := 2031;
        ELSIF x = 9792 THEN
            sigmoid_f := 2031;
        ELSIF x = 9793 THEN
            sigmoid_f := 2031;
        ELSIF x = 9794 THEN
            sigmoid_f := 2031;
        ELSIF x = 9795 THEN
            sigmoid_f := 2031;
        ELSIF x = 9796 THEN
            sigmoid_f := 2031;
        ELSIF x = 9797 THEN
            sigmoid_f := 2031;
        ELSIF x = 9798 THEN
            sigmoid_f := 2031;
        ELSIF x = 9799 THEN
            sigmoid_f := 2031;
        ELSIF x = 9800 THEN
            sigmoid_f := 2031;
        ELSIF x = 9801 THEN
            sigmoid_f := 2031;
        ELSIF x = 9802 THEN
            sigmoid_f := 2031;
        ELSIF x = 9803 THEN
            sigmoid_f := 2031;
        ELSIF x = 9804 THEN
            sigmoid_f := 2031;
        ELSIF x = 9805 THEN
            sigmoid_f := 2031;
        ELSIF x = 9806 THEN
            sigmoid_f := 2031;
        ELSIF x = 9807 THEN
            sigmoid_f := 2031;
        ELSIF x = 9808 THEN
            sigmoid_f := 2031;
        ELSIF x = 9809 THEN
            sigmoid_f := 2031;
        ELSIF x = 9810 THEN
            sigmoid_f := 2031;
        ELSIF x = 9811 THEN
            sigmoid_f := 2031;
        ELSIF x = 9812 THEN
            sigmoid_f := 2031;
        ELSIF x = 9813 THEN
            sigmoid_f := 2031;
        ELSIF x = 9814 THEN
            sigmoid_f := 2031;
        ELSIF x = 9815 THEN
            sigmoid_f := 2031;
        ELSIF x = 9816 THEN
            sigmoid_f := 2031;
        ELSIF x = 9817 THEN
            sigmoid_f := 2031;
        ELSIF x = 9818 THEN
            sigmoid_f := 2031;
        ELSIF x = 9819 THEN
            sigmoid_f := 2031;
        ELSIF x = 9820 THEN
            sigmoid_f := 2031;
        ELSIF x = 9821 THEN
            sigmoid_f := 2031;
        ELSIF x = 9822 THEN
            sigmoid_f := 2031;
        ELSIF x = 9823 THEN
            sigmoid_f := 2031;
        ELSIF x = 9824 THEN
            sigmoid_f := 2031;
        ELSIF x = 9825 THEN
            sigmoid_f := 2031;
        ELSIF x = 9826 THEN
            sigmoid_f := 2031;
        ELSIF x = 9827 THEN
            sigmoid_f := 2031;
        ELSIF x = 9828 THEN
            sigmoid_f := 2031;
        ELSIF x = 9829 THEN
            sigmoid_f := 2031;
        ELSIF x = 9830 THEN
            sigmoid_f := 2031;
        ELSIF x = 9831 THEN
            sigmoid_f := 2031;
        ELSIF x = 9832 THEN
            sigmoid_f := 2031;
        ELSIF x = 9833 THEN
            sigmoid_f := 2031;
        ELSIF x = 9834 THEN
            sigmoid_f := 2031;
        ELSIF x = 9835 THEN
            sigmoid_f := 2031;
        ELSIF x = 9836 THEN
            sigmoid_f := 2031;
        ELSIF x = 9837 THEN
            sigmoid_f := 2031;
        ELSIF x = 9838 THEN
            sigmoid_f := 2031;
        ELSIF x = 9839 THEN
            sigmoid_f := 2031;
        ELSIF x = 9840 THEN
            sigmoid_f := 2031;
        ELSIF x = 9841 THEN
            sigmoid_f := 2031;
        ELSIF x = 9842 THEN
            sigmoid_f := 2031;
        ELSIF x = 9843 THEN
            sigmoid_f := 2031;
        ELSIF x = 9844 THEN
            sigmoid_f := 2031;
        ELSIF x = 9845 THEN
            sigmoid_f := 2031;
        ELSIF x = 9846 THEN
            sigmoid_f := 2031;
        ELSIF x = 9847 THEN
            sigmoid_f := 2031;
        ELSIF x = 9848 THEN
            sigmoid_f := 2031;
        ELSIF x = 9849 THEN
            sigmoid_f := 2031;
        ELSIF x = 9850 THEN
            sigmoid_f := 2031;
        ELSIF x = 9851 THEN
            sigmoid_f := 2031;
        ELSIF x = 9852 THEN
            sigmoid_f := 2031;
        ELSIF x = 9853 THEN
            sigmoid_f := 2031;
        ELSIF x = 9854 THEN
            sigmoid_f := 2031;
        ELSIF x = 9855 THEN
            sigmoid_f := 2031;
        ELSIF x = 9856 THEN
            sigmoid_f := 2031;
        ELSIF x = 9857 THEN
            sigmoid_f := 2031;
        ELSIF x = 9858 THEN
            sigmoid_f := 2031;
        ELSIF x = 9859 THEN
            sigmoid_f := 2031;
        ELSIF x = 9860 THEN
            sigmoid_f := 2031;
        ELSIF x = 9861 THEN
            sigmoid_f := 2031;
        ELSIF x = 9862 THEN
            sigmoid_f := 2031;
        ELSIF x = 9863 THEN
            sigmoid_f := 2031;
        ELSIF x = 9864 THEN
            sigmoid_f := 2031;
        ELSIF x = 9865 THEN
            sigmoid_f := 2031;
        ELSIF x = 9866 THEN
            sigmoid_f := 2031;
        ELSIF x = 9867 THEN
            sigmoid_f := 2031;
        ELSIF x = 9868 THEN
            sigmoid_f := 2031;
        ELSIF x = 9869 THEN
            sigmoid_f := 2031;
        ELSIF x = 9870 THEN
            sigmoid_f := 2031;
        ELSIF x = 9871 THEN
            sigmoid_f := 2031;
        ELSIF x = 9872 THEN
            sigmoid_f := 2031;
        ELSIF x = 9873 THEN
            sigmoid_f := 2031;
        ELSIF x = 9874 THEN
            sigmoid_f := 2031;
        ELSIF x = 9875 THEN
            sigmoid_f := 2031;
        ELSIF x = 9876 THEN
            sigmoid_f := 2031;
        ELSIF x = 9877 THEN
            sigmoid_f := 2031;
        ELSIF x = 9878 THEN
            sigmoid_f := 2031;
        ELSIF x = 9879 THEN
            sigmoid_f := 2031;
        ELSIF x = 9880 THEN
            sigmoid_f := 2031;
        ELSIF x = 9881 THEN
            sigmoid_f := 2031;
        ELSIF x = 9882 THEN
            sigmoid_f := 2031;
        ELSIF x = 9883 THEN
            sigmoid_f := 2031;
        ELSIF x = 9884 THEN
            sigmoid_f := 2031;
        ELSIF x = 9885 THEN
            sigmoid_f := 2031;
        ELSIF x = 9886 THEN
            sigmoid_f := 2031;
        ELSIF x = 9887 THEN
            sigmoid_f := 2031;
        ELSIF x = 9888 THEN
            sigmoid_f := 2031;
        ELSIF x = 9889 THEN
            sigmoid_f := 2031;
        ELSIF x = 9890 THEN
            sigmoid_f := 2031;
        ELSIF x = 9891 THEN
            sigmoid_f := 2031;
        ELSIF x = 9892 THEN
            sigmoid_f := 2031;
        ELSIF x = 9893 THEN
            sigmoid_f := 2031;
        ELSIF x = 9894 THEN
            sigmoid_f := 2031;
        ELSIF x = 9895 THEN
            sigmoid_f := 2031;
        ELSIF x = 9896 THEN
            sigmoid_f := 2031;
        ELSIF x = 9897 THEN
            sigmoid_f := 2031;
        ELSIF x = 9898 THEN
            sigmoid_f := 2031;
        ELSIF x = 9899 THEN
            sigmoid_f := 2031;
        ELSIF x = 9900 THEN
            sigmoid_f := 2031;
        ELSIF x = 9901 THEN
            sigmoid_f := 2031;
        ELSIF x = 9902 THEN
            sigmoid_f := 2031;
        ELSIF x = 9903 THEN
            sigmoid_f := 2031;
        ELSIF x = 9904 THEN
            sigmoid_f := 2031;
        ELSIF x = 9905 THEN
            sigmoid_f := 2031;
        ELSIF x = 9906 THEN
            sigmoid_f := 2031;
        ELSIF x = 9907 THEN
            sigmoid_f := 2031;
        ELSIF x = 9908 THEN
            sigmoid_f := 2031;
        ELSIF x = 9909 THEN
            sigmoid_f := 2031;
        ELSIF x = 9910 THEN
            sigmoid_f := 2031;
        ELSIF x = 9911 THEN
            sigmoid_f := 2031;
        ELSIF x = 9912 THEN
            sigmoid_f := 2031;
        ELSIF x = 9913 THEN
            sigmoid_f := 2031;
        ELSIF x = 9914 THEN
            sigmoid_f := 2031;
        ELSIF x = 9915 THEN
            sigmoid_f := 2031;
        ELSIF x = 9916 THEN
            sigmoid_f := 2031;
        ELSIF x = 9917 THEN
            sigmoid_f := 2031;
        ELSIF x = 9918 THEN
            sigmoid_f := 2031;
        ELSIF x = 9919 THEN
            sigmoid_f := 2031;
        ELSIF x = 9920 THEN
            sigmoid_f := 2031;
        ELSIF x = 9921 THEN
            sigmoid_f := 2031;
        ELSIF x = 9922 THEN
            sigmoid_f := 2031;
        ELSIF x = 9923 THEN
            sigmoid_f := 2031;
        ELSIF x = 9924 THEN
            sigmoid_f := 2031;
        ELSIF x = 9925 THEN
            sigmoid_f := 2032;
        ELSIF x = 9926 THEN
            sigmoid_f := 2032;
        ELSIF x = 9927 THEN
            sigmoid_f := 2032;
        ELSIF x = 9928 THEN
            sigmoid_f := 2032;
        ELSIF x = 9929 THEN
            sigmoid_f := 2032;
        ELSIF x = 9930 THEN
            sigmoid_f := 2032;
        ELSIF x = 9931 THEN
            sigmoid_f := 2032;
        ELSIF x = 9932 THEN
            sigmoid_f := 2032;
        ELSIF x = 9933 THEN
            sigmoid_f := 2032;
        ELSIF x = 9934 THEN
            sigmoid_f := 2032;
        ELSIF x = 9935 THEN
            sigmoid_f := 2032;
        ELSIF x = 9936 THEN
            sigmoid_f := 2032;
        ELSIF x = 9937 THEN
            sigmoid_f := 2032;
        ELSIF x = 9938 THEN
            sigmoid_f := 2032;
        ELSIF x = 9939 THEN
            sigmoid_f := 2032;
        ELSIF x = 9940 THEN
            sigmoid_f := 2032;
        ELSIF x = 9941 THEN
            sigmoid_f := 2032;
        ELSIF x = 9942 THEN
            sigmoid_f := 2032;
        ELSIF x = 9943 THEN
            sigmoid_f := 2032;
        ELSIF x = 9944 THEN
            sigmoid_f := 2032;
        ELSIF x = 9945 THEN
            sigmoid_f := 2032;
        ELSIF x = 9946 THEN
            sigmoid_f := 2032;
        ELSIF x = 9947 THEN
            sigmoid_f := 2032;
        ELSIF x = 9948 THEN
            sigmoid_f := 2032;
        ELSIF x = 9949 THEN
            sigmoid_f := 2032;
        ELSIF x = 9950 THEN
            sigmoid_f := 2032;
        ELSIF x = 9951 THEN
            sigmoid_f := 2032;
        ELSIF x = 9952 THEN
            sigmoid_f := 2032;
        ELSIF x = 9953 THEN
            sigmoid_f := 2032;
        ELSIF x = 9954 THEN
            sigmoid_f := 2032;
        ELSIF x = 9955 THEN
            sigmoid_f := 2032;
        ELSIF x = 9956 THEN
            sigmoid_f := 2032;
        ELSIF x = 9957 THEN
            sigmoid_f := 2032;
        ELSIF x = 9958 THEN
            sigmoid_f := 2032;
        ELSIF x = 9959 THEN
            sigmoid_f := 2032;
        ELSIF x = 9960 THEN
            sigmoid_f := 2032;
        ELSIF x = 9961 THEN
            sigmoid_f := 2032;
        ELSIF x = 9962 THEN
            sigmoid_f := 2032;
        ELSIF x = 9963 THEN
            sigmoid_f := 2032;
        ELSIF x = 9964 THEN
            sigmoid_f := 2032;
        ELSIF x = 9965 THEN
            sigmoid_f := 2032;
        ELSIF x = 9966 THEN
            sigmoid_f := 2032;
        ELSIF x = 9967 THEN
            sigmoid_f := 2032;
        ELSIF x = 9968 THEN
            sigmoid_f := 2032;
        ELSIF x = 9969 THEN
            sigmoid_f := 2032;
        ELSIF x = 9970 THEN
            sigmoid_f := 2032;
        ELSIF x = 9971 THEN
            sigmoid_f := 2032;
        ELSIF x = 9972 THEN
            sigmoid_f := 2032;
        ELSIF x = 9973 THEN
            sigmoid_f := 2032;
        ELSIF x = 9974 THEN
            sigmoid_f := 2032;
        ELSIF x = 9975 THEN
            sigmoid_f := 2032;
        ELSIF x = 9976 THEN
            sigmoid_f := 2032;
        ELSIF x = 9977 THEN
            sigmoid_f := 2032;
        ELSIF x = 9978 THEN
            sigmoid_f := 2032;
        ELSIF x = 9979 THEN
            sigmoid_f := 2032;
        ELSIF x = 9980 THEN
            sigmoid_f := 2032;
        ELSIF x = 9981 THEN
            sigmoid_f := 2032;
        ELSIF x = 9982 THEN
            sigmoid_f := 2032;
        ELSIF x = 9983 THEN
            sigmoid_f := 2032;
        ELSIF x = 9984 THEN
            sigmoid_f := 2032;
        ELSIF x = 9985 THEN
            sigmoid_f := 2032;
        ELSIF x = 9986 THEN
            sigmoid_f := 2032;
        ELSIF x = 9987 THEN
            sigmoid_f := 2032;
        ELSIF x = 9988 THEN
            sigmoid_f := 2032;
        ELSIF x = 9989 THEN
            sigmoid_f := 2032;
        ELSIF x = 9990 THEN
            sigmoid_f := 2032;
        ELSIF x = 9991 THEN
            sigmoid_f := 2032;
        ELSIF x = 9992 THEN
            sigmoid_f := 2032;
        ELSIF x = 9993 THEN
            sigmoid_f := 2032;
        ELSIF x = 9994 THEN
            sigmoid_f := 2032;
        ELSIF x = 9995 THEN
            sigmoid_f := 2032;
        ELSIF x = 9996 THEN
            sigmoid_f := 2032;
        ELSIF x = 9997 THEN
            sigmoid_f := 2032;
        ELSIF x = 9998 THEN
            sigmoid_f := 2032;
        ELSIF x = 9999 THEN
            sigmoid_f := 2032;
        ELSIF x = 10000 THEN
            sigmoid_f := 2032;
        ELSIF x = 10001 THEN
            sigmoid_f := 2032;
        ELSIF x = 10002 THEN
            sigmoid_f := 2032;
        ELSIF x = 10003 THEN
            sigmoid_f := 2032;
        ELSIF x = 10004 THEN
            sigmoid_f := 2032;
        ELSIF x = 10005 THEN
            sigmoid_f := 2032;
        ELSIF x = 10006 THEN
            sigmoid_f := 2032;
        ELSIF x = 10007 THEN
            sigmoid_f := 2032;
        ELSIF x = 10008 THEN
            sigmoid_f := 2032;
        ELSIF x = 10009 THEN
            sigmoid_f := 2032;
        ELSIF x = 10010 THEN
            sigmoid_f := 2032;
        ELSIF x = 10011 THEN
            sigmoid_f := 2032;
        ELSIF x = 10012 THEN
            sigmoid_f := 2032;
        ELSIF x = 10013 THEN
            sigmoid_f := 2032;
        ELSIF x = 10014 THEN
            sigmoid_f := 2032;
        ELSIF x = 10015 THEN
            sigmoid_f := 2032;
        ELSIF x = 10016 THEN
            sigmoid_f := 2032;
        ELSIF x = 10017 THEN
            sigmoid_f := 2032;
        ELSIF x = 10018 THEN
            sigmoid_f := 2032;
        ELSIF x = 10019 THEN
            sigmoid_f := 2032;
        ELSIF x = 10020 THEN
            sigmoid_f := 2032;
        ELSIF x = 10021 THEN
            sigmoid_f := 2032;
        ELSIF x = 10022 THEN
            sigmoid_f := 2032;
        ELSIF x = 10023 THEN
            sigmoid_f := 2032;
        ELSIF x = 10024 THEN
            sigmoid_f := 2032;
        ELSIF x = 10025 THEN
            sigmoid_f := 2032;
        ELSIF x = 10026 THEN
            sigmoid_f := 2032;
        ELSIF x = 10027 THEN
            sigmoid_f := 2032;
        ELSIF x = 10028 THEN
            sigmoid_f := 2032;
        ELSIF x = 10029 THEN
            sigmoid_f := 2032;
        ELSIF x = 10030 THEN
            sigmoid_f := 2032;
        ELSIF x = 10031 THEN
            sigmoid_f := 2032;
        ELSIF x = 10032 THEN
            sigmoid_f := 2032;
        ELSIF x = 10033 THEN
            sigmoid_f := 2032;
        ELSIF x = 10034 THEN
            sigmoid_f := 2032;
        ELSIF x = 10035 THEN
            sigmoid_f := 2032;
        ELSIF x = 10036 THEN
            sigmoid_f := 2032;
        ELSIF x = 10037 THEN
            sigmoid_f := 2032;
        ELSIF x = 10038 THEN
            sigmoid_f := 2032;
        ELSIF x = 10039 THEN
            sigmoid_f := 2032;
        ELSIF x = 10040 THEN
            sigmoid_f := 2032;
        ELSIF x = 10041 THEN
            sigmoid_f := 2032;
        ELSIF x = 10042 THEN
            sigmoid_f := 2032;
        ELSIF x = 10043 THEN
            sigmoid_f := 2032;
        ELSIF x = 10044 THEN
            sigmoid_f := 2032;
        ELSIF x = 10045 THEN
            sigmoid_f := 2032;
        ELSIF x = 10046 THEN
            sigmoid_f := 2032;
        ELSIF x = 10047 THEN
            sigmoid_f := 2032;
        ELSIF x = 10048 THEN
            sigmoid_f := 2032;
        ELSIF x = 10049 THEN
            sigmoid_f := 2032;
        ELSIF x = 10050 THEN
            sigmoid_f := 2032;
        ELSIF x = 10051 THEN
            sigmoid_f := 2032;
        ELSIF x = 10052 THEN
            sigmoid_f := 2032;
        ELSIF x = 10053 THEN
            sigmoid_f := 2032;
        ELSIF x = 10054 THEN
            sigmoid_f := 2032;
        ELSIF x = 10055 THEN
            sigmoid_f := 2032;
        ELSIF x = 10056 THEN
            sigmoid_f := 2032;
        ELSIF x = 10057 THEN
            sigmoid_f := 2032;
        ELSIF x = 10058 THEN
            sigmoid_f := 2032;
        ELSIF x = 10059 THEN
            sigmoid_f := 2032;
        ELSIF x = 10060 THEN
            sigmoid_f := 2032;
        ELSIF x = 10061 THEN
            sigmoid_f := 2032;
        ELSIF x = 10062 THEN
            sigmoid_f := 2032;
        ELSIF x = 10063 THEN
            sigmoid_f := 2032;
        ELSIF x = 10064 THEN
            sigmoid_f := 2032;
        ELSIF x = 10065 THEN
            sigmoid_f := 2032;
        ELSIF x = 10066 THEN
            sigmoid_f := 2032;
        ELSIF x = 10067 THEN
            sigmoid_f := 2032;
        ELSIF x = 10068 THEN
            sigmoid_f := 2032;
        ELSIF x = 10069 THEN
            sigmoid_f := 2032;
        ELSIF x = 10070 THEN
            sigmoid_f := 2032;
        ELSIF x = 10071 THEN
            sigmoid_f := 2032;
        ELSIF x = 10072 THEN
            sigmoid_f := 2032;
        ELSIF x = 10073 THEN
            sigmoid_f := 2032;
        ELSIF x = 10074 THEN
            sigmoid_f := 2032;
        ELSIF x = 10075 THEN
            sigmoid_f := 2032;
        ELSIF x = 10076 THEN
            sigmoid_f := 2032;
        ELSIF x = 10077 THEN
            sigmoid_f := 2032;
        ELSIF x = 10078 THEN
            sigmoid_f := 2032;
        ELSIF x = 10079 THEN
            sigmoid_f := 2032;
        ELSIF x = 10080 THEN
            sigmoid_f := 2032;
        ELSIF x = 10081 THEN
            sigmoid_f := 2032;
        ELSIF x = 10082 THEN
            sigmoid_f := 2032;
        ELSIF x = 10083 THEN
            sigmoid_f := 2033;
        ELSIF x = 10084 THEN
            sigmoid_f := 2033;
        ELSIF x = 10085 THEN
            sigmoid_f := 2033;
        ELSIF x = 10086 THEN
            sigmoid_f := 2033;
        ELSIF x = 10087 THEN
            sigmoid_f := 2033;
        ELSIF x = 10088 THEN
            sigmoid_f := 2033;
        ELSIF x = 10089 THEN
            sigmoid_f := 2033;
        ELSIF x = 10090 THEN
            sigmoid_f := 2033;
        ELSIF x = 10091 THEN
            sigmoid_f := 2033;
        ELSIF x = 10092 THEN
            sigmoid_f := 2033;
        ELSIF x = 10093 THEN
            sigmoid_f := 2033;
        ELSIF x = 10094 THEN
            sigmoid_f := 2033;
        ELSIF x = 10095 THEN
            sigmoid_f := 2033;
        ELSIF x = 10096 THEN
            sigmoid_f := 2033;
        ELSIF x = 10097 THEN
            sigmoid_f := 2033;
        ELSIF x = 10098 THEN
            sigmoid_f := 2033;
        ELSIF x = 10099 THEN
            sigmoid_f := 2033;
        ELSIF x = 10100 THEN
            sigmoid_f := 2033;
        ELSIF x = 10101 THEN
            sigmoid_f := 2033;
        ELSIF x = 10102 THEN
            sigmoid_f := 2033;
        ELSIF x = 10103 THEN
            sigmoid_f := 2033;
        ELSIF x = 10104 THEN
            sigmoid_f := 2033;
        ELSIF x = 10105 THEN
            sigmoid_f := 2033;
        ELSIF x = 10106 THEN
            sigmoid_f := 2033;
        ELSIF x = 10107 THEN
            sigmoid_f := 2033;
        ELSIF x = 10108 THEN
            sigmoid_f := 2033;
        ELSIF x = 10109 THEN
            sigmoid_f := 2033;
        ELSIF x = 10110 THEN
            sigmoid_f := 2033;
        ELSIF x = 10111 THEN
            sigmoid_f := 2033;
        ELSIF x = 10112 THEN
            sigmoid_f := 2033;
        ELSIF x = 10113 THEN
            sigmoid_f := 2033;
        ELSIF x = 10114 THEN
            sigmoid_f := 2033;
        ELSIF x = 10115 THEN
            sigmoid_f := 2033;
        ELSIF x = 10116 THEN
            sigmoid_f := 2033;
        ELSIF x = 10117 THEN
            sigmoid_f := 2033;
        ELSIF x = 10118 THEN
            sigmoid_f := 2033;
        ELSIF x = 10119 THEN
            sigmoid_f := 2033;
        ELSIF x = 10120 THEN
            sigmoid_f := 2033;
        ELSIF x = 10121 THEN
            sigmoid_f := 2033;
        ELSIF x = 10122 THEN
            sigmoid_f := 2033;
        ELSIF x = 10123 THEN
            sigmoid_f := 2033;
        ELSIF x = 10124 THEN
            sigmoid_f := 2033;
        ELSIF x = 10125 THEN
            sigmoid_f := 2033;
        ELSIF x = 10126 THEN
            sigmoid_f := 2033;
        ELSIF x = 10127 THEN
            sigmoid_f := 2033;
        ELSIF x = 10128 THEN
            sigmoid_f := 2033;
        ELSIF x = 10129 THEN
            sigmoid_f := 2033;
        ELSIF x = 10130 THEN
            sigmoid_f := 2033;
        ELSIF x = 10131 THEN
            sigmoid_f := 2033;
        ELSIF x = 10132 THEN
            sigmoid_f := 2033;
        ELSIF x = 10133 THEN
            sigmoid_f := 2033;
        ELSIF x = 10134 THEN
            sigmoid_f := 2033;
        ELSIF x = 10135 THEN
            sigmoid_f := 2033;
        ELSIF x = 10136 THEN
            sigmoid_f := 2033;
        ELSIF x = 10137 THEN
            sigmoid_f := 2033;
        ELSIF x = 10138 THEN
            sigmoid_f := 2033;
        ELSIF x = 10139 THEN
            sigmoid_f := 2033;
        ELSIF x = 10140 THEN
            sigmoid_f := 2033;
        ELSIF x = 10141 THEN
            sigmoid_f := 2033;
        ELSIF x = 10142 THEN
            sigmoid_f := 2033;
        ELSIF x = 10143 THEN
            sigmoid_f := 2033;
        ELSIF x = 10144 THEN
            sigmoid_f := 2033;
        ELSIF x = 10145 THEN
            sigmoid_f := 2033;
        ELSIF x = 10146 THEN
            sigmoid_f := 2033;
        ELSIF x = 10147 THEN
            sigmoid_f := 2033;
        ELSIF x = 10148 THEN
            sigmoid_f := 2033;
        ELSIF x = 10149 THEN
            sigmoid_f := 2033;
        ELSIF x = 10150 THEN
            sigmoid_f := 2033;
        ELSIF x = 10151 THEN
            sigmoid_f := 2033;
        ELSIF x = 10152 THEN
            sigmoid_f := 2033;
        ELSIF x = 10153 THEN
            sigmoid_f := 2033;
        ELSIF x = 10154 THEN
            sigmoid_f := 2033;
        ELSIF x = 10155 THEN
            sigmoid_f := 2033;
        ELSIF x = 10156 THEN
            sigmoid_f := 2033;
        ELSIF x = 10157 THEN
            sigmoid_f := 2033;
        ELSIF x = 10158 THEN
            sigmoid_f := 2033;
        ELSIF x = 10159 THEN
            sigmoid_f := 2033;
        ELSIF x = 10160 THEN
            sigmoid_f := 2033;
        ELSIF x = 10161 THEN
            sigmoid_f := 2033;
        ELSIF x = 10162 THEN
            sigmoid_f := 2033;
        ELSIF x = 10163 THEN
            sigmoid_f := 2033;
        ELSIF x = 10164 THEN
            sigmoid_f := 2033;
        ELSIF x = 10165 THEN
            sigmoid_f := 2033;
        ELSIF x = 10166 THEN
            sigmoid_f := 2033;
        ELSIF x = 10167 THEN
            sigmoid_f := 2033;
        ELSIF x = 10168 THEN
            sigmoid_f := 2033;
        ELSIF x = 10169 THEN
            sigmoid_f := 2033;
        ELSIF x = 10170 THEN
            sigmoid_f := 2033;
        ELSIF x = 10171 THEN
            sigmoid_f := 2033;
        ELSIF x = 10172 THEN
            sigmoid_f := 2033;
        ELSIF x = 10173 THEN
            sigmoid_f := 2033;
        ELSIF x = 10174 THEN
            sigmoid_f := 2033;
        ELSIF x = 10175 THEN
            sigmoid_f := 2033;
        ELSIF x = 10176 THEN
            sigmoid_f := 2033;
        ELSIF x = 10177 THEN
            sigmoid_f := 2033;
        ELSIF x = 10178 THEN
            sigmoid_f := 2033;
        ELSIF x = 10179 THEN
            sigmoid_f := 2033;
        ELSIF x = 10180 THEN
            sigmoid_f := 2033;
        ELSIF x = 10181 THEN
            sigmoid_f := 2033;
        ELSIF x = 10182 THEN
            sigmoid_f := 2033;
        ELSIF x = 10183 THEN
            sigmoid_f := 2033;
        ELSIF x = 10184 THEN
            sigmoid_f := 2033;
        ELSIF x = 10185 THEN
            sigmoid_f := 2033;
        ELSIF x = 10186 THEN
            sigmoid_f := 2033;
        ELSIF x = 10187 THEN
            sigmoid_f := 2033;
        ELSIF x = 10188 THEN
            sigmoid_f := 2033;
        ELSIF x = 10189 THEN
            sigmoid_f := 2033;
        ELSIF x = 10190 THEN
            sigmoid_f := 2033;
        ELSIF x = 10191 THEN
            sigmoid_f := 2033;
        ELSIF x = 10192 THEN
            sigmoid_f := 2033;
        ELSIF x = 10193 THEN
            sigmoid_f := 2033;
        ELSIF x = 10194 THEN
            sigmoid_f := 2033;
        ELSIF x = 10195 THEN
            sigmoid_f := 2033;
        ELSIF x = 10196 THEN
            sigmoid_f := 2033;
        ELSIF x = 10197 THEN
            sigmoid_f := 2033;
        ELSIF x = 10198 THEN
            sigmoid_f := 2033;
        ELSIF x = 10199 THEN
            sigmoid_f := 2033;
        ELSIF x = 10200 THEN
            sigmoid_f := 2033;
        ELSIF x = 10201 THEN
            sigmoid_f := 2033;
        ELSIF x = 10202 THEN
            sigmoid_f := 2033;
        ELSIF x = 10203 THEN
            sigmoid_f := 2033;
        ELSIF x = 10204 THEN
            sigmoid_f := 2033;
        ELSIF x = 10205 THEN
            sigmoid_f := 2033;
        ELSIF x = 10206 THEN
            sigmoid_f := 2033;
        ELSIF x = 10207 THEN
            sigmoid_f := 2033;
        ELSIF x = 10208 THEN
            sigmoid_f := 2033;
        ELSIF x = 10209 THEN
            sigmoid_f := 2033;
        ELSIF x = 10210 THEN
            sigmoid_f := 2033;
        ELSIF x = 10211 THEN
            sigmoid_f := 2033;
        ELSIF x = 10212 THEN
            sigmoid_f := 2033;
        ELSIF x = 10213 THEN
            sigmoid_f := 2033;
        ELSIF x = 10214 THEN
            sigmoid_f := 2033;
        ELSIF x = 10215 THEN
            sigmoid_f := 2033;
        ELSIF x = 10216 THEN
            sigmoid_f := 2033;
        ELSIF x = 10217 THEN
            sigmoid_f := 2033;
        ELSIF x = 10218 THEN
            sigmoid_f := 2033;
        ELSIF x = 10219 THEN
            sigmoid_f := 2033;
        ELSIF x = 10220 THEN
            sigmoid_f := 2033;
        ELSIF x = 10221 THEN
            sigmoid_f := 2033;
        ELSIF x = 10222 THEN
            sigmoid_f := 2033;
        ELSIF x = 10223 THEN
            sigmoid_f := 2033;
        ELSIF x = 10224 THEN
            sigmoid_f := 2033;
        ELSIF x = 10225 THEN
            sigmoid_f := 2033;
        ELSIF x = 10226 THEN
            sigmoid_f := 2033;
        ELSIF x = 10227 THEN
            sigmoid_f := 2033;
        ELSIF x = 10228 THEN
            sigmoid_f := 2033;
        ELSIF x = 10229 THEN
            sigmoid_f := 2033;
        ELSIF x = 10230 THEN
            sigmoid_f := 2033;
        ELSIF x = 10231 THEN
            sigmoid_f := 2033;
        ELSIF x = 10232 THEN
            sigmoid_f := 2033;
        ELSIF x = 10233 THEN
            sigmoid_f := 2033;
        ELSIF x = 10234 THEN
            sigmoid_f := 2033;
        ELSIF x = 10235 THEN
            sigmoid_f := 2033;
        ELSIF x = 10236 THEN
            sigmoid_f := 2033;
        ELSIF x = 10237 THEN
            sigmoid_f := 2033;
        ELSIF x = 10238 THEN
            sigmoid_f := 2033;
        ELSIF x = 10239 THEN
            sigmoid_f := 2033;
        ELSIF x = 10240 THEN
            sigmoid_f := 2034;
        ELSIF x = 10241 THEN
            sigmoid_f := 2034;
        ELSIF x = 10242 THEN
            sigmoid_f := 2034;
        ELSIF x = 10243 THEN
            sigmoid_f := 2034;
        ELSIF x = 10244 THEN
            sigmoid_f := 2034;
        ELSIF x = 10245 THEN
            sigmoid_f := 2034;
        ELSIF x = 10246 THEN
            sigmoid_f := 2034;
        ELSIF x = 10247 THEN
            sigmoid_f := 2034;
        ELSIF x = 10248 THEN
            sigmoid_f := 2034;
        ELSIF x = 10249 THEN
            sigmoid_f := 2034;
        ELSIF x = 10250 THEN
            sigmoid_f := 2034;
        ELSIF x = 10251 THEN
            sigmoid_f := 2034;
        ELSIF x = 10252 THEN
            sigmoid_f := 2034;
        ELSIF x = 10253 THEN
            sigmoid_f := 2034;
        ELSIF x = 10254 THEN
            sigmoid_f := 2034;
        ELSIF x = 10255 THEN
            sigmoid_f := 2034;
        ELSIF x = 10256 THEN
            sigmoid_f := 2034;
        ELSIF x = 10257 THEN
            sigmoid_f := 2034;
        ELSIF x = 10258 THEN
            sigmoid_f := 2034;
        ELSIF x = 10259 THEN
            sigmoid_f := 2034;
        ELSIF x = 10260 THEN
            sigmoid_f := 2034;
        ELSIF x = 10261 THEN
            sigmoid_f := 2034;
        ELSIF x = 10262 THEN
            sigmoid_f := 2034;
        ELSIF x = 10263 THEN
            sigmoid_f := 2034;
        ELSIF x = 10264 THEN
            sigmoid_f := 2034;
        ELSIF x = 10265 THEN
            sigmoid_f := 2034;
        ELSIF x = 10266 THEN
            sigmoid_f := 2034;
        ELSIF x = 10267 THEN
            sigmoid_f := 2034;
        ELSIF x = 10268 THEN
            sigmoid_f := 2034;
        ELSIF x = 10269 THEN
            sigmoid_f := 2034;
        ELSIF x = 10270 THEN
            sigmoid_f := 2034;
        ELSIF x = 10271 THEN
            sigmoid_f := 2034;
        ELSIF x = 10272 THEN
            sigmoid_f := 2034;
        ELSIF x = 10273 THEN
            sigmoid_f := 2034;
        ELSIF x = 10274 THEN
            sigmoid_f := 2034;
        ELSIF x = 10275 THEN
            sigmoid_f := 2034;
        ELSIF x = 10276 THEN
            sigmoid_f := 2034;
        ELSIF x = 10277 THEN
            sigmoid_f := 2034;
        ELSIF x = 10278 THEN
            sigmoid_f := 2034;
        ELSIF x = 10279 THEN
            sigmoid_f := 2034;
        ELSIF x = 10280 THEN
            sigmoid_f := 2034;
        ELSIF x = 10281 THEN
            sigmoid_f := 2034;
        ELSIF x = 10282 THEN
            sigmoid_f := 2034;
        ELSIF x = 10283 THEN
            sigmoid_f := 2034;
        ELSIF x = 10284 THEN
            sigmoid_f := 2034;
        ELSIF x = 10285 THEN
            sigmoid_f := 2034;
        ELSIF x = 10286 THEN
            sigmoid_f := 2034;
        ELSIF x = 10287 THEN
            sigmoid_f := 2034;
        ELSIF x = 10288 THEN
            sigmoid_f := 2034;
        ELSIF x = 10289 THEN
            sigmoid_f := 2034;
        ELSIF x = 10290 THEN
            sigmoid_f := 2034;
        ELSIF x = 10291 THEN
            sigmoid_f := 2034;
        ELSIF x = 10292 THEN
            sigmoid_f := 2034;
        ELSIF x = 10293 THEN
            sigmoid_f := 2034;
        ELSIF x = 10294 THEN
            sigmoid_f := 2034;
        ELSIF x = 10295 THEN
            sigmoid_f := 2034;
        ELSIF x = 10296 THEN
            sigmoid_f := 2034;
        ELSIF x = 10297 THEN
            sigmoid_f := 2034;
        ELSIF x = 10298 THEN
            sigmoid_f := 2034;
        ELSIF x = 10299 THEN
            sigmoid_f := 2034;
        ELSIF x = 10300 THEN
            sigmoid_f := 2034;
        ELSIF x = 10301 THEN
            sigmoid_f := 2034;
        ELSIF x = 10302 THEN
            sigmoid_f := 2034;
        ELSIF x = 10303 THEN
            sigmoid_f := 2034;
        ELSIF x = 10304 THEN
            sigmoid_f := 2034;
        ELSIF x = 10305 THEN
            sigmoid_f := 2034;
        ELSIF x = 10306 THEN
            sigmoid_f := 2034;
        ELSIF x = 10307 THEN
            sigmoid_f := 2034;
        ELSIF x = 10308 THEN
            sigmoid_f := 2034;
        ELSIF x = 10309 THEN
            sigmoid_f := 2034;
        ELSIF x = 10310 THEN
            sigmoid_f := 2034;
        ELSIF x = 10311 THEN
            sigmoid_f := 2034;
        ELSIF x = 10312 THEN
            sigmoid_f := 2034;
        ELSIF x = 10313 THEN
            sigmoid_f := 2034;
        ELSIF x = 10314 THEN
            sigmoid_f := 2034;
        ELSIF x = 10315 THEN
            sigmoid_f := 2034;
        ELSIF x = 10316 THEN
            sigmoid_f := 2034;
        ELSIF x = 10317 THEN
            sigmoid_f := 2034;
        ELSIF x = 10318 THEN
            sigmoid_f := 2034;
        ELSIF x = 10319 THEN
            sigmoid_f := 2034;
        ELSIF x = 10320 THEN
            sigmoid_f := 2034;
        ELSIF x = 10321 THEN
            sigmoid_f := 2034;
        ELSIF x = 10322 THEN
            sigmoid_f := 2034;
        ELSIF x = 10323 THEN
            sigmoid_f := 2034;
        ELSIF x = 10324 THEN
            sigmoid_f := 2034;
        ELSIF x = 10325 THEN
            sigmoid_f := 2034;
        ELSIF x = 10326 THEN
            sigmoid_f := 2034;
        ELSIF x = 10327 THEN
            sigmoid_f := 2034;
        ELSIF x = 10328 THEN
            sigmoid_f := 2034;
        ELSIF x = 10329 THEN
            sigmoid_f := 2034;
        ELSIF x = 10330 THEN
            sigmoid_f := 2034;
        ELSIF x = 10331 THEN
            sigmoid_f := 2034;
        ELSIF x = 10332 THEN
            sigmoid_f := 2034;
        ELSIF x = 10333 THEN
            sigmoid_f := 2034;
        ELSIF x = 10334 THEN
            sigmoid_f := 2034;
        ELSIF x = 10335 THEN
            sigmoid_f := 2034;
        ELSIF x = 10336 THEN
            sigmoid_f := 2034;
        ELSIF x = 10337 THEN
            sigmoid_f := 2034;
        ELSIF x = 10338 THEN
            sigmoid_f := 2034;
        ELSIF x = 10339 THEN
            sigmoid_f := 2034;
        ELSIF x = 10340 THEN
            sigmoid_f := 2034;
        ELSIF x = 10341 THEN
            sigmoid_f := 2034;
        ELSIF x = 10342 THEN
            sigmoid_f := 2034;
        ELSIF x = 10343 THEN
            sigmoid_f := 2034;
        ELSIF x = 10344 THEN
            sigmoid_f := 2034;
        ELSIF x = 10345 THEN
            sigmoid_f := 2034;
        ELSIF x = 10346 THEN
            sigmoid_f := 2034;
        ELSIF x = 10347 THEN
            sigmoid_f := 2034;
        ELSIF x = 10348 THEN
            sigmoid_f := 2034;
        ELSIF x = 10349 THEN
            sigmoid_f := 2034;
        ELSIF x = 10350 THEN
            sigmoid_f := 2034;
        ELSIF x = 10351 THEN
            sigmoid_f := 2034;
        ELSIF x = 10352 THEN
            sigmoid_f := 2034;
        ELSIF x = 10353 THEN
            sigmoid_f := 2034;
        ELSIF x = 10354 THEN
            sigmoid_f := 2034;
        ELSIF x = 10355 THEN
            sigmoid_f := 2034;
        ELSIF x = 10356 THEN
            sigmoid_f := 2034;
        ELSIF x = 10357 THEN
            sigmoid_f := 2034;
        ELSIF x = 10358 THEN
            sigmoid_f := 2034;
        ELSIF x = 10359 THEN
            sigmoid_f := 2034;
        ELSIF x = 10360 THEN
            sigmoid_f := 2034;
        ELSIF x = 10361 THEN
            sigmoid_f := 2034;
        ELSIF x = 10362 THEN
            sigmoid_f := 2034;
        ELSIF x = 10363 THEN
            sigmoid_f := 2034;
        ELSIF x = 10364 THEN
            sigmoid_f := 2034;
        ELSIF x = 10365 THEN
            sigmoid_f := 2034;
        ELSIF x = 10366 THEN
            sigmoid_f := 2034;
        ELSIF x = 10367 THEN
            sigmoid_f := 2034;
        ELSIF x = 10368 THEN
            sigmoid_f := 2034;
        ELSIF x = 10369 THEN
            sigmoid_f := 2034;
        ELSIF x = 10370 THEN
            sigmoid_f := 2034;
        ELSIF x = 10371 THEN
            sigmoid_f := 2034;
        ELSIF x = 10372 THEN
            sigmoid_f := 2034;
        ELSIF x = 10373 THEN
            sigmoid_f := 2034;
        ELSIF x = 10374 THEN
            sigmoid_f := 2034;
        ELSIF x = 10375 THEN
            sigmoid_f := 2034;
        ELSIF x = 10376 THEN
            sigmoid_f := 2034;
        ELSIF x = 10377 THEN
            sigmoid_f := 2034;
        ELSIF x = 10378 THEN
            sigmoid_f := 2034;
        ELSIF x = 10379 THEN
            sigmoid_f := 2034;
        ELSIF x = 10380 THEN
            sigmoid_f := 2034;
        ELSIF x = 10381 THEN
            sigmoid_f := 2034;
        ELSIF x = 10382 THEN
            sigmoid_f := 2034;
        ELSIF x = 10383 THEN
            sigmoid_f := 2034;
        ELSIF x = 10384 THEN
            sigmoid_f := 2034;
        ELSIF x = 10385 THEN
            sigmoid_f := 2034;
        ELSIF x = 10386 THEN
            sigmoid_f := 2034;
        ELSIF x = 10387 THEN
            sigmoid_f := 2035;
        ELSIF x = 10388 THEN
            sigmoid_f := 2035;
        ELSIF x = 10389 THEN
            sigmoid_f := 2035;
        ELSIF x = 10390 THEN
            sigmoid_f := 2035;
        ELSIF x = 10391 THEN
            sigmoid_f := 2035;
        ELSIF x = 10392 THEN
            sigmoid_f := 2035;
        ELSIF x = 10393 THEN
            sigmoid_f := 2035;
        ELSIF x = 10394 THEN
            sigmoid_f := 2035;
        ELSIF x = 10395 THEN
            sigmoid_f := 2035;
        ELSIF x = 10396 THEN
            sigmoid_f := 2035;
        ELSIF x = 10397 THEN
            sigmoid_f := 2035;
        ELSIF x = 10398 THEN
            sigmoid_f := 2035;
        ELSIF x = 10399 THEN
            sigmoid_f := 2035;
        ELSIF x = 10400 THEN
            sigmoid_f := 2035;
        ELSIF x = 10401 THEN
            sigmoid_f := 2035;
        ELSIF x = 10402 THEN
            sigmoid_f := 2035;
        ELSIF x = 10403 THEN
            sigmoid_f := 2035;
        ELSIF x = 10404 THEN
            sigmoid_f := 2035;
        ELSIF x = 10405 THEN
            sigmoid_f := 2035;
        ELSIF x = 10406 THEN
            sigmoid_f := 2035;
        ELSIF x = 10407 THEN
            sigmoid_f := 2035;
        ELSIF x = 10408 THEN
            sigmoid_f := 2035;
        ELSIF x = 10409 THEN
            sigmoid_f := 2035;
        ELSIF x = 10410 THEN
            sigmoid_f := 2035;
        ELSIF x = 10411 THEN
            sigmoid_f := 2035;
        ELSIF x = 10412 THEN
            sigmoid_f := 2035;
        ELSIF x = 10413 THEN
            sigmoid_f := 2035;
        ELSIF x = 10414 THEN
            sigmoid_f := 2035;
        ELSIF x = 10415 THEN
            sigmoid_f := 2035;
        ELSIF x = 10416 THEN
            sigmoid_f := 2035;
        ELSIF x = 10417 THEN
            sigmoid_f := 2035;
        ELSIF x = 10418 THEN
            sigmoid_f := 2035;
        ELSIF x = 10419 THEN
            sigmoid_f := 2035;
        ELSIF x = 10420 THEN
            sigmoid_f := 2035;
        ELSIF x = 10421 THEN
            sigmoid_f := 2035;
        ELSIF x = 10422 THEN
            sigmoid_f := 2035;
        ELSIF x = 10423 THEN
            sigmoid_f := 2035;
        ELSIF x = 10424 THEN
            sigmoid_f := 2035;
        ELSIF x = 10425 THEN
            sigmoid_f := 2035;
        ELSIF x = 10426 THEN
            sigmoid_f := 2035;
        ELSIF x = 10427 THEN
            sigmoid_f := 2035;
        ELSIF x = 10428 THEN
            sigmoid_f := 2035;
        ELSIF x = 10429 THEN
            sigmoid_f := 2035;
        ELSIF x = 10430 THEN
            sigmoid_f := 2035;
        ELSIF x = 10431 THEN
            sigmoid_f := 2035;
        ELSIF x = 10432 THEN
            sigmoid_f := 2035;
        ELSIF x = 10433 THEN
            sigmoid_f := 2035;
        ELSIF x = 10434 THEN
            sigmoid_f := 2035;
        ELSIF x = 10435 THEN
            sigmoid_f := 2035;
        ELSIF x = 10436 THEN
            sigmoid_f := 2035;
        ELSIF x = 10437 THEN
            sigmoid_f := 2035;
        ELSIF x = 10438 THEN
            sigmoid_f := 2035;
        ELSIF x = 10439 THEN
            sigmoid_f := 2035;
        ELSIF x = 10440 THEN
            sigmoid_f := 2035;
        ELSIF x = 10441 THEN
            sigmoid_f := 2035;
        ELSIF x = 10442 THEN
            sigmoid_f := 2035;
        ELSIF x = 10443 THEN
            sigmoid_f := 2035;
        ELSIF x = 10444 THEN
            sigmoid_f := 2035;
        ELSIF x = 10445 THEN
            sigmoid_f := 2035;
        ELSIF x = 10446 THEN
            sigmoid_f := 2035;
        ELSIF x = 10447 THEN
            sigmoid_f := 2035;
        ELSIF x = 10448 THEN
            sigmoid_f := 2035;
        ELSIF x = 10449 THEN
            sigmoid_f := 2035;
        ELSIF x = 10450 THEN
            sigmoid_f := 2035;
        ELSIF x = 10451 THEN
            sigmoid_f := 2035;
        ELSIF x = 10452 THEN
            sigmoid_f := 2035;
        ELSIF x = 10453 THEN
            sigmoid_f := 2035;
        ELSIF x = 10454 THEN
            sigmoid_f := 2035;
        ELSIF x = 10455 THEN
            sigmoid_f := 2035;
        ELSIF x = 10456 THEN
            sigmoid_f := 2035;
        ELSIF x = 10457 THEN
            sigmoid_f := 2035;
        ELSIF x = 10458 THEN
            sigmoid_f := 2035;
        ELSIF x = 10459 THEN
            sigmoid_f := 2035;
        ELSIF x = 10460 THEN
            sigmoid_f := 2035;
        ELSIF x = 10461 THEN
            sigmoid_f := 2035;
        ELSIF x = 10462 THEN
            sigmoid_f := 2035;
        ELSIF x = 10463 THEN
            sigmoid_f := 2035;
        ELSIF x = 10464 THEN
            sigmoid_f := 2035;
        ELSIF x = 10465 THEN
            sigmoid_f := 2035;
        ELSIF x = 10466 THEN
            sigmoid_f := 2035;
        ELSIF x = 10467 THEN
            sigmoid_f := 2035;
        ELSIF x = 10468 THEN
            sigmoid_f := 2035;
        ELSIF x = 10469 THEN
            sigmoid_f := 2035;
        ELSIF x = 10470 THEN
            sigmoid_f := 2035;
        ELSIF x = 10471 THEN
            sigmoid_f := 2035;
        ELSIF x = 10472 THEN
            sigmoid_f := 2035;
        ELSIF x = 10473 THEN
            sigmoid_f := 2035;
        ELSIF x = 10474 THEN
            sigmoid_f := 2035;
        ELSIF x = 10475 THEN
            sigmoid_f := 2035;
        ELSIF x = 10476 THEN
            sigmoid_f := 2035;
        ELSIF x = 10477 THEN
            sigmoid_f := 2035;
        ELSIF x = 10478 THEN
            sigmoid_f := 2035;
        ELSIF x = 10479 THEN
            sigmoid_f := 2035;
        ELSIF x = 10480 THEN
            sigmoid_f := 2035;
        ELSIF x = 10481 THEN
            sigmoid_f := 2035;
        ELSIF x = 10482 THEN
            sigmoid_f := 2035;
        ELSIF x = 10483 THEN
            sigmoid_f := 2035;
        ELSIF x = 10484 THEN
            sigmoid_f := 2035;
        ELSIF x = 10485 THEN
            sigmoid_f := 2035;
        ELSIF x = 10486 THEN
            sigmoid_f := 2035;
        ELSIF x = 10487 THEN
            sigmoid_f := 2035;
        ELSIF x = 10488 THEN
            sigmoid_f := 2035;
        ELSIF x = 10489 THEN
            sigmoid_f := 2035;
        ELSIF x = 10490 THEN
            sigmoid_f := 2035;
        ELSIF x = 10491 THEN
            sigmoid_f := 2035;
        ELSIF x = 10492 THEN
            sigmoid_f := 2035;
        ELSIF x = 10493 THEN
            sigmoid_f := 2035;
        ELSIF x = 10494 THEN
            sigmoid_f := 2035;
        ELSIF x = 10495 THEN
            sigmoid_f := 2035;
        ELSIF x = 10496 THEN
            sigmoid_f := 2035;
        ELSIF x = 10497 THEN
            sigmoid_f := 2035;
        ELSIF x = 10498 THEN
            sigmoid_f := 2035;
        ELSIF x = 10499 THEN
            sigmoid_f := 2035;
        ELSIF x = 10500 THEN
            sigmoid_f := 2035;
        ELSIF x = 10501 THEN
            sigmoid_f := 2035;
        ELSIF x = 10502 THEN
            sigmoid_f := 2035;
        ELSIF x = 10503 THEN
            sigmoid_f := 2035;
        ELSIF x = 10504 THEN
            sigmoid_f := 2035;
        ELSIF x = 10505 THEN
            sigmoid_f := 2035;
        ELSIF x = 10506 THEN
            sigmoid_f := 2035;
        ELSIF x = 10507 THEN
            sigmoid_f := 2035;
        ELSIF x = 10508 THEN
            sigmoid_f := 2035;
        ELSIF x = 10509 THEN
            sigmoid_f := 2035;
        ELSIF x = 10510 THEN
            sigmoid_f := 2035;
        ELSIF x = 10511 THEN
            sigmoid_f := 2035;
        ELSIF x = 10512 THEN
            sigmoid_f := 2035;
        ELSIF x = 10513 THEN
            sigmoid_f := 2035;
        ELSIF x = 10514 THEN
            sigmoid_f := 2035;
        ELSIF x = 10515 THEN
            sigmoid_f := 2035;
        ELSIF x = 10516 THEN
            sigmoid_f := 2035;
        ELSIF x = 10517 THEN
            sigmoid_f := 2035;
        ELSIF x = 10518 THEN
            sigmoid_f := 2035;
        ELSIF x = 10519 THEN
            sigmoid_f := 2035;
        ELSIF x = 10520 THEN
            sigmoid_f := 2035;
        ELSIF x = 10521 THEN
            sigmoid_f := 2035;
        ELSIF x = 10522 THEN
            sigmoid_f := 2035;
        ELSIF x = 10523 THEN
            sigmoid_f := 2035;
        ELSIF x = 10524 THEN
            sigmoid_f := 2035;
        ELSIF x = 10525 THEN
            sigmoid_f := 2035;
        ELSIF x = 10526 THEN
            sigmoid_f := 2035;
        ELSIF x = 10527 THEN
            sigmoid_f := 2035;
        ELSIF x = 10528 THEN
            sigmoid_f := 2035;
        ELSIF x = 10529 THEN
            sigmoid_f := 2035;
        ELSIF x = 10530 THEN
            sigmoid_f := 2035;
        ELSIF x = 10531 THEN
            sigmoid_f := 2035;
        ELSIF x = 10532 THEN
            sigmoid_f := 2035;
        ELSIF x = 10533 THEN
            sigmoid_f := 2036;
        ELSIF x = 10534 THEN
            sigmoid_f := 2036;
        ELSIF x = 10535 THEN
            sigmoid_f := 2036;
        ELSIF x = 10536 THEN
            sigmoid_f := 2036;
        ELSIF x = 10537 THEN
            sigmoid_f := 2036;
        ELSIF x = 10538 THEN
            sigmoid_f := 2036;
        ELSIF x = 10539 THEN
            sigmoid_f := 2036;
        ELSIF x = 10540 THEN
            sigmoid_f := 2036;
        ELSIF x = 10541 THEN
            sigmoid_f := 2036;
        ELSIF x = 10542 THEN
            sigmoid_f := 2036;
        ELSIF x = 10543 THEN
            sigmoid_f := 2036;
        ELSIF x = 10544 THEN
            sigmoid_f := 2036;
        ELSIF x = 10545 THEN
            sigmoid_f := 2036;
        ELSIF x = 10546 THEN
            sigmoid_f := 2036;
        ELSIF x = 10547 THEN
            sigmoid_f := 2036;
        ELSIF x = 10548 THEN
            sigmoid_f := 2036;
        ELSIF x = 10549 THEN
            sigmoid_f := 2036;
        ELSIF x = 10550 THEN
            sigmoid_f := 2036;
        ELSIF x = 10551 THEN
            sigmoid_f := 2036;
        ELSIF x = 10552 THEN
            sigmoid_f := 2036;
        ELSIF x = 10553 THEN
            sigmoid_f := 2036;
        ELSIF x = 10554 THEN
            sigmoid_f := 2036;
        ELSIF x = 10555 THEN
            sigmoid_f := 2036;
        ELSIF x = 10556 THEN
            sigmoid_f := 2036;
        ELSIF x = 10557 THEN
            sigmoid_f := 2036;
        ELSIF x = 10558 THEN
            sigmoid_f := 2036;
        ELSIF x = 10559 THEN
            sigmoid_f := 2036;
        ELSIF x = 10560 THEN
            sigmoid_f := 2036;
        ELSIF x = 10561 THEN
            sigmoid_f := 2036;
        ELSIF x = 10562 THEN
            sigmoid_f := 2036;
        ELSIF x = 10563 THEN
            sigmoid_f := 2036;
        ELSIF x = 10564 THEN
            sigmoid_f := 2036;
        ELSIF x = 10565 THEN
            sigmoid_f := 2036;
        ELSIF x = 10566 THEN
            sigmoid_f := 2036;
        ELSIF x = 10567 THEN
            sigmoid_f := 2036;
        ELSIF x = 10568 THEN
            sigmoid_f := 2036;
        ELSIF x = 10569 THEN
            sigmoid_f := 2036;
        ELSIF x = 10570 THEN
            sigmoid_f := 2036;
        ELSIF x = 10571 THEN
            sigmoid_f := 2036;
        ELSIF x = 10572 THEN
            sigmoid_f := 2036;
        ELSIF x = 10573 THEN
            sigmoid_f := 2036;
        ELSIF x = 10574 THEN
            sigmoid_f := 2036;
        ELSIF x = 10575 THEN
            sigmoid_f := 2036;
        ELSIF x = 10576 THEN
            sigmoid_f := 2036;
        ELSIF x = 10577 THEN
            sigmoid_f := 2036;
        ELSIF x = 10578 THEN
            sigmoid_f := 2036;
        ELSIF x = 10579 THEN
            sigmoid_f := 2036;
        ELSIF x = 10580 THEN
            sigmoid_f := 2036;
        ELSIF x = 10581 THEN
            sigmoid_f := 2036;
        ELSIF x = 10582 THEN
            sigmoid_f := 2036;
        ELSIF x = 10583 THEN
            sigmoid_f := 2036;
        ELSIF x = 10584 THEN
            sigmoid_f := 2036;
        ELSIF x = 10585 THEN
            sigmoid_f := 2036;
        ELSIF x = 10586 THEN
            sigmoid_f := 2036;
        ELSIF x = 10587 THEN
            sigmoid_f := 2036;
        ELSIF x = 10588 THEN
            sigmoid_f := 2036;
        ELSIF x = 10589 THEN
            sigmoid_f := 2036;
        ELSIF x = 10590 THEN
            sigmoid_f := 2036;
        ELSIF x = 10591 THEN
            sigmoid_f := 2036;
        ELSIF x = 10592 THEN
            sigmoid_f := 2036;
        ELSIF x = 10593 THEN
            sigmoid_f := 2036;
        ELSIF x = 10594 THEN
            sigmoid_f := 2036;
        ELSIF x = 10595 THEN
            sigmoid_f := 2036;
        ELSIF x = 10596 THEN
            sigmoid_f := 2036;
        ELSIF x = 10597 THEN
            sigmoid_f := 2036;
        ELSIF x = 10598 THEN
            sigmoid_f := 2036;
        ELSIF x = 10599 THEN
            sigmoid_f := 2036;
        ELSIF x = 10600 THEN
            sigmoid_f := 2036;
        ELSIF x = 10601 THEN
            sigmoid_f := 2036;
        ELSIF x = 10602 THEN
            sigmoid_f := 2036;
        ELSIF x = 10603 THEN
            sigmoid_f := 2036;
        ELSIF x = 10604 THEN
            sigmoid_f := 2036;
        ELSIF x = 10605 THEN
            sigmoid_f := 2036;
        ELSIF x = 10606 THEN
            sigmoid_f := 2036;
        ELSIF x = 10607 THEN
            sigmoid_f := 2036;
        ELSIF x = 10608 THEN
            sigmoid_f := 2036;
        ELSIF x = 10609 THEN
            sigmoid_f := 2036;
        ELSIF x = 10610 THEN
            sigmoid_f := 2036;
        ELSIF x = 10611 THEN
            sigmoid_f := 2036;
        ELSIF x = 10612 THEN
            sigmoid_f := 2036;
        ELSIF x = 10613 THEN
            sigmoid_f := 2036;
        ELSIF x = 10614 THEN
            sigmoid_f := 2036;
        ELSIF x = 10615 THEN
            sigmoid_f := 2036;
        ELSIF x = 10616 THEN
            sigmoid_f := 2036;
        ELSIF x = 10617 THEN
            sigmoid_f := 2036;
        ELSIF x = 10618 THEN
            sigmoid_f := 2036;
        ELSIF x = 10619 THEN
            sigmoid_f := 2036;
        ELSIF x = 10620 THEN
            sigmoid_f := 2036;
        ELSIF x = 10621 THEN
            sigmoid_f := 2036;
        ELSIF x = 10622 THEN
            sigmoid_f := 2036;
        ELSIF x = 10623 THEN
            sigmoid_f := 2036;
        ELSIF x = 10624 THEN
            sigmoid_f := 2036;
        ELSIF x = 10625 THEN
            sigmoid_f := 2036;
        ELSIF x = 10626 THEN
            sigmoid_f := 2036;
        ELSIF x = 10627 THEN
            sigmoid_f := 2036;
        ELSIF x = 10628 THEN
            sigmoid_f := 2036;
        ELSIF x = 10629 THEN
            sigmoid_f := 2036;
        ELSIF x = 10630 THEN
            sigmoid_f := 2036;
        ELSIF x = 10631 THEN
            sigmoid_f := 2036;
        ELSIF x = 10632 THEN
            sigmoid_f := 2036;
        ELSIF x = 10633 THEN
            sigmoid_f := 2036;
        ELSIF x = 10634 THEN
            sigmoid_f := 2036;
        ELSIF x = 10635 THEN
            sigmoid_f := 2036;
        ELSIF x = 10636 THEN
            sigmoid_f := 2036;
        ELSIF x = 10637 THEN
            sigmoid_f := 2036;
        ELSIF x = 10638 THEN
            sigmoid_f := 2036;
        ELSIF x = 10639 THEN
            sigmoid_f := 2036;
        ELSIF x = 10640 THEN
            sigmoid_f := 2036;
        ELSIF x = 10641 THEN
            sigmoid_f := 2036;
        ELSIF x = 10642 THEN
            sigmoid_f := 2036;
        ELSIF x = 10643 THEN
            sigmoid_f := 2036;
        ELSIF x = 10644 THEN
            sigmoid_f := 2036;
        ELSIF x = 10645 THEN
            sigmoid_f := 2036;
        ELSIF x = 10646 THEN
            sigmoid_f := 2036;
        ELSIF x = 10647 THEN
            sigmoid_f := 2036;
        ELSIF x = 10648 THEN
            sigmoid_f := 2036;
        ELSIF x = 10649 THEN
            sigmoid_f := 2036;
        ELSIF x = 10650 THEN
            sigmoid_f := 2036;
        ELSIF x = 10651 THEN
            sigmoid_f := 2036;
        ELSIF x = 10652 THEN
            sigmoid_f := 2036;
        ELSIF x = 10653 THEN
            sigmoid_f := 2036;
        ELSIF x = 10654 THEN
            sigmoid_f := 2036;
        ELSIF x = 10655 THEN
            sigmoid_f := 2036;
        ELSIF x = 10656 THEN
            sigmoid_f := 2036;
        ELSIF x = 10657 THEN
            sigmoid_f := 2036;
        ELSIF x = 10658 THEN
            sigmoid_f := 2036;
        ELSIF x = 10659 THEN
            sigmoid_f := 2036;
        ELSIF x = 10660 THEN
            sigmoid_f := 2036;
        ELSIF x = 10661 THEN
            sigmoid_f := 2036;
        ELSIF x = 10662 THEN
            sigmoid_f := 2036;
        ELSIF x = 10663 THEN
            sigmoid_f := 2036;
        ELSIF x = 10664 THEN
            sigmoid_f := 2036;
        ELSIF x = 10665 THEN
            sigmoid_f := 2036;
        ELSIF x = 10666 THEN
            sigmoid_f := 2036;
        ELSIF x = 10667 THEN
            sigmoid_f := 2036;
        ELSIF x = 10668 THEN
            sigmoid_f := 2036;
        ELSIF x = 10669 THEN
            sigmoid_f := 2036;
        ELSIF x = 10670 THEN
            sigmoid_f := 2036;
        ELSIF x = 10671 THEN
            sigmoid_f := 2036;
        ELSIF x = 10672 THEN
            sigmoid_f := 2036;
        ELSIF x = 10673 THEN
            sigmoid_f := 2036;
        ELSIF x = 10674 THEN
            sigmoid_f := 2036;
        ELSIF x = 10675 THEN
            sigmoid_f := 2036;
        ELSIF x = 10676 THEN
            sigmoid_f := 2036;
        ELSIF x = 10677 THEN
            sigmoid_f := 2036;
        ELSIF x = 10678 THEN
            sigmoid_f := 2036;
        ELSIF x = 10679 THEN
            sigmoid_f := 2037;
        ELSIF x = 10680 THEN
            sigmoid_f := 2037;
        ELSIF x = 10681 THEN
            sigmoid_f := 2037;
        ELSIF x = 10682 THEN
            sigmoid_f := 2037;
        ELSIF x = 10683 THEN
            sigmoid_f := 2037;
        ELSIF x = 10684 THEN
            sigmoid_f := 2037;
        ELSIF x = 10685 THEN
            sigmoid_f := 2037;
        ELSIF x = 10686 THEN
            sigmoid_f := 2037;
        ELSIF x = 10687 THEN
            sigmoid_f := 2037;
        ELSIF x = 10688 THEN
            sigmoid_f := 2037;
        ELSIF x = 10689 THEN
            sigmoid_f := 2037;
        ELSIF x = 10690 THEN
            sigmoid_f := 2037;
        ELSIF x = 10691 THEN
            sigmoid_f := 2037;
        ELSIF x = 10692 THEN
            sigmoid_f := 2037;
        ELSIF x = 10693 THEN
            sigmoid_f := 2037;
        ELSIF x = 10694 THEN
            sigmoid_f := 2037;
        ELSIF x = 10695 THEN
            sigmoid_f := 2037;
        ELSIF x = 10696 THEN
            sigmoid_f := 2037;
        ELSIF x = 10697 THEN
            sigmoid_f := 2037;
        ELSIF x = 10698 THEN
            sigmoid_f := 2037;
        ELSIF x = 10699 THEN
            sigmoid_f := 2037;
        ELSIF x = 10700 THEN
            sigmoid_f := 2037;
        ELSIF x = 10701 THEN
            sigmoid_f := 2037;
        ELSIF x = 10702 THEN
            sigmoid_f := 2037;
        ELSIF x = 10703 THEN
            sigmoid_f := 2037;
        ELSIF x = 10704 THEN
            sigmoid_f := 2037;
        ELSIF x = 10705 THEN
            sigmoid_f := 2037;
        ELSIF x = 10706 THEN
            sigmoid_f := 2037;
        ELSIF x = 10707 THEN
            sigmoid_f := 2037;
        ELSIF x = 10708 THEN
            sigmoid_f := 2037;
        ELSIF x = 10709 THEN
            sigmoid_f := 2037;
        ELSIF x = 10710 THEN
            sigmoid_f := 2037;
        ELSIF x = 10711 THEN
            sigmoid_f := 2037;
        ELSIF x = 10712 THEN
            sigmoid_f := 2037;
        ELSIF x = 10713 THEN
            sigmoid_f := 2037;
        ELSIF x = 10714 THEN
            sigmoid_f := 2037;
        ELSIF x = 10715 THEN
            sigmoid_f := 2037;
        ELSIF x = 10716 THEN
            sigmoid_f := 2037;
        ELSIF x = 10717 THEN
            sigmoid_f := 2037;
        ELSIF x = 10718 THEN
            sigmoid_f := 2037;
        ELSIF x = 10719 THEN
            sigmoid_f := 2037;
        ELSIF x = 10720 THEN
            sigmoid_f := 2037;
        ELSIF x = 10721 THEN
            sigmoid_f := 2037;
        ELSIF x = 10722 THEN
            sigmoid_f := 2037;
        ELSIF x = 10723 THEN
            sigmoid_f := 2037;
        ELSIF x = 10724 THEN
            sigmoid_f := 2037;
        ELSIF x = 10725 THEN
            sigmoid_f := 2037;
        ELSIF x = 10726 THEN
            sigmoid_f := 2037;
        ELSIF x = 10727 THEN
            sigmoid_f := 2037;
        ELSIF x = 10728 THEN
            sigmoid_f := 2037;
        ELSIF x = 10729 THEN
            sigmoid_f := 2037;
        ELSIF x = 10730 THEN
            sigmoid_f := 2037;
        ELSIF x = 10731 THEN
            sigmoid_f := 2037;
        ELSIF x = 10732 THEN
            sigmoid_f := 2037;
        ELSIF x = 10733 THEN
            sigmoid_f := 2037;
        ELSIF x = 10734 THEN
            sigmoid_f := 2037;
        ELSIF x = 10735 THEN
            sigmoid_f := 2037;
        ELSIF x = 10736 THEN
            sigmoid_f := 2037;
        ELSIF x = 10737 THEN
            sigmoid_f := 2037;
        ELSIF x = 10738 THEN
            sigmoid_f := 2037;
        ELSIF x = 10739 THEN
            sigmoid_f := 2037;
        ELSIF x = 10740 THEN
            sigmoid_f := 2037;
        ELSIF x = 10741 THEN
            sigmoid_f := 2037;
        ELSIF x = 10742 THEN
            sigmoid_f := 2037;
        ELSIF x = 10743 THEN
            sigmoid_f := 2037;
        ELSIF x = 10744 THEN
            sigmoid_f := 2037;
        ELSIF x = 10745 THEN
            sigmoid_f := 2037;
        ELSIF x = 10746 THEN
            sigmoid_f := 2037;
        ELSIF x = 10747 THEN
            sigmoid_f := 2037;
        ELSIF x = 10748 THEN
            sigmoid_f := 2037;
        ELSIF x = 10749 THEN
            sigmoid_f := 2037;
        ELSIF x = 10750 THEN
            sigmoid_f := 2037;
        ELSIF x = 10751 THEN
            sigmoid_f := 2037;
        ELSIF x = 10752 THEN
            sigmoid_f := 2037;
        ELSIF x = 10753 THEN
            sigmoid_f := 2037;
        ELSIF x = 10754 THEN
            sigmoid_f := 2037;
        ELSIF x = 10755 THEN
            sigmoid_f := 2037;
        ELSIF x = 10756 THEN
            sigmoid_f := 2037;
        ELSIF x = 10757 THEN
            sigmoid_f := 2037;
        ELSIF x = 10758 THEN
            sigmoid_f := 2037;
        ELSIF x = 10759 THEN
            sigmoid_f := 2037;
        ELSIF x = 10760 THEN
            sigmoid_f := 2037;
        ELSIF x = 10761 THEN
            sigmoid_f := 2037;
        ELSIF x = 10762 THEN
            sigmoid_f := 2037;
        ELSIF x = 10763 THEN
            sigmoid_f := 2037;
        ELSIF x = 10764 THEN
            sigmoid_f := 2037;
        ELSIF x = 10765 THEN
            sigmoid_f := 2037;
        ELSIF x = 10766 THEN
            sigmoid_f := 2037;
        ELSIF x = 10767 THEN
            sigmoid_f := 2037;
        ELSIF x = 10768 THEN
            sigmoid_f := 2037;
        ELSIF x = 10769 THEN
            sigmoid_f := 2037;
        ELSIF x = 10770 THEN
            sigmoid_f := 2037;
        ELSIF x = 10771 THEN
            sigmoid_f := 2037;
        ELSIF x = 10772 THEN
            sigmoid_f := 2037;
        ELSIF x = 10773 THEN
            sigmoid_f := 2037;
        ELSIF x = 10774 THEN
            sigmoid_f := 2037;
        ELSIF x = 10775 THEN
            sigmoid_f := 2037;
        ELSIF x = 10776 THEN
            sigmoid_f := 2037;
        ELSIF x = 10777 THEN
            sigmoid_f := 2037;
        ELSIF x = 10778 THEN
            sigmoid_f := 2037;
        ELSIF x = 10779 THEN
            sigmoid_f := 2037;
        ELSIF x = 10780 THEN
            sigmoid_f := 2037;
        ELSIF x = 10781 THEN
            sigmoid_f := 2037;
        ELSIF x = 10782 THEN
            sigmoid_f := 2037;
        ELSIF x = 10783 THEN
            sigmoid_f := 2037;
        ELSIF x = 10784 THEN
            sigmoid_f := 2037;
        ELSIF x = 10785 THEN
            sigmoid_f := 2037;
        ELSIF x = 10786 THEN
            sigmoid_f := 2037;
        ELSIF x = 10787 THEN
            sigmoid_f := 2037;
        ELSIF x = 10788 THEN
            sigmoid_f := 2037;
        ELSIF x = 10789 THEN
            sigmoid_f := 2037;
        ELSIF x = 10790 THEN
            sigmoid_f := 2037;
        ELSIF x = 10791 THEN
            sigmoid_f := 2037;
        ELSIF x = 10792 THEN
            sigmoid_f := 2037;
        ELSIF x = 10793 THEN
            sigmoid_f := 2037;
        ELSIF x = 10794 THEN
            sigmoid_f := 2037;
        ELSIF x = 10795 THEN
            sigmoid_f := 2037;
        ELSIF x = 10796 THEN
            sigmoid_f := 2037;
        ELSIF x = 10797 THEN
            sigmoid_f := 2037;
        ELSIF x = 10798 THEN
            sigmoid_f := 2037;
        ELSIF x = 10799 THEN
            sigmoid_f := 2037;
        ELSIF x = 10800 THEN
            sigmoid_f := 2037;
        ELSIF x = 10801 THEN
            sigmoid_f := 2037;
        ELSIF x = 10802 THEN
            sigmoid_f := 2037;
        ELSIF x = 10803 THEN
            sigmoid_f := 2037;
        ELSIF x = 10804 THEN
            sigmoid_f := 2037;
        ELSIF x = 10805 THEN
            sigmoid_f := 2037;
        ELSIF x = 10806 THEN
            sigmoid_f := 2037;
        ELSIF x = 10807 THEN
            sigmoid_f := 2037;
        ELSIF x = 10808 THEN
            sigmoid_f := 2037;
        ELSIF x = 10809 THEN
            sigmoid_f := 2037;
        ELSIF x = 10810 THEN
            sigmoid_f := 2037;
        ELSIF x = 10811 THEN
            sigmoid_f := 2037;
        ELSIF x = 10812 THEN
            sigmoid_f := 2037;
        ELSIF x = 10813 THEN
            sigmoid_f := 2037;
        ELSIF x = 10814 THEN
            sigmoid_f := 2037;
        ELSIF x = 10815 THEN
            sigmoid_f := 2037;
        ELSIF x = 10816 THEN
            sigmoid_f := 2037;
        ELSIF x = 10817 THEN
            sigmoid_f := 2037;
        ELSIF x = 10818 THEN
            sigmoid_f := 2037;
        ELSIF x = 10819 THEN
            sigmoid_f := 2037;
        ELSIF x = 10820 THEN
            sigmoid_f := 2037;
        ELSIF x = 10821 THEN
            sigmoid_f := 2037;
        ELSIF x = 10822 THEN
            sigmoid_f := 2037;
        ELSIF x = 10823 THEN
            sigmoid_f := 2037;
        ELSIF x = 10824 THEN
            sigmoid_f := 2037;
        ELSIF x = 10825 THEN
            sigmoid_f := 2037;
        ELSIF x = 10826 THEN
            sigmoid_f := 2037;
        ELSIF x = 10827 THEN
            sigmoid_f := 2037;
        ELSIF x = 10828 THEN
            sigmoid_f := 2037;
        ELSIF x = 10829 THEN
            sigmoid_f := 2037;
        ELSIF x = 10830 THEN
            sigmoid_f := 2037;
        ELSIF x = 10831 THEN
            sigmoid_f := 2037;
        ELSIF x = 10832 THEN
            sigmoid_f := 2037;
        ELSIF x = 10833 THEN
            sigmoid_f := 2037;
        ELSIF x = 10834 THEN
            sigmoid_f := 2037;
        ELSIF x = 10835 THEN
            sigmoid_f := 2037;
        ELSIF x = 10836 THEN
            sigmoid_f := 2037;
        ELSIF x = 10837 THEN
            sigmoid_f := 2037;
        ELSIF x = 10838 THEN
            sigmoid_f := 2037;
        ELSIF x = 10839 THEN
            sigmoid_f := 2037;
        ELSIF x = 10840 THEN
            sigmoid_f := 2037;
        ELSIF x = 10841 THEN
            sigmoid_f := 2037;
        ELSIF x = 10842 THEN
            sigmoid_f := 2037;
        ELSIF x = 10843 THEN
            sigmoid_f := 2037;
        ELSIF x = 10844 THEN
            sigmoid_f := 2037;
        ELSIF x = 10845 THEN
            sigmoid_f := 2037;
        ELSIF x = 10846 THEN
            sigmoid_f := 2037;
        ELSIF x = 10847 THEN
            sigmoid_f := 2037;
        ELSIF x = 10848 THEN
            sigmoid_f := 2037;
        ELSIF x = 10849 THEN
            sigmoid_f := 2037;
        ELSIF x = 10850 THEN
            sigmoid_f := 2037;
        ELSIF x = 10851 THEN
            sigmoid_f := 2037;
        ELSIF x = 10852 THEN
            sigmoid_f := 2037;
        ELSIF x = 10853 THEN
            sigmoid_f := 2037;
        ELSIF x = 10854 THEN
            sigmoid_f := 2037;
        ELSIF x = 10855 THEN
            sigmoid_f := 2037;
        ELSIF x = 10856 THEN
            sigmoid_f := 2037;
        ELSIF x = 10857 THEN
            sigmoid_f := 2037;
        ELSIF x = 10858 THEN
            sigmoid_f := 2037;
        ELSIF x = 10859 THEN
            sigmoid_f := 2037;
        ELSIF x = 10860 THEN
            sigmoid_f := 2037;
        ELSIF x = 10861 THEN
            sigmoid_f := 2037;
        ELSIF x = 10862 THEN
            sigmoid_f := 2037;
        ELSIF x = 10863 THEN
            sigmoid_f := 2037;
        ELSIF x = 10864 THEN
            sigmoid_f := 2037;
        ELSIF x = 10865 THEN
            sigmoid_f := 2037;
        ELSIF x = 10866 THEN
            sigmoid_f := 2037;
        ELSIF x = 10867 THEN
            sigmoid_f := 2037;
        ELSIF x = 10868 THEN
            sigmoid_f := 2037;
        ELSIF x = 10869 THEN
            sigmoid_f := 2037;
        ELSIF x = 10870 THEN
            sigmoid_f := 2037;
        ELSIF x = 10871 THEN
            sigmoid_f := 2037;
        ELSIF x = 10872 THEN
            sigmoid_f := 2037;
        ELSIF x = 10873 THEN
            sigmoid_f := 2037;
        ELSIF x = 10874 THEN
            sigmoid_f := 2037;
        ELSIF x = 10875 THEN
            sigmoid_f := 2037;
        ELSIF x = 10876 THEN
            sigmoid_f := 2037;
        ELSIF x = 10877 THEN
            sigmoid_f := 2037;
        ELSIF x = 10878 THEN
            sigmoid_f := 2037;
        ELSIF x = 10879 THEN
            sigmoid_f := 2037;
        ELSIF x = 10880 THEN
            sigmoid_f := 2037;
        ELSIF x = 10881 THEN
            sigmoid_f := 2037;
        ELSIF x = 10882 THEN
            sigmoid_f := 2037;
        ELSIF x = 10883 THEN
            sigmoid_f := 2037;
        ELSIF x = 10884 THEN
            sigmoid_f := 2037;
        ELSIF x = 10885 THEN
            sigmoid_f := 2037;
        ELSIF x = 10886 THEN
            sigmoid_f := 2037;
        ELSIF x = 10887 THEN
            sigmoid_f := 2037;
        ELSIF x = 10888 THEN
            sigmoid_f := 2037;
        ELSIF x = 10889 THEN
            sigmoid_f := 2037;
        ELSIF x = 10890 THEN
            sigmoid_f := 2037;
        ELSIF x = 10891 THEN
            sigmoid_f := 2037;
        ELSIF x = 10892 THEN
            sigmoid_f := 2037;
        ELSIF x = 10893 THEN
            sigmoid_f := 2037;
        ELSIF x = 10894 THEN
            sigmoid_f := 2037;
        ELSIF x = 10895 THEN
            sigmoid_f := 2037;
        ELSIF x = 10896 THEN
            sigmoid_f := 2037;
        ELSIF x = 10897 THEN
            sigmoid_f := 2037;
        ELSIF x = 10898 THEN
            sigmoid_f := 2037;
        ELSIF x = 10899 THEN
            sigmoid_f := 2037;
        ELSIF x = 10900 THEN
            sigmoid_f := 2037;
        ELSIF x = 10901 THEN
            sigmoid_f := 2037;
        ELSIF x = 10902 THEN
            sigmoid_f := 2037;
        ELSIF x = 10903 THEN
            sigmoid_f := 2037;
        ELSIF x = 10904 THEN
            sigmoid_f := 2037;
        ELSIF x = 10905 THEN
            sigmoid_f := 2037;
        ELSIF x = 10906 THEN
            sigmoid_f := 2037;
        ELSIF x = 10907 THEN
            sigmoid_f := 2037;
        ELSIF x = 10908 THEN
            sigmoid_f := 2037;
        ELSIF x = 10909 THEN
            sigmoid_f := 2037;
        ELSIF x = 10910 THEN
            sigmoid_f := 2037;
        ELSIF x = 10911 THEN
            sigmoid_f := 2037;
        ELSIF x = 10912 THEN
            sigmoid_f := 2037;
        ELSIF x = 10913 THEN
            sigmoid_f := 2037;
        ELSIF x = 10914 THEN
            sigmoid_f := 2037;
        ELSIF x = 10915 THEN
            sigmoid_f := 2037;
        ELSIF x = 10916 THEN
            sigmoid_f := 2037;
        ELSIF x = 10917 THEN
            sigmoid_f := 2037;
        ELSIF x = 10918 THEN
            sigmoid_f := 2037;
        ELSIF x = 10919 THEN
            sigmoid_f := 2037;
        ELSIF x = 10920 THEN
            sigmoid_f := 2037;
        ELSIF x = 10921 THEN
            sigmoid_f := 2037;
        ELSIF x = 10922 THEN
            sigmoid_f := 2037;
        ELSIF x = 10923 THEN
            sigmoid_f := 2038;
        ELSIF x = 10924 THEN
            sigmoid_f := 2038;
        ELSIF x = 10925 THEN
            sigmoid_f := 2038;
        ELSIF x = 10926 THEN
            sigmoid_f := 2038;
        ELSIF x = 10927 THEN
            sigmoid_f := 2038;
        ELSIF x = 10928 THEN
            sigmoid_f := 2038;
        ELSIF x = 10929 THEN
            sigmoid_f := 2038;
        ELSIF x = 10930 THEN
            sigmoid_f := 2038;
        ELSIF x = 10931 THEN
            sigmoid_f := 2038;
        ELSIF x = 10932 THEN
            sigmoid_f := 2038;
        ELSIF x = 10933 THEN
            sigmoid_f := 2038;
        ELSIF x = 10934 THEN
            sigmoid_f := 2038;
        ELSIF x = 10935 THEN
            sigmoid_f := 2038;
        ELSIF x = 10936 THEN
            sigmoid_f := 2038;
        ELSIF x = 10937 THEN
            sigmoid_f := 2038;
        ELSIF x = 10938 THEN
            sigmoid_f := 2038;
        ELSIF x = 10939 THEN
            sigmoid_f := 2038;
        ELSIF x = 10940 THEN
            sigmoid_f := 2038;
        ELSIF x = 10941 THEN
            sigmoid_f := 2038;
        ELSIF x = 10942 THEN
            sigmoid_f := 2038;
        ELSIF x = 10943 THEN
            sigmoid_f := 2038;
        ELSIF x = 10944 THEN
            sigmoid_f := 2038;
        ELSIF x = 10945 THEN
            sigmoid_f := 2038;
        ELSIF x = 10946 THEN
            sigmoid_f := 2038;
        ELSIF x = 10947 THEN
            sigmoid_f := 2038;
        ELSIF x = 10948 THEN
            sigmoid_f := 2038;
        ELSIF x = 10949 THEN
            sigmoid_f := 2038;
        ELSIF x = 10950 THEN
            sigmoid_f := 2038;
        ELSIF x = 10951 THEN
            sigmoid_f := 2038;
        ELSIF x = 10952 THEN
            sigmoid_f := 2038;
        ELSIF x = 10953 THEN
            sigmoid_f := 2038;
        ELSIF x = 10954 THEN
            sigmoid_f := 2038;
        ELSIF x = 10955 THEN
            sigmoid_f := 2038;
        ELSIF x = 10956 THEN
            sigmoid_f := 2038;
        ELSIF x = 10957 THEN
            sigmoid_f := 2038;
        ELSIF x = 10958 THEN
            sigmoid_f := 2038;
        ELSIF x = 10959 THEN
            sigmoid_f := 2038;
        ELSIF x = 10960 THEN
            sigmoid_f := 2038;
        ELSIF x = 10961 THEN
            sigmoid_f := 2038;
        ELSIF x = 10962 THEN
            sigmoid_f := 2038;
        ELSIF x = 10963 THEN
            sigmoid_f := 2038;
        ELSIF x = 10964 THEN
            sigmoid_f := 2038;
        ELSIF x = 10965 THEN
            sigmoid_f := 2038;
        ELSIF x = 10966 THEN
            sigmoid_f := 2038;
        ELSIF x = 10967 THEN
            sigmoid_f := 2038;
        ELSIF x = 10968 THEN
            sigmoid_f := 2038;
        ELSIF x = 10969 THEN
            sigmoid_f := 2038;
        ELSIF x = 10970 THEN
            sigmoid_f := 2038;
        ELSIF x = 10971 THEN
            sigmoid_f := 2038;
        ELSIF x = 10972 THEN
            sigmoid_f := 2038;
        ELSIF x = 10973 THEN
            sigmoid_f := 2038;
        ELSIF x = 10974 THEN
            sigmoid_f := 2038;
        ELSIF x = 10975 THEN
            sigmoid_f := 2038;
        ELSIF x = 10976 THEN
            sigmoid_f := 2038;
        ELSIF x = 10977 THEN
            sigmoid_f := 2038;
        ELSIF x = 10978 THEN
            sigmoid_f := 2038;
        ELSIF x = 10979 THEN
            sigmoid_f := 2038;
        ELSIF x = 10980 THEN
            sigmoid_f := 2038;
        ELSIF x = 10981 THEN
            sigmoid_f := 2038;
        ELSIF x = 10982 THEN
            sigmoid_f := 2038;
        ELSIF x = 10983 THEN
            sigmoid_f := 2038;
        ELSIF x = 10984 THEN
            sigmoid_f := 2038;
        ELSIF x = 10985 THEN
            sigmoid_f := 2038;
        ELSIF x = 10986 THEN
            sigmoid_f := 2038;
        ELSIF x = 10987 THEN
            sigmoid_f := 2038;
        ELSIF x = 10988 THEN
            sigmoid_f := 2038;
        ELSIF x = 10989 THEN
            sigmoid_f := 2038;
        ELSIF x = 10990 THEN
            sigmoid_f := 2038;
        ELSIF x = 10991 THEN
            sigmoid_f := 2038;
        ELSIF x = 10992 THEN
            sigmoid_f := 2038;
        ELSIF x = 10993 THEN
            sigmoid_f := 2038;
        ELSIF x = 10994 THEN
            sigmoid_f := 2038;
        ELSIF x = 10995 THEN
            sigmoid_f := 2038;
        ELSIF x = 10996 THEN
            sigmoid_f := 2038;
        ELSIF x = 10997 THEN
            sigmoid_f := 2038;
        ELSIF x = 10998 THEN
            sigmoid_f := 2038;
        ELSIF x = 10999 THEN
            sigmoid_f := 2038;
        ELSIF x = 11000 THEN
            sigmoid_f := 2038;
        ELSIF x = 11001 THEN
            sigmoid_f := 2038;
        ELSIF x = 11002 THEN
            sigmoid_f := 2038;
        ELSIF x = 11003 THEN
            sigmoid_f := 2038;
        ELSIF x = 11004 THEN
            sigmoid_f := 2038;
        ELSIF x = 11005 THEN
            sigmoid_f := 2038;
        ELSIF x = 11006 THEN
            sigmoid_f := 2038;
        ELSIF x = 11007 THEN
            sigmoid_f := 2038;
        ELSIF x = 11008 THEN
            sigmoid_f := 2038;
        ELSIF x = 11009 THEN
            sigmoid_f := 2038;
        ELSIF x = 11010 THEN
            sigmoid_f := 2038;
        ELSIF x = 11011 THEN
            sigmoid_f := 2038;
        ELSIF x = 11012 THEN
            sigmoid_f := 2038;
        ELSIF x = 11013 THEN
            sigmoid_f := 2038;
        ELSIF x = 11014 THEN
            sigmoid_f := 2038;
        ELSIF x = 11015 THEN
            sigmoid_f := 2038;
        ELSIF x = 11016 THEN
            sigmoid_f := 2038;
        ELSIF x = 11017 THEN
            sigmoid_f := 2038;
        ELSIF x = 11018 THEN
            sigmoid_f := 2038;
        ELSIF x = 11019 THEN
            sigmoid_f := 2038;
        ELSIF x = 11020 THEN
            sigmoid_f := 2038;
        ELSIF x = 11021 THEN
            sigmoid_f := 2038;
        ELSIF x = 11022 THEN
            sigmoid_f := 2038;
        ELSIF x = 11023 THEN
            sigmoid_f := 2038;
        ELSIF x = 11024 THEN
            sigmoid_f := 2038;
        ELSIF x = 11025 THEN
            sigmoid_f := 2038;
        ELSIF x = 11026 THEN
            sigmoid_f := 2038;
        ELSIF x = 11027 THEN
            sigmoid_f := 2038;
        ELSIF x = 11028 THEN
            sigmoid_f := 2038;
        ELSIF x = 11029 THEN
            sigmoid_f := 2038;
        ELSIF x = 11030 THEN
            sigmoid_f := 2038;
        ELSIF x = 11031 THEN
            sigmoid_f := 2038;
        ELSIF x = 11032 THEN
            sigmoid_f := 2038;
        ELSIF x = 11033 THEN
            sigmoid_f := 2038;
        ELSIF x = 11034 THEN
            sigmoid_f := 2038;
        ELSIF x = 11035 THEN
            sigmoid_f := 2038;
        ELSIF x = 11036 THEN
            sigmoid_f := 2038;
        ELSIF x = 11037 THEN
            sigmoid_f := 2038;
        ELSIF x = 11038 THEN
            sigmoid_f := 2038;
        ELSIF x = 11039 THEN
            sigmoid_f := 2038;
        ELSIF x = 11040 THEN
            sigmoid_f := 2038;
        ELSIF x = 11041 THEN
            sigmoid_f := 2038;
        ELSIF x = 11042 THEN
            sigmoid_f := 2038;
        ELSIF x = 11043 THEN
            sigmoid_f := 2038;
        ELSIF x = 11044 THEN
            sigmoid_f := 2038;
        ELSIF x = 11045 THEN
            sigmoid_f := 2038;
        ELSIF x = 11046 THEN
            sigmoid_f := 2038;
        ELSIF x = 11047 THEN
            sigmoid_f := 2038;
        ELSIF x = 11048 THEN
            sigmoid_f := 2038;
        ELSIF x = 11049 THEN
            sigmoid_f := 2038;
        ELSIF x = 11050 THEN
            sigmoid_f := 2038;
        ELSIF x = 11051 THEN
            sigmoid_f := 2038;
        ELSIF x = 11052 THEN
            sigmoid_f := 2038;
        ELSIF x = 11053 THEN
            sigmoid_f := 2038;
        ELSIF x = 11054 THEN
            sigmoid_f := 2038;
        ELSIF x = 11055 THEN
            sigmoid_f := 2038;
        ELSIF x = 11056 THEN
            sigmoid_f := 2038;
        ELSIF x = 11057 THEN
            sigmoid_f := 2038;
        ELSIF x = 11058 THEN
            sigmoid_f := 2038;
        ELSIF x = 11059 THEN
            sigmoid_f := 2038;
        ELSIF x = 11060 THEN
            sigmoid_f := 2038;
        ELSIF x = 11061 THEN
            sigmoid_f := 2038;
        ELSIF x = 11062 THEN
            sigmoid_f := 2038;
        ELSIF x = 11063 THEN
            sigmoid_f := 2038;
        ELSIF x = 11064 THEN
            sigmoid_f := 2038;
        ELSIF x = 11065 THEN
            sigmoid_f := 2038;
        ELSIF x = 11066 THEN
            sigmoid_f := 2038;
        ELSIF x = 11067 THEN
            sigmoid_f := 2038;
        ELSIF x = 11068 THEN
            sigmoid_f := 2038;
        ELSIF x = 11069 THEN
            sigmoid_f := 2038;
        ELSIF x = 11070 THEN
            sigmoid_f := 2038;
        ELSIF x = 11071 THEN
            sigmoid_f := 2038;
        ELSIF x = 11072 THEN
            sigmoid_f := 2038;
        ELSIF x = 11073 THEN
            sigmoid_f := 2038;
        ELSIF x = 11074 THEN
            sigmoid_f := 2038;
        ELSIF x = 11075 THEN
            sigmoid_f := 2038;
        ELSIF x = 11076 THEN
            sigmoid_f := 2038;
        ELSIF x = 11077 THEN
            sigmoid_f := 2038;
        ELSIF x = 11078 THEN
            sigmoid_f := 2038;
        ELSIF x = 11079 THEN
            sigmoid_f := 2038;
        ELSIF x = 11080 THEN
            sigmoid_f := 2038;
        ELSIF x = 11081 THEN
            sigmoid_f := 2038;
        ELSIF x = 11082 THEN
            sigmoid_f := 2038;
        ELSIF x = 11083 THEN
            sigmoid_f := 2038;
        ELSIF x = 11084 THEN
            sigmoid_f := 2038;
        ELSIF x = 11085 THEN
            sigmoid_f := 2038;
        ELSIF x = 11086 THEN
            sigmoid_f := 2038;
        ELSIF x = 11087 THEN
            sigmoid_f := 2038;
        ELSIF x = 11088 THEN
            sigmoid_f := 2038;
        ELSIF x = 11089 THEN
            sigmoid_f := 2038;
        ELSIF x = 11090 THEN
            sigmoid_f := 2038;
        ELSIF x = 11091 THEN
            sigmoid_f := 2038;
        ELSIF x = 11092 THEN
            sigmoid_f := 2038;
        ELSIF x = 11093 THEN
            sigmoid_f := 2038;
        ELSIF x = 11094 THEN
            sigmoid_f := 2039;
        ELSIF x = 11095 THEN
            sigmoid_f := 2039;
        ELSIF x = 11096 THEN
            sigmoid_f := 2039;
        ELSIF x = 11097 THEN
            sigmoid_f := 2039;
        ELSIF x = 11098 THEN
            sigmoid_f := 2039;
        ELSIF x = 11099 THEN
            sigmoid_f := 2039;
        ELSIF x = 11100 THEN
            sigmoid_f := 2039;
        ELSIF x = 11101 THEN
            sigmoid_f := 2039;
        ELSIF x = 11102 THEN
            sigmoid_f := 2039;
        ELSIF x = 11103 THEN
            sigmoid_f := 2039;
        ELSIF x = 11104 THEN
            sigmoid_f := 2039;
        ELSIF x = 11105 THEN
            sigmoid_f := 2039;
        ELSIF x = 11106 THEN
            sigmoid_f := 2039;
        ELSIF x = 11107 THEN
            sigmoid_f := 2039;
        ELSIF x = 11108 THEN
            sigmoid_f := 2039;
        ELSIF x = 11109 THEN
            sigmoid_f := 2039;
        ELSIF x = 11110 THEN
            sigmoid_f := 2039;
        ELSIF x = 11111 THEN
            sigmoid_f := 2039;
        ELSIF x = 11112 THEN
            sigmoid_f := 2039;
        ELSIF x = 11113 THEN
            sigmoid_f := 2039;
        ELSIF x = 11114 THEN
            sigmoid_f := 2039;
        ELSIF x = 11115 THEN
            sigmoid_f := 2039;
        ELSIF x = 11116 THEN
            sigmoid_f := 2039;
        ELSIF x = 11117 THEN
            sigmoid_f := 2039;
        ELSIF x = 11118 THEN
            sigmoid_f := 2039;
        ELSIF x = 11119 THEN
            sigmoid_f := 2039;
        ELSIF x = 11120 THEN
            sigmoid_f := 2039;
        ELSIF x = 11121 THEN
            sigmoid_f := 2039;
        ELSIF x = 11122 THEN
            sigmoid_f := 2039;
        ELSIF x = 11123 THEN
            sigmoid_f := 2039;
        ELSIF x = 11124 THEN
            sigmoid_f := 2039;
        ELSIF x = 11125 THEN
            sigmoid_f := 2039;
        ELSIF x = 11126 THEN
            sigmoid_f := 2039;
        ELSIF x = 11127 THEN
            sigmoid_f := 2039;
        ELSIF x = 11128 THEN
            sigmoid_f := 2039;
        ELSIF x = 11129 THEN
            sigmoid_f := 2039;
        ELSIF x = 11130 THEN
            sigmoid_f := 2039;
        ELSIF x = 11131 THEN
            sigmoid_f := 2039;
        ELSIF x = 11132 THEN
            sigmoid_f := 2039;
        ELSIF x = 11133 THEN
            sigmoid_f := 2039;
        ELSIF x = 11134 THEN
            sigmoid_f := 2039;
        ELSIF x = 11135 THEN
            sigmoid_f := 2039;
        ELSIF x = 11136 THEN
            sigmoid_f := 2039;
        ELSIF x = 11137 THEN
            sigmoid_f := 2039;
        ELSIF x = 11138 THEN
            sigmoid_f := 2039;
        ELSIF x = 11139 THEN
            sigmoid_f := 2039;
        ELSIF x = 11140 THEN
            sigmoid_f := 2039;
        ELSIF x = 11141 THEN
            sigmoid_f := 2039;
        ELSIF x = 11142 THEN
            sigmoid_f := 2039;
        ELSIF x = 11143 THEN
            sigmoid_f := 2039;
        ELSIF x = 11144 THEN
            sigmoid_f := 2039;
        ELSIF x = 11145 THEN
            sigmoid_f := 2039;
        ELSIF x = 11146 THEN
            sigmoid_f := 2039;
        ELSIF x = 11147 THEN
            sigmoid_f := 2039;
        ELSIF x = 11148 THEN
            sigmoid_f := 2039;
        ELSIF x = 11149 THEN
            sigmoid_f := 2039;
        ELSIF x = 11150 THEN
            sigmoid_f := 2039;
        ELSIF x = 11151 THEN
            sigmoid_f := 2039;
        ELSIF x = 11152 THEN
            sigmoid_f := 2039;
        ELSIF x = 11153 THEN
            sigmoid_f := 2039;
        ELSIF x = 11154 THEN
            sigmoid_f := 2039;
        ELSIF x = 11155 THEN
            sigmoid_f := 2039;
        ELSIF x = 11156 THEN
            sigmoid_f := 2039;
        ELSIF x = 11157 THEN
            sigmoid_f := 2039;
        ELSIF x = 11158 THEN
            sigmoid_f := 2039;
        ELSIF x = 11159 THEN
            sigmoid_f := 2039;
        ELSIF x = 11160 THEN
            sigmoid_f := 2039;
        ELSIF x = 11161 THEN
            sigmoid_f := 2039;
        ELSIF x = 11162 THEN
            sigmoid_f := 2039;
        ELSIF x = 11163 THEN
            sigmoid_f := 2039;
        ELSIF x = 11164 THEN
            sigmoid_f := 2039;
        ELSIF x = 11165 THEN
            sigmoid_f := 2039;
        ELSIF x = 11166 THEN
            sigmoid_f := 2039;
        ELSIF x = 11167 THEN
            sigmoid_f := 2039;
        ELSIF x = 11168 THEN
            sigmoid_f := 2039;
        ELSIF x = 11169 THEN
            sigmoid_f := 2039;
        ELSIF x = 11170 THEN
            sigmoid_f := 2039;
        ELSIF x = 11171 THEN
            sigmoid_f := 2039;
        ELSIF x = 11172 THEN
            sigmoid_f := 2039;
        ELSIF x = 11173 THEN
            sigmoid_f := 2039;
        ELSIF x = 11174 THEN
            sigmoid_f := 2039;
        ELSIF x = 11175 THEN
            sigmoid_f := 2039;
        ELSIF x = 11176 THEN
            sigmoid_f := 2039;
        ELSIF x = 11177 THEN
            sigmoid_f := 2039;
        ELSIF x = 11178 THEN
            sigmoid_f := 2039;
        ELSIF x = 11179 THEN
            sigmoid_f := 2039;
        ELSIF x = 11180 THEN
            sigmoid_f := 2039;
        ELSIF x = 11181 THEN
            sigmoid_f := 2039;
        ELSIF x = 11182 THEN
            sigmoid_f := 2039;
        ELSIF x = 11183 THEN
            sigmoid_f := 2039;
        ELSIF x = 11184 THEN
            sigmoid_f := 2039;
        ELSIF x = 11185 THEN
            sigmoid_f := 2039;
        ELSIF x = 11186 THEN
            sigmoid_f := 2039;
        ELSIF x = 11187 THEN
            sigmoid_f := 2039;
        ELSIF x = 11188 THEN
            sigmoid_f := 2039;
        ELSIF x = 11189 THEN
            sigmoid_f := 2039;
        ELSIF x = 11190 THEN
            sigmoid_f := 2039;
        ELSIF x = 11191 THEN
            sigmoid_f := 2039;
        ELSIF x = 11192 THEN
            sigmoid_f := 2039;
        ELSIF x = 11193 THEN
            sigmoid_f := 2039;
        ELSIF x = 11194 THEN
            sigmoid_f := 2039;
        ELSIF x = 11195 THEN
            sigmoid_f := 2039;
        ELSIF x = 11196 THEN
            sigmoid_f := 2039;
        ELSIF x = 11197 THEN
            sigmoid_f := 2039;
        ELSIF x = 11198 THEN
            sigmoid_f := 2039;
        ELSIF x = 11199 THEN
            sigmoid_f := 2039;
        ELSIF x = 11200 THEN
            sigmoid_f := 2039;
        ELSIF x = 11201 THEN
            sigmoid_f := 2039;
        ELSIF x = 11202 THEN
            sigmoid_f := 2039;
        ELSIF x = 11203 THEN
            sigmoid_f := 2039;
        ELSIF x = 11204 THEN
            sigmoid_f := 2039;
        ELSIF x = 11205 THEN
            sigmoid_f := 2039;
        ELSIF x = 11206 THEN
            sigmoid_f := 2039;
        ELSIF x = 11207 THEN
            sigmoid_f := 2039;
        ELSIF x = 11208 THEN
            sigmoid_f := 2039;
        ELSIF x = 11209 THEN
            sigmoid_f := 2039;
        ELSIF x = 11210 THEN
            sigmoid_f := 2039;
        ELSIF x = 11211 THEN
            sigmoid_f := 2039;
        ELSIF x = 11212 THEN
            sigmoid_f := 2039;
        ELSIF x = 11213 THEN
            sigmoid_f := 2039;
        ELSIF x = 11214 THEN
            sigmoid_f := 2039;
        ELSIF x = 11215 THEN
            sigmoid_f := 2039;
        ELSIF x = 11216 THEN
            sigmoid_f := 2039;
        ELSIF x = 11217 THEN
            sigmoid_f := 2039;
        ELSIF x = 11218 THEN
            sigmoid_f := 2039;
        ELSIF x = 11219 THEN
            sigmoid_f := 2039;
        ELSIF x = 11220 THEN
            sigmoid_f := 2039;
        ELSIF x = 11221 THEN
            sigmoid_f := 2039;
        ELSIF x = 11222 THEN
            sigmoid_f := 2039;
        ELSIF x = 11223 THEN
            sigmoid_f := 2039;
        ELSIF x = 11224 THEN
            sigmoid_f := 2039;
        ELSIF x = 11225 THEN
            sigmoid_f := 2039;
        ELSIF x = 11226 THEN
            sigmoid_f := 2039;
        ELSIF x = 11227 THEN
            sigmoid_f := 2039;
        ELSIF x = 11228 THEN
            sigmoid_f := 2039;
        ELSIF x = 11229 THEN
            sigmoid_f := 2039;
        ELSIF x = 11230 THEN
            sigmoid_f := 2039;
        ELSIF x = 11231 THEN
            sigmoid_f := 2039;
        ELSIF x = 11232 THEN
            sigmoid_f := 2039;
        ELSIF x = 11233 THEN
            sigmoid_f := 2039;
        ELSIF x = 11234 THEN
            sigmoid_f := 2039;
        ELSIF x = 11235 THEN
            sigmoid_f := 2039;
        ELSIF x = 11236 THEN
            sigmoid_f := 2039;
        ELSIF x = 11237 THEN
            sigmoid_f := 2039;
        ELSIF x = 11238 THEN
            sigmoid_f := 2039;
        ELSIF x = 11239 THEN
            sigmoid_f := 2039;
        ELSIF x = 11240 THEN
            sigmoid_f := 2039;
        ELSIF x = 11241 THEN
            sigmoid_f := 2039;
        ELSIF x = 11242 THEN
            sigmoid_f := 2039;
        ELSIF x = 11243 THEN
            sigmoid_f := 2039;
        ELSIF x = 11244 THEN
            sigmoid_f := 2039;
        ELSIF x = 11245 THEN
            sigmoid_f := 2039;
        ELSIF x = 11246 THEN
            sigmoid_f := 2039;
        ELSIF x = 11247 THEN
            sigmoid_f := 2039;
        ELSIF x = 11248 THEN
            sigmoid_f := 2039;
        ELSIF x = 11249 THEN
            sigmoid_f := 2039;
        ELSIF x = 11250 THEN
            sigmoid_f := 2039;
        ELSIF x = 11251 THEN
            sigmoid_f := 2039;
        ELSIF x = 11252 THEN
            sigmoid_f := 2039;
        ELSIF x = 11253 THEN
            sigmoid_f := 2039;
        ELSIF x = 11254 THEN
            sigmoid_f := 2039;
        ELSIF x = 11255 THEN
            sigmoid_f := 2039;
        ELSIF x = 11256 THEN
            sigmoid_f := 2039;
        ELSIF x = 11257 THEN
            sigmoid_f := 2039;
        ELSIF x = 11258 THEN
            sigmoid_f := 2039;
        ELSIF x = 11259 THEN
            sigmoid_f := 2039;
        ELSIF x = 11260 THEN
            sigmoid_f := 2039;
        ELSIF x = 11261 THEN
            sigmoid_f := 2039;
        ELSIF x = 11262 THEN
            sigmoid_f := 2039;
        ELSIF x = 11263 THEN
            sigmoid_f := 2039;
        ELSIF x = 11264 THEN
            sigmoid_f := 2039;
        ELSIF x = 11265 THEN
            sigmoid_f := 2039;
        ELSIF x = 11266 THEN
            sigmoid_f := 2039;
        ELSIF x = 11267 THEN
            sigmoid_f := 2039;
        ELSIF x = 11268 THEN
            sigmoid_f := 2039;
        ELSIF x = 11269 THEN
            sigmoid_f := 2039;
        ELSIF x = 11270 THEN
            sigmoid_f := 2039;
        ELSIF x = 11271 THEN
            sigmoid_f := 2039;
        ELSIF x = 11272 THEN
            sigmoid_f := 2039;
        ELSIF x = 11273 THEN
            sigmoid_f := 2039;
        ELSIF x = 11274 THEN
            sigmoid_f := 2039;
        ELSIF x = 11275 THEN
            sigmoid_f := 2039;
        ELSIF x = 11276 THEN
            sigmoid_f := 2039;
        ELSIF x = 11277 THEN
            sigmoid_f := 2039;
        ELSIF x = 11278 THEN
            sigmoid_f := 2039;
        ELSIF x = 11279 THEN
            sigmoid_f := 2039;
        ELSIF x = 11280 THEN
            sigmoid_f := 2039;
        ELSIF x = 11281 THEN
            sigmoid_f := 2039;
        ELSIF x = 11282 THEN
            sigmoid_f := 2039;
        ELSIF x = 11283 THEN
            sigmoid_f := 2039;
        ELSIF x = 11284 THEN
            sigmoid_f := 2039;
        ELSIF x = 11285 THEN
            sigmoid_f := 2039;
        ELSIF x = 11286 THEN
            sigmoid_f := 2039;
        ELSIF x = 11287 THEN
            sigmoid_f := 2039;
        ELSIF x = 11288 THEN
            sigmoid_f := 2039;
        ELSIF x = 11289 THEN
            sigmoid_f := 2039;
        ELSIF x = 11290 THEN
            sigmoid_f := 2039;
        ELSIF x = 11291 THEN
            sigmoid_f := 2039;
        ELSIF x = 11292 THEN
            sigmoid_f := 2039;
        ELSIF x = 11293 THEN
            sigmoid_f := 2039;
        ELSIF x = 11294 THEN
            sigmoid_f := 2039;
        ELSIF x = 11295 THEN
            sigmoid_f := 2039;
        ELSIF x = 11296 THEN
            sigmoid_f := 2039;
        ELSIF x = 11297 THEN
            sigmoid_f := 2039;
        ELSIF x = 11298 THEN
            sigmoid_f := 2039;
        ELSIF x = 11299 THEN
            sigmoid_f := 2039;
        ELSIF x = 11300 THEN
            sigmoid_f := 2039;
        ELSIF x = 11301 THEN
            sigmoid_f := 2039;
        ELSIF x = 11302 THEN
            sigmoid_f := 2039;
        ELSIF x = 11303 THEN
            sigmoid_f := 2039;
        ELSIF x = 11304 THEN
            sigmoid_f := 2039;
        ELSIF x = 11305 THEN
            sigmoid_f := 2039;
        ELSIF x = 11306 THEN
            sigmoid_f := 2039;
        ELSIF x = 11307 THEN
            sigmoid_f := 2039;
        ELSIF x = 11308 THEN
            sigmoid_f := 2039;
        ELSIF x = 11309 THEN
            sigmoid_f := 2039;
        ELSIF x = 11310 THEN
            sigmoid_f := 2039;
        ELSIF x = 11311 THEN
            sigmoid_f := 2039;
        ELSIF x = 11312 THEN
            sigmoid_f := 2039;
        ELSIF x = 11313 THEN
            sigmoid_f := 2039;
        ELSIF x = 11314 THEN
            sigmoid_f := 2039;
        ELSIF x = 11315 THEN
            sigmoid_f := 2039;
        ELSIF x = 11316 THEN
            sigmoid_f := 2039;
        ELSIF x = 11317 THEN
            sigmoid_f := 2039;
        ELSIF x = 11318 THEN
            sigmoid_f := 2039;
        ELSIF x = 11319 THEN
            sigmoid_f := 2039;
        ELSIF x = 11320 THEN
            sigmoid_f := 2039;
        ELSIF x = 11321 THEN
            sigmoid_f := 2039;
        ELSIF x = 11322 THEN
            sigmoid_f := 2039;
        ELSIF x = 11323 THEN
            sigmoid_f := 2039;
        ELSIF x = 11324 THEN
            sigmoid_f := 2039;
        ELSIF x = 11325 THEN
            sigmoid_f := 2039;
        ELSIF x = 11326 THEN
            sigmoid_f := 2039;
        ELSIF x = 11327 THEN
            sigmoid_f := 2039;
        ELSIF x = 11328 THEN
            sigmoid_f := 2039;
        ELSIF x = 11329 THEN
            sigmoid_f := 2039;
        ELSIF x = 11330 THEN
            sigmoid_f := 2039;
        ELSIF x = 11331 THEN
            sigmoid_f := 2039;
        ELSIF x = 11332 THEN
            sigmoid_f := 2039;
        ELSIF x = 11333 THEN
            sigmoid_f := 2039;
        ELSIF x = 11334 THEN
            sigmoid_f := 2039;
        ELSIF x = 11335 THEN
            sigmoid_f := 2039;
        ELSIF x = 11336 THEN
            sigmoid_f := 2039;
        ELSIF x = 11337 THEN
            sigmoid_f := 2039;
        ELSIF x = 11338 THEN
            sigmoid_f := 2039;
        ELSIF x = 11339 THEN
            sigmoid_f := 2039;
        ELSIF x = 11340 THEN
            sigmoid_f := 2039;
        ELSIF x = 11341 THEN
            sigmoid_f := 2039;
        ELSIF x = 11342 THEN
            sigmoid_f := 2039;
        ELSIF x = 11343 THEN
            sigmoid_f := 2039;
        ELSIF x = 11344 THEN
            sigmoid_f := 2039;
        ELSIF x = 11345 THEN
            sigmoid_f := 2039;
        ELSIF x = 11346 THEN
            sigmoid_f := 2039;
        ELSIF x = 11347 THEN
            sigmoid_f := 2039;
        ELSIF x = 11348 THEN
            sigmoid_f := 2039;
        ELSIF x = 11349 THEN
            sigmoid_f := 2039;
        ELSIF x = 11350 THEN
            sigmoid_f := 2039;
        ELSIF x = 11351 THEN
            sigmoid_f := 2039;
        ELSIF x = 11352 THEN
            sigmoid_f := 2039;
        ELSIF x = 11353 THEN
            sigmoid_f := 2039;
        ELSIF x = 11354 THEN
            sigmoid_f := 2039;
        ELSIF x = 11355 THEN
            sigmoid_f := 2039;
        ELSIF x = 11356 THEN
            sigmoid_f := 2039;
        ELSIF x = 11357 THEN
            sigmoid_f := 2039;
        ELSIF x = 11358 THEN
            sigmoid_f := 2039;
        ELSIF x = 11359 THEN
            sigmoid_f := 2039;
        ELSIF x = 11360 THEN
            sigmoid_f := 2039;
        ELSIF x = 11361 THEN
            sigmoid_f := 2039;
        ELSIF x = 11362 THEN
            sigmoid_f := 2039;
        ELSIF x = 11363 THEN
            sigmoid_f := 2039;
        ELSIF x = 11364 THEN
            sigmoid_f := 2039;
        ELSIF x = 11365 THEN
            sigmoid_f := 2039;
        ELSIF x = 11366 THEN
            sigmoid_f := 2039;
        ELSIF x = 11367 THEN
            sigmoid_f := 2039;
        ELSIF x = 11368 THEN
            sigmoid_f := 2039;
        ELSIF x = 11369 THEN
            sigmoid_f := 2039;
        ELSIF x = 11370 THEN
            sigmoid_f := 2039;
        ELSIF x = 11371 THEN
            sigmoid_f := 2039;
        ELSIF x = 11372 THEN
            sigmoid_f := 2039;
        ELSIF x = 11373 THEN
            sigmoid_f := 2039;
        ELSIF x = 11374 THEN
            sigmoid_f := 2039;
        ELSIF x = 11375 THEN
            sigmoid_f := 2039;
        ELSIF x = 11376 THEN
            sigmoid_f := 2039;
        ELSIF x = 11377 THEN
            sigmoid_f := 2039;
        ELSIF x = 11378 THEN
            sigmoid_f := 2040;
        ELSIF x = 11379 THEN
            sigmoid_f := 2040;
        ELSIF x = 11380 THEN
            sigmoid_f := 2040;
        ELSIF x = 11381 THEN
            sigmoid_f := 2040;
        ELSIF x = 11382 THEN
            sigmoid_f := 2040;
        ELSIF x = 11383 THEN
            sigmoid_f := 2040;
        ELSIF x = 11384 THEN
            sigmoid_f := 2040;
        ELSIF x = 11385 THEN
            sigmoid_f := 2040;
        ELSIF x = 11386 THEN
            sigmoid_f := 2040;
        ELSIF x = 11387 THEN
            sigmoid_f := 2040;
        ELSIF x = 11388 THEN
            sigmoid_f := 2040;
        ELSIF x = 11389 THEN
            sigmoid_f := 2040;
        ELSIF x = 11390 THEN
            sigmoid_f := 2040;
        ELSIF x = 11391 THEN
            sigmoid_f := 2040;
        ELSIF x = 11392 THEN
            sigmoid_f := 2040;
        ELSIF x = 11393 THEN
            sigmoid_f := 2040;
        ELSIF x = 11394 THEN
            sigmoid_f := 2040;
        ELSIF x = 11395 THEN
            sigmoid_f := 2040;
        ELSIF x = 11396 THEN
            sigmoid_f := 2040;
        ELSIF x = 11397 THEN
            sigmoid_f := 2040;
        ELSIF x = 11398 THEN
            sigmoid_f := 2040;
        ELSIF x = 11399 THEN
            sigmoid_f := 2040;
        ELSIF x = 11400 THEN
            sigmoid_f := 2040;
        ELSIF x = 11401 THEN
            sigmoid_f := 2040;
        ELSIF x = 11402 THEN
            sigmoid_f := 2040;
        ELSIF x = 11403 THEN
            sigmoid_f := 2040;
        ELSIF x = 11404 THEN
            sigmoid_f := 2040;
        ELSIF x = 11405 THEN
            sigmoid_f := 2040;
        ELSIF x = 11406 THEN
            sigmoid_f := 2040;
        ELSIF x = 11407 THEN
            sigmoid_f := 2040;
        ELSIF x = 11408 THEN
            sigmoid_f := 2040;
        ELSIF x = 11409 THEN
            sigmoid_f := 2040;
        ELSIF x = 11410 THEN
            sigmoid_f := 2040;
        ELSIF x = 11411 THEN
            sigmoid_f := 2040;
        ELSIF x = 11412 THEN
            sigmoid_f := 2040;
        ELSIF x = 11413 THEN
            sigmoid_f := 2040;
        ELSIF x = 11414 THEN
            sigmoid_f := 2040;
        ELSIF x = 11415 THEN
            sigmoid_f := 2040;
        ELSIF x = 11416 THEN
            sigmoid_f := 2040;
        ELSIF x = 11417 THEN
            sigmoid_f := 2040;
        ELSIF x = 11418 THEN
            sigmoid_f := 2040;
        ELSIF x = 11419 THEN
            sigmoid_f := 2040;
        ELSIF x = 11420 THEN
            sigmoid_f := 2040;
        ELSIF x = 11421 THEN
            sigmoid_f := 2040;
        ELSIF x = 11422 THEN
            sigmoid_f := 2040;
        ELSIF x = 11423 THEN
            sigmoid_f := 2040;
        ELSIF x = 11424 THEN
            sigmoid_f := 2040;
        ELSIF x = 11425 THEN
            sigmoid_f := 2040;
        ELSIF x = 11426 THEN
            sigmoid_f := 2040;
        ELSIF x = 11427 THEN
            sigmoid_f := 2040;
        ELSIF x = 11428 THEN
            sigmoid_f := 2040;
        ELSIF x = 11429 THEN
            sigmoid_f := 2040;
        ELSIF x = 11430 THEN
            sigmoid_f := 2040;
        ELSIF x = 11431 THEN
            sigmoid_f := 2040;
        ELSIF x = 11432 THEN
            sigmoid_f := 2040;
        ELSIF x = 11433 THEN
            sigmoid_f := 2040;
        ELSIF x = 11434 THEN
            sigmoid_f := 2040;
        ELSIF x = 11435 THEN
            sigmoid_f := 2040;
        ELSIF x = 11436 THEN
            sigmoid_f := 2040;
        ELSIF x = 11437 THEN
            sigmoid_f := 2040;
        ELSIF x = 11438 THEN
            sigmoid_f := 2040;
        ELSIF x = 11439 THEN
            sigmoid_f := 2040;
        ELSIF x = 11440 THEN
            sigmoid_f := 2040;
        ELSIF x = 11441 THEN
            sigmoid_f := 2040;
        ELSIF x = 11442 THEN
            sigmoid_f := 2040;
        ELSIF x = 11443 THEN
            sigmoid_f := 2040;
        ELSIF x = 11444 THEN
            sigmoid_f := 2040;
        ELSIF x = 11445 THEN
            sigmoid_f := 2040;
        ELSIF x = 11446 THEN
            sigmoid_f := 2040;
        ELSIF x = 11447 THEN
            sigmoid_f := 2040;
        ELSIF x = 11448 THEN
            sigmoid_f := 2040;
        ELSIF x = 11449 THEN
            sigmoid_f := 2040;
        ELSIF x = 11450 THEN
            sigmoid_f := 2040;
        ELSIF x = 11451 THEN
            sigmoid_f := 2040;
        ELSIF x = 11452 THEN
            sigmoid_f := 2040;
        ELSIF x = 11453 THEN
            sigmoid_f := 2040;
        ELSIF x = 11454 THEN
            sigmoid_f := 2040;
        ELSIF x = 11455 THEN
            sigmoid_f := 2040;
        ELSIF x = 11456 THEN
            sigmoid_f := 2040;
        ELSIF x = 11457 THEN
            sigmoid_f := 2040;
        ELSIF x = 11458 THEN
            sigmoid_f := 2040;
        ELSIF x = 11459 THEN
            sigmoid_f := 2040;
        ELSIF x = 11460 THEN
            sigmoid_f := 2040;
        ELSIF x = 11461 THEN
            sigmoid_f := 2040;
        ELSIF x = 11462 THEN
            sigmoid_f := 2040;
        ELSIF x = 11463 THEN
            sigmoid_f := 2040;
        ELSIF x = 11464 THEN
            sigmoid_f := 2040;
        ELSIF x = 11465 THEN
            sigmoid_f := 2040;
        ELSIF x = 11466 THEN
            sigmoid_f := 2040;
        ELSIF x = 11467 THEN
            sigmoid_f := 2040;
        ELSIF x = 11468 THEN
            sigmoid_f := 2040;
        ELSIF x = 11469 THEN
            sigmoid_f := 2040;
        ELSIF x = 11470 THEN
            sigmoid_f := 2040;
        ELSIF x = 11471 THEN
            sigmoid_f := 2040;
        ELSIF x = 11472 THEN
            sigmoid_f := 2040;
        ELSIF x = 11473 THEN
            sigmoid_f := 2040;
        ELSIF x = 11474 THEN
            sigmoid_f := 2040;
        ELSIF x = 11475 THEN
            sigmoid_f := 2040;
        ELSIF x = 11476 THEN
            sigmoid_f := 2040;
        ELSIF x = 11477 THEN
            sigmoid_f := 2040;
        ELSIF x = 11478 THEN
            sigmoid_f := 2040;
        ELSIF x = 11479 THEN
            sigmoid_f := 2040;
        ELSIF x = 11480 THEN
            sigmoid_f := 2040;
        ELSIF x = 11481 THEN
            sigmoid_f := 2040;
        ELSIF x = 11482 THEN
            sigmoid_f := 2040;
        ELSIF x = 11483 THEN
            sigmoid_f := 2040;
        ELSIF x = 11484 THEN
            sigmoid_f := 2040;
        ELSIF x = 11485 THEN
            sigmoid_f := 2040;
        ELSIF x = 11486 THEN
            sigmoid_f := 2040;
        ELSIF x = 11487 THEN
            sigmoid_f := 2040;
        ELSIF x = 11488 THEN
            sigmoid_f := 2040;
        ELSIF x = 11489 THEN
            sigmoid_f := 2040;
        ELSIF x = 11490 THEN
            sigmoid_f := 2040;
        ELSIF x = 11491 THEN
            sigmoid_f := 2040;
        ELSIF x = 11492 THEN
            sigmoid_f := 2040;
        ELSIF x = 11493 THEN
            sigmoid_f := 2040;
        ELSIF x = 11494 THEN
            sigmoid_f := 2040;
        ELSIF x = 11495 THEN
            sigmoid_f := 2040;
        ELSIF x = 11496 THEN
            sigmoid_f := 2040;
        ELSIF x = 11497 THEN
            sigmoid_f := 2040;
        ELSIF x = 11498 THEN
            sigmoid_f := 2040;
        ELSIF x = 11499 THEN
            sigmoid_f := 2040;
        ELSIF x = 11500 THEN
            sigmoid_f := 2040;
        ELSIF x = 11501 THEN
            sigmoid_f := 2040;
        ELSIF x = 11502 THEN
            sigmoid_f := 2040;
        ELSIF x = 11503 THEN
            sigmoid_f := 2040;
        ELSIF x = 11504 THEN
            sigmoid_f := 2040;
        ELSIF x = 11505 THEN
            sigmoid_f := 2040;
        ELSIF x = 11506 THEN
            sigmoid_f := 2040;
        ELSIF x = 11507 THEN
            sigmoid_f := 2040;
        ELSIF x = 11508 THEN
            sigmoid_f := 2040;
        ELSIF x = 11509 THEN
            sigmoid_f := 2040;
        ELSIF x = 11510 THEN
            sigmoid_f := 2040;
        ELSIF x = 11511 THEN
            sigmoid_f := 2040;
        ELSIF x = 11512 THEN
            sigmoid_f := 2040;
        ELSIF x = 11513 THEN
            sigmoid_f := 2040;
        ELSIF x = 11514 THEN
            sigmoid_f := 2040;
        ELSIF x = 11515 THEN
            sigmoid_f := 2040;
        ELSIF x = 11516 THEN
            sigmoid_f := 2040;
        ELSIF x = 11517 THEN
            sigmoid_f := 2040;
        ELSIF x = 11518 THEN
            sigmoid_f := 2040;
        ELSIF x = 11519 THEN
            sigmoid_f := 2040;
        ELSIF x = 11520 THEN
            sigmoid_f := 2040;
        ELSIF x = 11521 THEN
            sigmoid_f := 2040;
        ELSIF x = 11522 THEN
            sigmoid_f := 2040;
        ELSIF x = 11523 THEN
            sigmoid_f := 2040;
        ELSIF x = 11524 THEN
            sigmoid_f := 2040;
        ELSIF x = 11525 THEN
            sigmoid_f := 2040;
        ELSIF x = 11526 THEN
            sigmoid_f := 2040;
        ELSIF x = 11527 THEN
            sigmoid_f := 2040;
        ELSIF x = 11528 THEN
            sigmoid_f := 2040;
        ELSIF x = 11529 THEN
            sigmoid_f := 2040;
        ELSIF x = 11530 THEN
            sigmoid_f := 2040;
        ELSIF x = 11531 THEN
            sigmoid_f := 2040;
        ELSIF x = 11532 THEN
            sigmoid_f := 2040;
        ELSIF x = 11533 THEN
            sigmoid_f := 2040;
        ELSIF x = 11534 THEN
            sigmoid_f := 2040;
        ELSIF x = 11535 THEN
            sigmoid_f := 2040;
        ELSIF x = 11536 THEN
            sigmoid_f := 2040;
        ELSIF x = 11537 THEN
            sigmoid_f := 2040;
        ELSIF x = 11538 THEN
            sigmoid_f := 2040;
        ELSIF x = 11539 THEN
            sigmoid_f := 2040;
        ELSIF x = 11540 THEN
            sigmoid_f := 2040;
        ELSIF x = 11541 THEN
            sigmoid_f := 2040;
        ELSIF x = 11542 THEN
            sigmoid_f := 2040;
        ELSIF x = 11543 THEN
            sigmoid_f := 2040;
        ELSIF x = 11544 THEN
            sigmoid_f := 2040;
        ELSIF x = 11545 THEN
            sigmoid_f := 2040;
        ELSIF x = 11546 THEN
            sigmoid_f := 2040;
        ELSIF x = 11547 THEN
            sigmoid_f := 2040;
        ELSIF x = 11548 THEN
            sigmoid_f := 2040;
        ELSIF x = 11549 THEN
            sigmoid_f := 2040;
        ELSIF x = 11550 THEN
            sigmoid_f := 2040;
        ELSIF x = 11551 THEN
            sigmoid_f := 2040;
        ELSIF x = 11552 THEN
            sigmoid_f := 2040;
        ELSIF x = 11553 THEN
            sigmoid_f := 2040;
        ELSIF x = 11554 THEN
            sigmoid_f := 2040;
        ELSIF x = 11555 THEN
            sigmoid_f := 2040;
        ELSIF x = 11556 THEN
            sigmoid_f := 2040;
        ELSIF x = 11557 THEN
            sigmoid_f := 2040;
        ELSIF x = 11558 THEN
            sigmoid_f := 2040;
        ELSIF x = 11559 THEN
            sigmoid_f := 2040;
        ELSIF x = 11560 THEN
            sigmoid_f := 2040;
        ELSIF x = 11561 THEN
            sigmoid_f := 2040;
        ELSIF x = 11562 THEN
            sigmoid_f := 2040;
        ELSIF x = 11563 THEN
            sigmoid_f := 2040;
        ELSIF x = 11564 THEN
            sigmoid_f := 2040;
        ELSIF x = 11565 THEN
            sigmoid_f := 2040;
        ELSIF x = 11566 THEN
            sigmoid_f := 2040;
        ELSIF x = 11567 THEN
            sigmoid_f := 2040;
        ELSIF x = 11568 THEN
            sigmoid_f := 2040;
        ELSIF x = 11569 THEN
            sigmoid_f := 2040;
        ELSIF x = 11570 THEN
            sigmoid_f := 2040;
        ELSIF x = 11571 THEN
            sigmoid_f := 2040;
        ELSIF x = 11572 THEN
            sigmoid_f := 2040;
        ELSIF x = 11573 THEN
            sigmoid_f := 2040;
        ELSIF x = 11574 THEN
            sigmoid_f := 2040;
        ELSIF x = 11575 THEN
            sigmoid_f := 2040;
        ELSIF x = 11576 THEN
            sigmoid_f := 2040;
        ELSIF x = 11577 THEN
            sigmoid_f := 2040;
        ELSIF x = 11578 THEN
            sigmoid_f := 2040;
        ELSIF x = 11579 THEN
            sigmoid_f := 2040;
        ELSIF x = 11580 THEN
            sigmoid_f := 2040;
        ELSIF x = 11581 THEN
            sigmoid_f := 2040;
        ELSIF x = 11582 THEN
            sigmoid_f := 2040;
        ELSIF x = 11583 THEN
            sigmoid_f := 2040;
        ELSIF x = 11584 THEN
            sigmoid_f := 2040;
        ELSIF x = 11585 THEN
            sigmoid_f := 2040;
        ELSIF x = 11586 THEN
            sigmoid_f := 2040;
        ELSIF x = 11587 THEN
            sigmoid_f := 2040;
        ELSIF x = 11588 THEN
            sigmoid_f := 2040;
        ELSIF x = 11589 THEN
            sigmoid_f := 2040;
        ELSIF x = 11590 THEN
            sigmoid_f := 2040;
        ELSIF x = 11591 THEN
            sigmoid_f := 2040;
        ELSIF x = 11592 THEN
            sigmoid_f := 2040;
        ELSIF x = 11593 THEN
            sigmoid_f := 2040;
        ELSIF x = 11594 THEN
            sigmoid_f := 2040;
        ELSIF x = 11595 THEN
            sigmoid_f := 2040;
        ELSIF x = 11596 THEN
            sigmoid_f := 2040;
        ELSIF x = 11597 THEN
            sigmoid_f := 2040;
        ELSIF x = 11598 THEN
            sigmoid_f := 2040;
        ELSIF x = 11599 THEN
            sigmoid_f := 2040;
        ELSIF x = 11600 THEN
            sigmoid_f := 2040;
        ELSIF x = 11601 THEN
            sigmoid_f := 2040;
        ELSIF x = 11602 THEN
            sigmoid_f := 2040;
        ELSIF x = 11603 THEN
            sigmoid_f := 2040;
        ELSIF x = 11604 THEN
            sigmoid_f := 2040;
        ELSIF x = 11605 THEN
            sigmoid_f := 2040;
        ELSIF x = 11606 THEN
            sigmoid_f := 2041;
        ELSIF x = 11607 THEN
            sigmoid_f := 2041;
        ELSIF x = 11608 THEN
            sigmoid_f := 2041;
        ELSIF x = 11609 THEN
            sigmoid_f := 2041;
        ELSIF x = 11610 THEN
            sigmoid_f := 2041;
        ELSIF x = 11611 THEN
            sigmoid_f := 2041;
        ELSIF x = 11612 THEN
            sigmoid_f := 2041;
        ELSIF x = 11613 THEN
            sigmoid_f := 2041;
        ELSIF x = 11614 THEN
            sigmoid_f := 2041;
        ELSIF x = 11615 THEN
            sigmoid_f := 2041;
        ELSIF x = 11616 THEN
            sigmoid_f := 2041;
        ELSIF x = 11617 THEN
            sigmoid_f := 2041;
        ELSIF x = 11618 THEN
            sigmoid_f := 2041;
        ELSIF x = 11619 THEN
            sigmoid_f := 2041;
        ELSIF x = 11620 THEN
            sigmoid_f := 2041;
        ELSIF x = 11621 THEN
            sigmoid_f := 2041;
        ELSIF x = 11622 THEN
            sigmoid_f := 2041;
        ELSIF x = 11623 THEN
            sigmoid_f := 2041;
        ELSIF x = 11624 THEN
            sigmoid_f := 2041;
        ELSIF x = 11625 THEN
            sigmoid_f := 2041;
        ELSIF x = 11626 THEN
            sigmoid_f := 2041;
        ELSIF x = 11627 THEN
            sigmoid_f := 2041;
        ELSIF x = 11628 THEN
            sigmoid_f := 2041;
        ELSIF x = 11629 THEN
            sigmoid_f := 2041;
        ELSIF x = 11630 THEN
            sigmoid_f := 2041;
        ELSIF x = 11631 THEN
            sigmoid_f := 2041;
        ELSIF x = 11632 THEN
            sigmoid_f := 2041;
        ELSIF x = 11633 THEN
            sigmoid_f := 2041;
        ELSIF x = 11634 THEN
            sigmoid_f := 2041;
        ELSIF x = 11635 THEN
            sigmoid_f := 2041;
        ELSIF x = 11636 THEN
            sigmoid_f := 2041;
        ELSIF x = 11637 THEN
            sigmoid_f := 2041;
        ELSIF x = 11638 THEN
            sigmoid_f := 2041;
        ELSIF x = 11639 THEN
            sigmoid_f := 2041;
        ELSIF x = 11640 THEN
            sigmoid_f := 2041;
        ELSIF x = 11641 THEN
            sigmoid_f := 2041;
        ELSIF x = 11642 THEN
            sigmoid_f := 2041;
        ELSIF x = 11643 THEN
            sigmoid_f := 2041;
        ELSIF x = 11644 THEN
            sigmoid_f := 2041;
        ELSIF x = 11645 THEN
            sigmoid_f := 2041;
        ELSIF x = 11646 THEN
            sigmoid_f := 2041;
        ELSIF x = 11647 THEN
            sigmoid_f := 2041;
        ELSIF x = 11648 THEN
            sigmoid_f := 2041;
        ELSIF x = 11649 THEN
            sigmoid_f := 2041;
        ELSIF x = 11650 THEN
            sigmoid_f := 2041;
        ELSIF x = 11651 THEN
            sigmoid_f := 2041;
        ELSIF x = 11652 THEN
            sigmoid_f := 2041;
        ELSIF x = 11653 THEN
            sigmoid_f := 2041;
        ELSIF x = 11654 THEN
            sigmoid_f := 2041;
        ELSIF x = 11655 THEN
            sigmoid_f := 2041;
        ELSIF x = 11656 THEN
            sigmoid_f := 2041;
        ELSIF x = 11657 THEN
            sigmoid_f := 2041;
        ELSIF x = 11658 THEN
            sigmoid_f := 2041;
        ELSIF x = 11659 THEN
            sigmoid_f := 2041;
        ELSIF x = 11660 THEN
            sigmoid_f := 2041;
        ELSIF x = 11661 THEN
            sigmoid_f := 2041;
        ELSIF x = 11662 THEN
            sigmoid_f := 2041;
        ELSIF x = 11663 THEN
            sigmoid_f := 2041;
        ELSIF x = 11664 THEN
            sigmoid_f := 2041;
        ELSIF x = 11665 THEN
            sigmoid_f := 2041;
        ELSIF x = 11666 THEN
            sigmoid_f := 2041;
        ELSIF x = 11667 THEN
            sigmoid_f := 2041;
        ELSIF x = 11668 THEN
            sigmoid_f := 2041;
        ELSIF x = 11669 THEN
            sigmoid_f := 2041;
        ELSIF x = 11670 THEN
            sigmoid_f := 2041;
        ELSIF x = 11671 THEN
            sigmoid_f := 2041;
        ELSIF x = 11672 THEN
            sigmoid_f := 2041;
        ELSIF x = 11673 THEN
            sigmoid_f := 2041;
        ELSIF x = 11674 THEN
            sigmoid_f := 2041;
        ELSIF x = 11675 THEN
            sigmoid_f := 2041;
        ELSIF x = 11676 THEN
            sigmoid_f := 2041;
        ELSIF x = 11677 THEN
            sigmoid_f := 2041;
        ELSIF x = 11678 THEN
            sigmoid_f := 2041;
        ELSIF x = 11679 THEN
            sigmoid_f := 2041;
        ELSIF x = 11680 THEN
            sigmoid_f := 2041;
        ELSIF x = 11681 THEN
            sigmoid_f := 2041;
        ELSIF x = 11682 THEN
            sigmoid_f := 2041;
        ELSIF x = 11683 THEN
            sigmoid_f := 2041;
        ELSIF x = 11684 THEN
            sigmoid_f := 2041;
        ELSIF x = 11685 THEN
            sigmoid_f := 2041;
        ELSIF x = 11686 THEN
            sigmoid_f := 2041;
        ELSIF x = 11687 THEN
            sigmoid_f := 2041;
        ELSIF x = 11688 THEN
            sigmoid_f := 2041;
        ELSIF x = 11689 THEN
            sigmoid_f := 2041;
        ELSIF x = 11690 THEN
            sigmoid_f := 2041;
        ELSIF x = 11691 THEN
            sigmoid_f := 2041;
        ELSIF x = 11692 THEN
            sigmoid_f := 2041;
        ELSIF x = 11693 THEN
            sigmoid_f := 2041;
        ELSIF x = 11694 THEN
            sigmoid_f := 2041;
        ELSIF x = 11695 THEN
            sigmoid_f := 2041;
        ELSIF x = 11696 THEN
            sigmoid_f := 2041;
        ELSIF x = 11697 THEN
            sigmoid_f := 2041;
        ELSIF x = 11698 THEN
            sigmoid_f := 2041;
        ELSIF x = 11699 THEN
            sigmoid_f := 2041;
        ELSIF x = 11700 THEN
            sigmoid_f := 2041;
        ELSIF x = 11701 THEN
            sigmoid_f := 2041;
        ELSIF x = 11702 THEN
            sigmoid_f := 2041;
        ELSIF x = 11703 THEN
            sigmoid_f := 2041;
        ELSIF x = 11704 THEN
            sigmoid_f := 2041;
        ELSIF x = 11705 THEN
            sigmoid_f := 2041;
        ELSIF x = 11706 THEN
            sigmoid_f := 2041;
        ELSIF x = 11707 THEN
            sigmoid_f := 2041;
        ELSIF x = 11708 THEN
            sigmoid_f := 2041;
        ELSIF x = 11709 THEN
            sigmoid_f := 2041;
        ELSIF x = 11710 THEN
            sigmoid_f := 2041;
        ELSIF x = 11711 THEN
            sigmoid_f := 2041;
        ELSIF x = 11712 THEN
            sigmoid_f := 2041;
        ELSIF x = 11713 THEN
            sigmoid_f := 2041;
        ELSIF x = 11714 THEN
            sigmoid_f := 2041;
        ELSIF x = 11715 THEN
            sigmoid_f := 2041;
        ELSIF x = 11716 THEN
            sigmoid_f := 2041;
        ELSIF x = 11717 THEN
            sigmoid_f := 2041;
        ELSIF x = 11718 THEN
            sigmoid_f := 2041;
        ELSIF x = 11719 THEN
            sigmoid_f := 2041;
        ELSIF x = 11720 THEN
            sigmoid_f := 2041;
        ELSIF x = 11721 THEN
            sigmoid_f := 2041;
        ELSIF x = 11722 THEN
            sigmoid_f := 2041;
        ELSIF x = 11723 THEN
            sigmoid_f := 2041;
        ELSIF x = 11724 THEN
            sigmoid_f := 2041;
        ELSIF x = 11725 THEN
            sigmoid_f := 2041;
        ELSIF x = 11726 THEN
            sigmoid_f := 2041;
        ELSIF x = 11727 THEN
            sigmoid_f := 2041;
        ELSIF x = 11728 THEN
            sigmoid_f := 2041;
        ELSIF x = 11729 THEN
            sigmoid_f := 2041;
        ELSIF x = 11730 THEN
            sigmoid_f := 2041;
        ELSIF x = 11731 THEN
            sigmoid_f := 2041;
        ELSIF x = 11732 THEN
            sigmoid_f := 2041;
        ELSIF x = 11733 THEN
            sigmoid_f := 2041;
        ELSIF x = 11734 THEN
            sigmoid_f := 2041;
        ELSIF x = 11735 THEN
            sigmoid_f := 2041;
        ELSIF x = 11736 THEN
            sigmoid_f := 2041;
        ELSIF x = 11737 THEN
            sigmoid_f := 2041;
        ELSIF x = 11738 THEN
            sigmoid_f := 2041;
        ELSIF x = 11739 THEN
            sigmoid_f := 2041;
        ELSIF x = 11740 THEN
            sigmoid_f := 2041;
        ELSIF x = 11741 THEN
            sigmoid_f := 2041;
        ELSIF x = 11742 THEN
            sigmoid_f := 2041;
        ELSIF x = 11743 THEN
            sigmoid_f := 2041;
        ELSIF x = 11744 THEN
            sigmoid_f := 2041;
        ELSIF x = 11745 THEN
            sigmoid_f := 2041;
        ELSIF x = 11746 THEN
            sigmoid_f := 2041;
        ELSIF x = 11747 THEN
            sigmoid_f := 2041;
        ELSIF x = 11748 THEN
            sigmoid_f := 2041;
        ELSIF x = 11749 THEN
            sigmoid_f := 2041;
        ELSIF x = 11750 THEN
            sigmoid_f := 2041;
        ELSIF x = 11751 THEN
            sigmoid_f := 2041;
        ELSIF x = 11752 THEN
            sigmoid_f := 2041;
        ELSIF x = 11753 THEN
            sigmoid_f := 2041;
        ELSIF x = 11754 THEN
            sigmoid_f := 2041;
        ELSIF x = 11755 THEN
            sigmoid_f := 2041;
        ELSIF x = 11756 THEN
            sigmoid_f := 2041;
        ELSIF x = 11757 THEN
            sigmoid_f := 2041;
        ELSIF x = 11758 THEN
            sigmoid_f := 2041;
        ELSIF x = 11759 THEN
            sigmoid_f := 2041;
        ELSIF x = 11760 THEN
            sigmoid_f := 2041;
        ELSIF x = 11761 THEN
            sigmoid_f := 2041;
        ELSIF x = 11762 THEN
            sigmoid_f := 2041;
        ELSIF x = 11763 THEN
            sigmoid_f := 2041;
        ELSIF x = 11764 THEN
            sigmoid_f := 2041;
        ELSIF x = 11765 THEN
            sigmoid_f := 2041;
        ELSIF x = 11766 THEN
            sigmoid_f := 2041;
        ELSIF x = 11767 THEN
            sigmoid_f := 2041;
        ELSIF x = 11768 THEN
            sigmoid_f := 2041;
        ELSIF x = 11769 THEN
            sigmoid_f := 2041;
        ELSIF x = 11770 THEN
            sigmoid_f := 2041;
        ELSIF x = 11771 THEN
            sigmoid_f := 2041;
        ELSIF x = 11772 THEN
            sigmoid_f := 2041;
        ELSIF x = 11773 THEN
            sigmoid_f := 2041;
        ELSIF x = 11774 THEN
            sigmoid_f := 2041;
        ELSIF x = 11775 THEN
            sigmoid_f := 2041;
        ELSIF x = 11776 THEN
            sigmoid_f := 2042;
        ELSIF x = 11777 THEN
            sigmoid_f := 2042;
        ELSIF x = 11778 THEN
            sigmoid_f := 2042;
        ELSIF x = 11779 THEN
            sigmoid_f := 2042;
        ELSIF x = 11780 THEN
            sigmoid_f := 2042;
        ELSIF x = 11781 THEN
            sigmoid_f := 2042;
        ELSIF x = 11782 THEN
            sigmoid_f := 2042;
        ELSIF x = 11783 THEN
            sigmoid_f := 2042;
        ELSIF x = 11784 THEN
            sigmoid_f := 2042;
        ELSIF x = 11785 THEN
            sigmoid_f := 2042;
        ELSIF x = 11786 THEN
            sigmoid_f := 2042;
        ELSIF x = 11787 THEN
            sigmoid_f := 2042;
        ELSIF x = 11788 THEN
            sigmoid_f := 2042;
        ELSIF x = 11789 THEN
            sigmoid_f := 2042;
        ELSIF x = 11790 THEN
            sigmoid_f := 2042;
        ELSIF x = 11791 THEN
            sigmoid_f := 2042;
        ELSIF x = 11792 THEN
            sigmoid_f := 2042;
        ELSIF x = 11793 THEN
            sigmoid_f := 2042;
        ELSIF x = 11794 THEN
            sigmoid_f := 2042;
        ELSIF x = 11795 THEN
            sigmoid_f := 2042;
        ELSIF x = 11796 THEN
            sigmoid_f := 2042;
        ELSIF x = 11797 THEN
            sigmoid_f := 2042;
        ELSIF x = 11798 THEN
            sigmoid_f := 2042;
        ELSIF x = 11799 THEN
            sigmoid_f := 2042;
        ELSIF x = 11800 THEN
            sigmoid_f := 2042;
        ELSIF x = 11801 THEN
            sigmoid_f := 2042;
        ELSIF x = 11802 THEN
            sigmoid_f := 2042;
        ELSIF x = 11803 THEN
            sigmoid_f := 2042;
        ELSIF x = 11804 THEN
            sigmoid_f := 2042;
        ELSIF x = 11805 THEN
            sigmoid_f := 2042;
        ELSIF x = 11806 THEN
            sigmoid_f := 2042;
        ELSIF x = 11807 THEN
            sigmoid_f := 2042;
        ELSIF x = 11808 THEN
            sigmoid_f := 2042;
        ELSIF x = 11809 THEN
            sigmoid_f := 2042;
        ELSIF x = 11810 THEN
            sigmoid_f := 2042;
        ELSIF x = 11811 THEN
            sigmoid_f := 2042;
        ELSIF x = 11812 THEN
            sigmoid_f := 2042;
        ELSIF x = 11813 THEN
            sigmoid_f := 2042;
        ELSIF x = 11814 THEN
            sigmoid_f := 2042;
        ELSIF x = 11815 THEN
            sigmoid_f := 2042;
        ELSIF x = 11816 THEN
            sigmoid_f := 2042;
        ELSIF x = 11817 THEN
            sigmoid_f := 2042;
        ELSIF x = 11818 THEN
            sigmoid_f := 2042;
        ELSIF x = 11819 THEN
            sigmoid_f := 2042;
        ELSIF x = 11820 THEN
            sigmoid_f := 2042;
        ELSIF x = 11821 THEN
            sigmoid_f := 2042;
        ELSIF x = 11822 THEN
            sigmoid_f := 2042;
        ELSIF x = 11823 THEN
            sigmoid_f := 2042;
        ELSIF x = 11824 THEN
            sigmoid_f := 2042;
        ELSIF x = 11825 THEN
            sigmoid_f := 2042;
        ELSIF x = 11826 THEN
            sigmoid_f := 2042;
        ELSIF x = 11827 THEN
            sigmoid_f := 2042;
        ELSIF x = 11828 THEN
            sigmoid_f := 2042;
        ELSIF x = 11829 THEN
            sigmoid_f := 2042;
        ELSIF x = 11830 THEN
            sigmoid_f := 2042;
        ELSIF x = 11831 THEN
            sigmoid_f := 2042;
        ELSIF x = 11832 THEN
            sigmoid_f := 2042;
        ELSIF x = 11833 THEN
            sigmoid_f := 2042;
        ELSIF x = 11834 THEN
            sigmoid_f := 2042;
        ELSIF x = 11835 THEN
            sigmoid_f := 2042;
        ELSIF x = 11836 THEN
            sigmoid_f := 2042;
        ELSIF x = 11837 THEN
            sigmoid_f := 2042;
        ELSIF x = 11838 THEN
            sigmoid_f := 2042;
        ELSIF x = 11839 THEN
            sigmoid_f := 2042;
        ELSIF x = 11840 THEN
            sigmoid_f := 2042;
        ELSIF x = 11841 THEN
            sigmoid_f := 2042;
        ELSIF x = 11842 THEN
            sigmoid_f := 2042;
        ELSIF x = 11843 THEN
            sigmoid_f := 2042;
        ELSIF x = 11844 THEN
            sigmoid_f := 2042;
        ELSIF x = 11845 THEN
            sigmoid_f := 2042;
        ELSIF x = 11846 THEN
            sigmoid_f := 2042;
        ELSIF x = 11847 THEN
            sigmoid_f := 2042;
        ELSIF x = 11848 THEN
            sigmoid_f := 2042;
        ELSIF x = 11849 THEN
            sigmoid_f := 2042;
        ELSIF x = 11850 THEN
            sigmoid_f := 2042;
        ELSIF x = 11851 THEN
            sigmoid_f := 2042;
        ELSIF x = 11852 THEN
            sigmoid_f := 2042;
        ELSIF x = 11853 THEN
            sigmoid_f := 2042;
        ELSIF x = 11854 THEN
            sigmoid_f := 2042;
        ELSIF x = 11855 THEN
            sigmoid_f := 2042;
        ELSIF x = 11856 THEN
            sigmoid_f := 2042;
        ELSIF x = 11857 THEN
            sigmoid_f := 2042;
        ELSIF x = 11858 THEN
            sigmoid_f := 2042;
        ELSIF x = 11859 THEN
            sigmoid_f := 2042;
        ELSIF x = 11860 THEN
            sigmoid_f := 2042;
        ELSIF x = 11861 THEN
            sigmoid_f := 2042;
        ELSIF x = 11862 THEN
            sigmoid_f := 2042;
        ELSIF x = 11863 THEN
            sigmoid_f := 2042;
        ELSIF x = 11864 THEN
            sigmoid_f := 2042;
        ELSIF x = 11865 THEN
            sigmoid_f := 2042;
        ELSIF x = 11866 THEN
            sigmoid_f := 2042;
        ELSIF x = 11867 THEN
            sigmoid_f := 2042;
        ELSIF x = 11868 THEN
            sigmoid_f := 2042;
        ELSIF x = 11869 THEN
            sigmoid_f := 2042;
        ELSIF x = 11870 THEN
            sigmoid_f := 2042;
        ELSIF x = 11871 THEN
            sigmoid_f := 2042;
        ELSIF x = 11872 THEN
            sigmoid_f := 2042;
        ELSIF x = 11873 THEN
            sigmoid_f := 2042;
        ELSIF x = 11874 THEN
            sigmoid_f := 2042;
        ELSIF x = 11875 THEN
            sigmoid_f := 2042;
        ELSIF x = 11876 THEN
            sigmoid_f := 2042;
        ELSIF x = 11877 THEN
            sigmoid_f := 2042;
        ELSIF x = 11878 THEN
            sigmoid_f := 2042;
        ELSIF x = 11879 THEN
            sigmoid_f := 2042;
        ELSIF x = 11880 THEN
            sigmoid_f := 2042;
        ELSIF x = 11881 THEN
            sigmoid_f := 2042;
        ELSIF x = 11882 THEN
            sigmoid_f := 2042;
        ELSIF x = 11883 THEN
            sigmoid_f := 2042;
        ELSIF x = 11884 THEN
            sigmoid_f := 2042;
        ELSIF x = 11885 THEN
            sigmoid_f := 2042;
        ELSIF x = 11886 THEN
            sigmoid_f := 2042;
        ELSIF x = 11887 THEN
            sigmoid_f := 2042;
        ELSIF x = 11888 THEN
            sigmoid_f := 2042;
        ELSIF x = 11889 THEN
            sigmoid_f := 2042;
        ELSIF x = 11890 THEN
            sigmoid_f := 2042;
        ELSIF x = 11891 THEN
            sigmoid_f := 2042;
        ELSIF x = 11892 THEN
            sigmoid_f := 2042;
        ELSIF x = 11893 THEN
            sigmoid_f := 2042;
        ELSIF x = 11894 THEN
            sigmoid_f := 2042;
        ELSIF x = 11895 THEN
            sigmoid_f := 2042;
        ELSIF x = 11896 THEN
            sigmoid_f := 2042;
        ELSIF x = 11897 THEN
            sigmoid_f := 2042;
        ELSIF x = 11898 THEN
            sigmoid_f := 2042;
        ELSIF x = 11899 THEN
            sigmoid_f := 2042;
        ELSIF x = 11900 THEN
            sigmoid_f := 2042;
        ELSIF x = 11901 THEN
            sigmoid_f := 2042;
        ELSIF x = 11902 THEN
            sigmoid_f := 2042;
        ELSIF x = 11903 THEN
            sigmoid_f := 2042;
        ELSIF x = 11904 THEN
            sigmoid_f := 2042;
        ELSIF x = 11905 THEN
            sigmoid_f := 2042;
        ELSIF x = 11906 THEN
            sigmoid_f := 2042;
        ELSIF x = 11907 THEN
            sigmoid_f := 2042;
        ELSIF x = 11908 THEN
            sigmoid_f := 2042;
        ELSIF x = 11909 THEN
            sigmoid_f := 2042;
        ELSIF x = 11910 THEN
            sigmoid_f := 2042;
        ELSIF x = 11911 THEN
            sigmoid_f := 2042;
        ELSIF x = 11912 THEN
            sigmoid_f := 2042;
        ELSIF x = 11913 THEN
            sigmoid_f := 2042;
        ELSIF x = 11914 THEN
            sigmoid_f := 2042;
        ELSIF x = 11915 THEN
            sigmoid_f := 2042;
        ELSIF x = 11916 THEN
            sigmoid_f := 2042;
        ELSIF x = 11917 THEN
            sigmoid_f := 2042;
        ELSIF x = 11918 THEN
            sigmoid_f := 2042;
        ELSIF x = 11919 THEN
            sigmoid_f := 2042;
        ELSIF x = 11920 THEN
            sigmoid_f := 2042;
        ELSIF x = 11921 THEN
            sigmoid_f := 2042;
        ELSIF x = 11922 THEN
            sigmoid_f := 2042;
        ELSIF x = 11923 THEN
            sigmoid_f := 2042;
        ELSIF x = 11924 THEN
            sigmoid_f := 2042;
        ELSIF x = 11925 THEN
            sigmoid_f := 2042;
        ELSIF x = 11926 THEN
            sigmoid_f := 2042;
        ELSIF x = 11927 THEN
            sigmoid_f := 2042;
        ELSIF x = 11928 THEN
            sigmoid_f := 2042;
        ELSIF x = 11929 THEN
            sigmoid_f := 2042;
        ELSIF x = 11930 THEN
            sigmoid_f := 2042;
        ELSIF x = 11931 THEN
            sigmoid_f := 2042;
        ELSIF x = 11932 THEN
            sigmoid_f := 2042;
        ELSIF x = 11933 THEN
            sigmoid_f := 2042;
        ELSIF x = 11934 THEN
            sigmoid_f := 2042;
        ELSIF x = 11935 THEN
            sigmoid_f := 2042;
        ELSIF x = 11936 THEN
            sigmoid_f := 2042;
        ELSIF x = 11937 THEN
            sigmoid_f := 2042;
        ELSIF x = 11938 THEN
            sigmoid_f := 2042;
        ELSIF x = 11939 THEN
            sigmoid_f := 2042;
        ELSIF x = 11940 THEN
            sigmoid_f := 2042;
        ELSIF x = 11941 THEN
            sigmoid_f := 2042;
        ELSIF x = 11942 THEN
            sigmoid_f := 2042;
        ELSIF x = 11943 THEN
            sigmoid_f := 2042;
        ELSIF x = 11944 THEN
            sigmoid_f := 2042;
        ELSIF x = 11945 THEN
            sigmoid_f := 2042;
        ELSIF x = 11946 THEN
            sigmoid_f := 2042;
        ELSIF x = 11947 THEN
            sigmoid_f := 2042;
        ELSIF x = 11948 THEN
            sigmoid_f := 2042;
        ELSIF x = 11949 THEN
            sigmoid_f := 2042;
        ELSIF x = 11950 THEN
            sigmoid_f := 2042;
        ELSIF x = 11951 THEN
            sigmoid_f := 2042;
        ELSIF x = 11952 THEN
            sigmoid_f := 2042;
        ELSIF x = 11953 THEN
            sigmoid_f := 2042;
        ELSIF x = 11954 THEN
            sigmoid_f := 2042;
        ELSIF x = 11955 THEN
            sigmoid_f := 2042;
        ELSIF x = 11956 THEN
            sigmoid_f := 2042;
        ELSIF x = 11957 THEN
            sigmoid_f := 2042;
        ELSIF x = 11958 THEN
            sigmoid_f := 2042;
        ELSIF x = 11959 THEN
            sigmoid_f := 2042;
        ELSIF x = 11960 THEN
            sigmoid_f := 2042;
        ELSIF x = 11961 THEN
            sigmoid_f := 2042;
        ELSIF x = 11962 THEN
            sigmoid_f := 2042;
        ELSIF x = 11963 THEN
            sigmoid_f := 2042;
        ELSIF x = 11964 THEN
            sigmoid_f := 2042;
        ELSIF x = 11965 THEN
            sigmoid_f := 2042;
        ELSIF x = 11966 THEN
            sigmoid_f := 2042;
        ELSIF x = 11967 THEN
            sigmoid_f := 2042;
        ELSIF x = 11968 THEN
            sigmoid_f := 2042;
        ELSIF x = 11969 THEN
            sigmoid_f := 2042;
        ELSIF x = 11970 THEN
            sigmoid_f := 2042;
        ELSIF x = 11971 THEN
            sigmoid_f := 2042;
        ELSIF x = 11972 THEN
            sigmoid_f := 2042;
        ELSIF x = 11973 THEN
            sigmoid_f := 2042;
        ELSIF x = 11974 THEN
            sigmoid_f := 2042;
        ELSIF x = 11975 THEN
            sigmoid_f := 2042;
        ELSIF x = 11976 THEN
            sigmoid_f := 2042;
        ELSIF x = 11977 THEN
            sigmoid_f := 2042;
        ELSIF x = 11978 THEN
            sigmoid_f := 2042;
        ELSIF x = 11979 THEN
            sigmoid_f := 2042;
        ELSIF x = 11980 THEN
            sigmoid_f := 2042;
        ELSIF x = 11981 THEN
            sigmoid_f := 2042;
        ELSIF x = 11982 THEN
            sigmoid_f := 2042;
        ELSIF x = 11983 THEN
            sigmoid_f := 2042;
        ELSIF x = 11984 THEN
            sigmoid_f := 2042;
        ELSIF x = 11985 THEN
            sigmoid_f := 2042;
        ELSIF x = 11986 THEN
            sigmoid_f := 2042;
        ELSIF x = 11987 THEN
            sigmoid_f := 2042;
        ELSIF x = 11988 THEN
            sigmoid_f := 2042;
        ELSIF x = 11989 THEN
            sigmoid_f := 2042;
        ELSIF x = 11990 THEN
            sigmoid_f := 2042;
        ELSIF x = 11991 THEN
            sigmoid_f := 2042;
        ELSIF x = 11992 THEN
            sigmoid_f := 2042;
        ELSIF x = 11993 THEN
            sigmoid_f := 2042;
        ELSIF x = 11994 THEN
            sigmoid_f := 2042;
        ELSIF x = 11995 THEN
            sigmoid_f := 2042;
        ELSIF x = 11996 THEN
            sigmoid_f := 2042;
        ELSIF x = 11997 THEN
            sigmoid_f := 2042;
        ELSIF x = 11998 THEN
            sigmoid_f := 2042;
        ELSIF x = 11999 THEN
            sigmoid_f := 2042;
        ELSIF x = 12000 THEN
            sigmoid_f := 2042;
        ELSIF x = 12001 THEN
            sigmoid_f := 2042;
        ELSIF x = 12002 THEN
            sigmoid_f := 2042;
        ELSIF x = 12003 THEN
            sigmoid_f := 2042;
        ELSIF x = 12004 THEN
            sigmoid_f := 2042;
        ELSIF x = 12005 THEN
            sigmoid_f := 2042;
        ELSIF x = 12006 THEN
            sigmoid_f := 2042;
        ELSIF x = 12007 THEN
            sigmoid_f := 2042;
        ELSIF x = 12008 THEN
            sigmoid_f := 2042;
        ELSIF x = 12009 THEN
            sigmoid_f := 2042;
        ELSIF x = 12010 THEN
            sigmoid_f := 2042;
        ELSIF x = 12011 THEN
            sigmoid_f := 2042;
        ELSIF x = 12012 THEN
            sigmoid_f := 2042;
        ELSIF x = 12013 THEN
            sigmoid_f := 2042;
        ELSIF x = 12014 THEN
            sigmoid_f := 2042;
        ELSIF x = 12015 THEN
            sigmoid_f := 2042;
        ELSIF x = 12016 THEN
            sigmoid_f := 2042;
        ELSIF x = 12017 THEN
            sigmoid_f := 2042;
        ELSIF x = 12018 THEN
            sigmoid_f := 2042;
        ELSIF x = 12019 THEN
            sigmoid_f := 2042;
        ELSIF x = 12020 THEN
            sigmoid_f := 2042;
        ELSIF x = 12021 THEN
            sigmoid_f := 2042;
        ELSIF x = 12022 THEN
            sigmoid_f := 2042;
        ELSIF x = 12023 THEN
            sigmoid_f := 2042;
        ELSIF x = 12024 THEN
            sigmoid_f := 2042;
        ELSIF x = 12025 THEN
            sigmoid_f := 2042;
        ELSIF x = 12026 THEN
            sigmoid_f := 2042;
        ELSIF x = 12027 THEN
            sigmoid_f := 2042;
        ELSIF x = 12028 THEN
            sigmoid_f := 2042;
        ELSIF x = 12029 THEN
            sigmoid_f := 2042;
        ELSIF x = 12030 THEN
            sigmoid_f := 2042;
        ELSIF x = 12031 THEN
            sigmoid_f := 2042;
        ELSIF x = 12032 THEN
            sigmoid_f := 2042;
        ELSIF x = 12033 THEN
            sigmoid_f := 2042;
        ELSIF x = 12034 THEN
            sigmoid_f := 2042;
        ELSIF x = 12035 THEN
            sigmoid_f := 2042;
        ELSIF x = 12036 THEN
            sigmoid_f := 2042;
        ELSIF x = 12037 THEN
            sigmoid_f := 2042;
        ELSIF x = 12038 THEN
            sigmoid_f := 2042;
        ELSIF x = 12039 THEN
            sigmoid_f := 2042;
        ELSIF x = 12040 THEN
            sigmoid_f := 2042;
        ELSIF x = 12041 THEN
            sigmoid_f := 2042;
        ELSIF x = 12042 THEN
            sigmoid_f := 2042;
        ELSIF x = 12043 THEN
            sigmoid_f := 2042;
        ELSIF x = 12044 THEN
            sigmoid_f := 2042;
        ELSIF x = 12045 THEN
            sigmoid_f := 2042;
        ELSIF x = 12046 THEN
            sigmoid_f := 2042;
        ELSIF x = 12047 THEN
            sigmoid_f := 2042;
        ELSIF x = 12048 THEN
            sigmoid_f := 2042;
        ELSIF x = 12049 THEN
            sigmoid_f := 2042;
        ELSIF x = 12050 THEN
            sigmoid_f := 2042;
        ELSIF x = 12051 THEN
            sigmoid_f := 2042;
        ELSIF x = 12052 THEN
            sigmoid_f := 2042;
        ELSIF x = 12053 THEN
            sigmoid_f := 2042;
        ELSIF x = 12054 THEN
            sigmoid_f := 2042;
        ELSIF x = 12055 THEN
            sigmoid_f := 2042;
        ELSIF x = 12056 THEN
            sigmoid_f := 2042;
        ELSIF x = 12057 THEN
            sigmoid_f := 2042;
        ELSIF x = 12058 THEN
            sigmoid_f := 2042;
        ELSIF x = 12059 THEN
            sigmoid_f := 2042;
        ELSIF x = 12060 THEN
            sigmoid_f := 2042;
        ELSIF x = 12061 THEN
            sigmoid_f := 2042;
        ELSIF x = 12062 THEN
            sigmoid_f := 2042;
        ELSIF x = 12063 THEN
            sigmoid_f := 2042;
        ELSIF x = 12064 THEN
            sigmoid_f := 2042;
        ELSIF x = 12065 THEN
            sigmoid_f := 2042;
        ELSIF x = 12066 THEN
            sigmoid_f := 2042;
        ELSIF x = 12067 THEN
            sigmoid_f := 2042;
        ELSIF x = 12068 THEN
            sigmoid_f := 2042;
        ELSIF x = 12069 THEN
            sigmoid_f := 2042;
        ELSIF x = 12070 THEN
            sigmoid_f := 2042;
        ELSIF x = 12071 THEN
            sigmoid_f := 2042;
        ELSIF x = 12072 THEN
            sigmoid_f := 2042;
        ELSIF x = 12073 THEN
            sigmoid_f := 2042;
        ELSIF x = 12074 THEN
            sigmoid_f := 2042;
        ELSIF x = 12075 THEN
            sigmoid_f := 2042;
        ELSIF x = 12076 THEN
            sigmoid_f := 2042;
        ELSIF x = 12077 THEN
            sigmoid_f := 2042;
        ELSIF x = 12078 THEN
            sigmoid_f := 2042;
        ELSIF x = 12079 THEN
            sigmoid_f := 2042;
        ELSIF x = 12080 THEN
            sigmoid_f := 2042;
        ELSIF x = 12081 THEN
            sigmoid_f := 2042;
        ELSIF x = 12082 THEN
            sigmoid_f := 2042;
        ELSIF x = 12083 THEN
            sigmoid_f := 2042;
        ELSIF x = 12084 THEN
            sigmoid_f := 2042;
        ELSIF x = 12085 THEN
            sigmoid_f := 2042;
        ELSIF x = 12086 THEN
            sigmoid_f := 2042;
        ELSIF x = 12087 THEN
            sigmoid_f := 2042;
        ELSIF x = 12088 THEN
            sigmoid_f := 2042;
        ELSIF x = 12089 THEN
            sigmoid_f := 2042;
        ELSIF x = 12090 THEN
            sigmoid_f := 2042;
        ELSIF x = 12091 THEN
            sigmoid_f := 2042;
        ELSIF x = 12092 THEN
            sigmoid_f := 2042;
        ELSIF x = 12093 THEN
            sigmoid_f := 2042;
        ELSIF x = 12094 THEN
            sigmoid_f := 2042;
        ELSIF x = 12095 THEN
            sigmoid_f := 2042;
        ELSIF x = 12096 THEN
            sigmoid_f := 2042;
        ELSIF x = 12097 THEN
            sigmoid_f := 2042;
        ELSIF x = 12098 THEN
            sigmoid_f := 2042;
        ELSIF x = 12099 THEN
            sigmoid_f := 2042;
        ELSIF x = 12100 THEN
            sigmoid_f := 2042;
        ELSIF x = 12101 THEN
            sigmoid_f := 2042;
        ELSIF x = 12102 THEN
            sigmoid_f := 2042;
        ELSIF x = 12103 THEN
            sigmoid_f := 2042;
        ELSIF x = 12104 THEN
            sigmoid_f := 2042;
        ELSIF x = 12105 THEN
            sigmoid_f := 2042;
        ELSIF x = 12106 THEN
            sigmoid_f := 2042;
        ELSIF x = 12107 THEN
            sigmoid_f := 2042;
        ELSIF x = 12108 THEN
            sigmoid_f := 2042;
        ELSIF x = 12109 THEN
            sigmoid_f := 2042;
        ELSIF x = 12110 THEN
            sigmoid_f := 2042;
        ELSIF x = 12111 THEN
            sigmoid_f := 2042;
        ELSIF x = 12112 THEN
            sigmoid_f := 2042;
        ELSIF x = 12113 THEN
            sigmoid_f := 2042;
        ELSIF x = 12114 THEN
            sigmoid_f := 2042;
        ELSIF x = 12115 THEN
            sigmoid_f := 2042;
        ELSIF x = 12116 THEN
            sigmoid_f := 2042;
        ELSIF x = 12117 THEN
            sigmoid_f := 2042;
        ELSIF x = 12118 THEN
            sigmoid_f := 2042;
        ELSIF x = 12119 THEN
            sigmoid_f := 2042;
        ELSIF x = 12120 THEN
            sigmoid_f := 2042;
        ELSIF x = 12121 THEN
            sigmoid_f := 2042;
        ELSIF x = 12122 THEN
            sigmoid_f := 2042;
        ELSIF x = 12123 THEN
            sigmoid_f := 2042;
        ELSIF x = 12124 THEN
            sigmoid_f := 2042;
        ELSIF x = 12125 THEN
            sigmoid_f := 2042;
        ELSIF x = 12126 THEN
            sigmoid_f := 2042;
        ELSIF x = 12127 THEN
            sigmoid_f := 2042;
        ELSIF x = 12128 THEN
            sigmoid_f := 2042;
        ELSIF x = 12129 THEN
            sigmoid_f := 2042;
        ELSIF x = 12130 THEN
            sigmoid_f := 2042;
        ELSIF x = 12131 THEN
            sigmoid_f := 2042;
        ELSIF x = 12132 THEN
            sigmoid_f := 2042;
        ELSIF x = 12133 THEN
            sigmoid_f := 2042;
        ELSIF x = 12134 THEN
            sigmoid_f := 2042;
        ELSIF x = 12135 THEN
            sigmoid_f := 2042;
        ELSIF x = 12136 THEN
            sigmoid_f := 2042;
        ELSIF x = 12137 THEN
            sigmoid_f := 2042;
        ELSIF x = 12138 THEN
            sigmoid_f := 2042;
        ELSIF x = 12139 THEN
            sigmoid_f := 2042;
        ELSIF x = 12140 THEN
            sigmoid_f := 2042;
        ELSIF x = 12141 THEN
            sigmoid_f := 2042;
        ELSIF x = 12142 THEN
            sigmoid_f := 2042;
        ELSIF x = 12143 THEN
            sigmoid_f := 2042;
        ELSIF x = 12144 THEN
            sigmoid_f := 2042;
        ELSIF x = 12145 THEN
            sigmoid_f := 2042;
        ELSIF x = 12146 THEN
            sigmoid_f := 2042;
        ELSIF x = 12147 THEN
            sigmoid_f := 2042;
        ELSIF x = 12148 THEN
            sigmoid_f := 2042;
        ELSIF x = 12149 THEN
            sigmoid_f := 2042;
        ELSIF x = 12150 THEN
            sigmoid_f := 2042;
        ELSIF x = 12151 THEN
            sigmoid_f := 2042;
        ELSIF x = 12152 THEN
            sigmoid_f := 2042;
        ELSIF x = 12153 THEN
            sigmoid_f := 2042;
        ELSIF x = 12154 THEN
            sigmoid_f := 2042;
        ELSIF x = 12155 THEN
            sigmoid_f := 2042;
        ELSIF x = 12156 THEN
            sigmoid_f := 2042;
        ELSIF x = 12157 THEN
            sigmoid_f := 2042;
        ELSIF x = 12158 THEN
            sigmoid_f := 2042;
        ELSIF x = 12159 THEN
            sigmoid_f := 2042;
        ELSIF x = 12160 THEN
            sigmoid_f := 2042;
        ELSIF x = 12161 THEN
            sigmoid_f := 2042;
        ELSIF x = 12162 THEN
            sigmoid_f := 2042;
        ELSIF x = 12163 THEN
            sigmoid_f := 2042;
        ELSIF x = 12164 THEN
            sigmoid_f := 2042;
        ELSIF x = 12165 THEN
            sigmoid_f := 2042;
        ELSIF x = 12166 THEN
            sigmoid_f := 2042;
        ELSIF x = 12167 THEN
            sigmoid_f := 2042;
        ELSIF x = 12168 THEN
            sigmoid_f := 2042;
        ELSIF x = 12169 THEN
            sigmoid_f := 2042;
        ELSIF x = 12170 THEN
            sigmoid_f := 2042;
        ELSIF x = 12171 THEN
            sigmoid_f := 2042;
        ELSIF x = 12172 THEN
            sigmoid_f := 2042;
        ELSIF x = 12173 THEN
            sigmoid_f := 2042;
        ELSIF x = 12174 THEN
            sigmoid_f := 2042;
        ELSIF x = 12175 THEN
            sigmoid_f := 2042;
        ELSIF x = 12176 THEN
            sigmoid_f := 2042;
        ELSIF x = 12177 THEN
            sigmoid_f := 2042;
        ELSIF x = 12178 THEN
            sigmoid_f := 2042;
        ELSIF x = 12179 THEN
            sigmoid_f := 2042;
        ELSIF x = 12180 THEN
            sigmoid_f := 2042;
        ELSIF x = 12181 THEN
            sigmoid_f := 2042;
        ELSIF x = 12182 THEN
            sigmoid_f := 2042;
        ELSIF x = 12183 THEN
            sigmoid_f := 2042;
        ELSIF x = 12184 THEN
            sigmoid_f := 2042;
        ELSIF x = 12185 THEN
            sigmoid_f := 2042;
        ELSIF x = 12186 THEN
            sigmoid_f := 2042;
        ELSIF x = 12187 THEN
            sigmoid_f := 2042;
        ELSIF x = 12188 THEN
            sigmoid_f := 2042;
        ELSIF x = 12189 THEN
            sigmoid_f := 2042;
        ELSIF x = 12190 THEN
            sigmoid_f := 2042;
        ELSIF x = 12191 THEN
            sigmoid_f := 2042;
        ELSIF x = 12192 THEN
            sigmoid_f := 2042;
        ELSIF x = 12193 THEN
            sigmoid_f := 2042;
        ELSIF x = 12194 THEN
            sigmoid_f := 2042;
        ELSIF x = 12195 THEN
            sigmoid_f := 2042;
        ELSIF x = 12196 THEN
            sigmoid_f := 2042;
        ELSIF x = 12197 THEN
            sigmoid_f := 2042;
        ELSIF x = 12198 THEN
            sigmoid_f := 2042;
        ELSIF x = 12199 THEN
            sigmoid_f := 2042;
        ELSIF x = 12200 THEN
            sigmoid_f := 2042;
        ELSIF x = 12201 THEN
            sigmoid_f := 2042;
        ELSIF x = 12202 THEN
            sigmoid_f := 2042;
        ELSIF x = 12203 THEN
            sigmoid_f := 2042;
        ELSIF x = 12204 THEN
            sigmoid_f := 2042;
        ELSIF x = 12205 THEN
            sigmoid_f := 2042;
        ELSIF x = 12206 THEN
            sigmoid_f := 2042;
        ELSIF x = 12207 THEN
            sigmoid_f := 2042;
        ELSIF x = 12208 THEN
            sigmoid_f := 2042;
        ELSIF x = 12209 THEN
            sigmoid_f := 2042;
        ELSIF x = 12210 THEN
            sigmoid_f := 2042;
        ELSIF x = 12211 THEN
            sigmoid_f := 2042;
        ELSIF x = 12212 THEN
            sigmoid_f := 2042;
        ELSIF x = 12213 THEN
            sigmoid_f := 2042;
        ELSIF x = 12214 THEN
            sigmoid_f := 2042;
        ELSIF x = 12215 THEN
            sigmoid_f := 2042;
        ELSIF x = 12216 THEN
            sigmoid_f := 2042;
        ELSIF x = 12217 THEN
            sigmoid_f := 2042;
        ELSIF x = 12218 THEN
            sigmoid_f := 2042;
        ELSIF x = 12219 THEN
            sigmoid_f := 2042;
        ELSIF x = 12220 THEN
            sigmoid_f := 2042;
        ELSIF x = 12221 THEN
            sigmoid_f := 2042;
        ELSIF x = 12222 THEN
            sigmoid_f := 2042;
        ELSIF x = 12223 THEN
            sigmoid_f := 2042;
        ELSIF x = 12224 THEN
            sigmoid_f := 2042;
        ELSIF x = 12225 THEN
            sigmoid_f := 2042;
        ELSIF x = 12226 THEN
            sigmoid_f := 2042;
        ELSIF x = 12227 THEN
            sigmoid_f := 2042;
        ELSIF x = 12228 THEN
            sigmoid_f := 2042;
        ELSIF x = 12229 THEN
            sigmoid_f := 2042;
        ELSIF x = 12230 THEN
            sigmoid_f := 2042;
        ELSIF x = 12231 THEN
            sigmoid_f := 2042;
        ELSIF x = 12232 THEN
            sigmoid_f := 2042;
        ELSIF x = 12233 THEN
            sigmoid_f := 2042;
        ELSIF x = 12234 THEN
            sigmoid_f := 2042;
        ELSIF x = 12235 THEN
            sigmoid_f := 2042;
        ELSIF x = 12236 THEN
            sigmoid_f := 2042;
        ELSIF x = 12237 THEN
            sigmoid_f := 2042;
        ELSIF x = 12238 THEN
            sigmoid_f := 2042;
        ELSIF x = 12239 THEN
            sigmoid_f := 2042;
        ELSIF x = 12240 THEN
            sigmoid_f := 2042;
        ELSIF x = 12241 THEN
            sigmoid_f := 2042;
        ELSIF x = 12242 THEN
            sigmoid_f := 2042;
        ELSIF x = 12243 THEN
            sigmoid_f := 2042;
        ELSIF x = 12244 THEN
            sigmoid_f := 2042;
        ELSIF x = 12245 THEN
            sigmoid_f := 2042;
        ELSIF x = 12246 THEN
            sigmoid_f := 2042;
        ELSIF x = 12247 THEN
            sigmoid_f := 2042;
        ELSIF x = 12248 THEN
            sigmoid_f := 2042;
        ELSIF x = 12249 THEN
            sigmoid_f := 2042;
        ELSIF x = 12250 THEN
            sigmoid_f := 2042;
        ELSIF x = 12251 THEN
            sigmoid_f := 2042;
        ELSIF x = 12252 THEN
            sigmoid_f := 2042;
        ELSIF x = 12253 THEN
            sigmoid_f := 2042;
        ELSIF x = 12254 THEN
            sigmoid_f := 2042;
        ELSIF x = 12255 THEN
            sigmoid_f := 2042;
        ELSIF x = 12256 THEN
            sigmoid_f := 2042;
        ELSIF x = 12257 THEN
            sigmoid_f := 2042;
        ELSIF x = 12258 THEN
            sigmoid_f := 2042;
        ELSIF x = 12259 THEN
            sigmoid_f := 2042;
        ELSIF x = 12260 THEN
            sigmoid_f := 2042;
        ELSIF x = 12261 THEN
            sigmoid_f := 2042;
        ELSIF x = 12262 THEN
            sigmoid_f := 2042;
        ELSIF x = 12263 THEN
            sigmoid_f := 2042;
        ELSIF x = 12264 THEN
            sigmoid_f := 2042;
        ELSIF x = 12265 THEN
            sigmoid_f := 2042;
        ELSIF x = 12266 THEN
            sigmoid_f := 2042;
        ELSIF x = 12267 THEN
            sigmoid_f := 2042;
        ELSIF x = 12268 THEN
            sigmoid_f := 2042;
        ELSIF x = 12269 THEN
            sigmoid_f := 2042;
        ELSIF x = 12270 THEN
            sigmoid_f := 2042;
        ELSIF x = 12271 THEN
            sigmoid_f := 2042;
        ELSIF x = 12272 THEN
            sigmoid_f := 2042;
        ELSIF x = 12273 THEN
            sigmoid_f := 2042;
        ELSIF x = 12274 THEN
            sigmoid_f := 2042;
        ELSIF x = 12275 THEN
            sigmoid_f := 2042;
        ELSIF x = 12276 THEN
            sigmoid_f := 2042;
        ELSIF x = 12277 THEN
            sigmoid_f := 2042;
        ELSIF x = 12278 THEN
            sigmoid_f := 2042;
        ELSIF x = 12279 THEN
            sigmoid_f := 2042;
        ELSIF x = 12280 THEN
            sigmoid_f := 2042;
        ELSIF x = 12281 THEN
            sigmoid_f := 2042;
        ELSIF x = 12282 THEN
            sigmoid_f := 2042;
        ELSIF x = 12283 THEN
            sigmoid_f := 2042;
        ELSIF x = 12284 THEN
            sigmoid_f := 2042;
        ELSIF x = 12285 THEN
            sigmoid_f := 2042;
        ELSIF x = 12286 THEN
            sigmoid_f := 2042;
        ELSIF x = 12287 THEN
            sigmoid_f := 2042;
        ELSIF x = 12288 THEN
            sigmoid_f := 2044;
        ELSIF x = 12289 THEN
            sigmoid_f := 2044;
        ELSIF x = 12290 THEN
            sigmoid_f := 2044;
        ELSIF x = 12291 THEN
            sigmoid_f := 2044;
        ELSIF x = 12292 THEN
            sigmoid_f := 2044;
        ELSIF x = 12293 THEN
            sigmoid_f := 2044;
        ELSIF x = 12294 THEN
            sigmoid_f := 2044;
        ELSIF x = 12295 THEN
            sigmoid_f := 2044;
        ELSIF x = 12296 THEN
            sigmoid_f := 2044;
        ELSIF x = 12297 THEN
            sigmoid_f := 2044;
        ELSIF x = 12298 THEN
            sigmoid_f := 2044;
        ELSIF x = 12299 THEN
            sigmoid_f := 2044;
        ELSIF x = 12300 THEN
            sigmoid_f := 2044;
        ELSIF x = 12301 THEN
            sigmoid_f := 2044;
        ELSIF x = 12302 THEN
            sigmoid_f := 2044;
        ELSIF x = 12303 THEN
            sigmoid_f := 2044;
        ELSIF x = 12304 THEN
            sigmoid_f := 2044;
        ELSIF x = 12305 THEN
            sigmoid_f := 2044;
        ELSIF x = 12306 THEN
            sigmoid_f := 2044;
        ELSIF x = 12307 THEN
            sigmoid_f := 2044;
        ELSIF x = 12308 THEN
            sigmoid_f := 2044;
        ELSIF x = 12309 THEN
            sigmoid_f := 2044;
        ELSIF x = 12310 THEN
            sigmoid_f := 2044;
        ELSIF x = 12311 THEN
            sigmoid_f := 2044;
        ELSIF x = 12312 THEN
            sigmoid_f := 2044;
        ELSIF x = 12313 THEN
            sigmoid_f := 2044;
        ELSIF x = 12314 THEN
            sigmoid_f := 2044;
        ELSIF x = 12315 THEN
            sigmoid_f := 2044;
        ELSIF x = 12316 THEN
            sigmoid_f := 2044;
        ELSIF x = 12317 THEN
            sigmoid_f := 2044;
        ELSIF x = 12318 THEN
            sigmoid_f := 2044;
        ELSIF x = 12319 THEN
            sigmoid_f := 2044;
        ELSIF x = 12320 THEN
            sigmoid_f := 2044;
        ELSIF x = 12321 THEN
            sigmoid_f := 2044;
        ELSIF x = 12322 THEN
            sigmoid_f := 2044;
        ELSIF x = 12323 THEN
            sigmoid_f := 2044;
        ELSIF x = 12324 THEN
            sigmoid_f := 2044;
        ELSIF x = 12325 THEN
            sigmoid_f := 2044;
        ELSIF x = 12326 THEN
            sigmoid_f := 2044;
        ELSIF x = 12327 THEN
            sigmoid_f := 2044;
        ELSIF x = 12328 THEN
            sigmoid_f := 2044;
        ELSIF x = 12329 THEN
            sigmoid_f := 2044;
        ELSIF x = 12330 THEN
            sigmoid_f := 2044;
        ELSIF x = 12331 THEN
            sigmoid_f := 2044;
        ELSIF x = 12332 THEN
            sigmoid_f := 2044;
        ELSIF x = 12333 THEN
            sigmoid_f := 2044;
        ELSIF x = 12334 THEN
            sigmoid_f := 2044;
        ELSIF x = 12335 THEN
            sigmoid_f := 2044;
        ELSIF x = 12336 THEN
            sigmoid_f := 2044;
        ELSIF x = 12337 THEN
            sigmoid_f := 2044;
        ELSIF x = 12338 THEN
            sigmoid_f := 2044;
        ELSIF x = 12339 THEN
            sigmoid_f := 2044;
        ELSIF x = 12340 THEN
            sigmoid_f := 2044;
        ELSIF x = 12341 THEN
            sigmoid_f := 2044;
        ELSIF x = 12342 THEN
            sigmoid_f := 2044;
        ELSIF x = 12343 THEN
            sigmoid_f := 2044;
        ELSIF x = 12344 THEN
            sigmoid_f := 2044;
        ELSIF x = 12345 THEN
            sigmoid_f := 2044;
        ELSIF x = 12346 THEN
            sigmoid_f := 2044;
        ELSIF x = 12347 THEN
            sigmoid_f := 2044;
        ELSIF x = 12348 THEN
            sigmoid_f := 2044;
        ELSIF x = 12349 THEN
            sigmoid_f := 2044;
        ELSIF x = 12350 THEN
            sigmoid_f := 2044;
        ELSIF x = 12351 THEN
            sigmoid_f := 2044;
        ELSIF x = 12352 THEN
            sigmoid_f := 2044;
        ELSIF x = 12353 THEN
            sigmoid_f := 2044;
        ELSIF x = 12354 THEN
            sigmoid_f := 2044;
        ELSIF x = 12355 THEN
            sigmoid_f := 2044;
        ELSIF x = 12356 THEN
            sigmoid_f := 2044;
        ELSIF x = 12357 THEN
            sigmoid_f := 2044;
        ELSIF x = 12358 THEN
            sigmoid_f := 2044;
        ELSIF x = 12359 THEN
            sigmoid_f := 2044;
        ELSIF x = 12360 THEN
            sigmoid_f := 2044;
        ELSIF x = 12361 THEN
            sigmoid_f := 2044;
        ELSIF x = 12362 THEN
            sigmoid_f := 2044;
        ELSIF x = 12363 THEN
            sigmoid_f := 2044;
        ELSIF x = 12364 THEN
            sigmoid_f := 2044;
        ELSIF x = 12365 THEN
            sigmoid_f := 2044;
        ELSIF x = 12366 THEN
            sigmoid_f := 2044;
        ELSIF x = 12367 THEN
            sigmoid_f := 2044;
        ELSIF x = 12368 THEN
            sigmoid_f := 2044;
        ELSIF x = 12369 THEN
            sigmoid_f := 2044;
        ELSIF x = 12370 THEN
            sigmoid_f := 2044;
        ELSIF x = 12371 THEN
            sigmoid_f := 2044;
        ELSIF x = 12372 THEN
            sigmoid_f := 2044;
        ELSIF x = 12373 THEN
            sigmoid_f := 2044;
        ELSIF x = 12374 THEN
            sigmoid_f := 2044;
        ELSIF x = 12375 THEN
            sigmoid_f := 2044;
        ELSIF x = 12376 THEN
            sigmoid_f := 2044;
        ELSIF x = 12377 THEN
            sigmoid_f := 2044;
        ELSIF x = 12378 THEN
            sigmoid_f := 2044;
        ELSIF x = 12379 THEN
            sigmoid_f := 2044;
        ELSIF x = 12380 THEN
            sigmoid_f := 2044;
        ELSIF x = 12381 THEN
            sigmoid_f := 2044;
        ELSIF x = 12382 THEN
            sigmoid_f := 2044;
        ELSIF x = 12383 THEN
            sigmoid_f := 2044;
        ELSIF x = 12384 THEN
            sigmoid_f := 2044;
        ELSIF x = 12385 THEN
            sigmoid_f := 2044;
        ELSIF x = 12386 THEN
            sigmoid_f := 2044;
        ELSIF x = 12387 THEN
            sigmoid_f := 2044;
        ELSIF x = 12388 THEN
            sigmoid_f := 2044;
        ELSIF x = 12389 THEN
            sigmoid_f := 2044;
        ELSIF x = 12390 THEN
            sigmoid_f := 2044;
        ELSIF x = 12391 THEN
            sigmoid_f := 2044;
        ELSIF x = 12392 THEN
            sigmoid_f := 2044;
        ELSIF x = 12393 THEN
            sigmoid_f := 2044;
        ELSIF x = 12394 THEN
            sigmoid_f := 2044;
        ELSIF x = 12395 THEN
            sigmoid_f := 2044;
        ELSIF x = 12396 THEN
            sigmoid_f := 2044;
        ELSIF x = 12397 THEN
            sigmoid_f := 2044;
        ELSIF x = 12398 THEN
            sigmoid_f := 2044;
        ELSIF x = 12399 THEN
            sigmoid_f := 2044;
        ELSIF x = 12400 THEN
            sigmoid_f := 2044;
        ELSIF x = 12401 THEN
            sigmoid_f := 2044;
        ELSIF x = 12402 THEN
            sigmoid_f := 2044;
        ELSIF x = 12403 THEN
            sigmoid_f := 2044;
        ELSIF x = 12404 THEN
            sigmoid_f := 2044;
        ELSIF x = 12405 THEN
            sigmoid_f := 2044;
        ELSIF x = 12406 THEN
            sigmoid_f := 2044;
        ELSIF x = 12407 THEN
            sigmoid_f := 2044;
        ELSIF x = 12408 THEN
            sigmoid_f := 2044;
        ELSIF x = 12409 THEN
            sigmoid_f := 2044;
        ELSIF x = 12410 THEN
            sigmoid_f := 2044;
        ELSIF x = 12411 THEN
            sigmoid_f := 2044;
        ELSIF x = 12412 THEN
            sigmoid_f := 2044;
        ELSIF x = 12413 THEN
            sigmoid_f := 2044;
        ELSIF x = 12414 THEN
            sigmoid_f := 2044;
        ELSIF x = 12415 THEN
            sigmoid_f := 2044;
        ELSIF x = 12416 THEN
            sigmoid_f := 2044;
        ELSIF x = 12417 THEN
            sigmoid_f := 2044;
        ELSIF x = 12418 THEN
            sigmoid_f := 2044;
        ELSIF x = 12419 THEN
            sigmoid_f := 2044;
        ELSIF x = 12420 THEN
            sigmoid_f := 2044;
        ELSIF x = 12421 THEN
            sigmoid_f := 2044;
        ELSIF x = 12422 THEN
            sigmoid_f := 2044;
        ELSIF x = 12423 THEN
            sigmoid_f := 2044;
        ELSIF x = 12424 THEN
            sigmoid_f := 2044;
        ELSIF x = 12425 THEN
            sigmoid_f := 2044;
        ELSIF x = 12426 THEN
            sigmoid_f := 2044;
        ELSIF x = 12427 THEN
            sigmoid_f := 2044;
        ELSIF x = 12428 THEN
            sigmoid_f := 2044;
        ELSIF x = 12429 THEN
            sigmoid_f := 2044;
        ELSIF x = 12430 THEN
            sigmoid_f := 2044;
        ELSIF x = 12431 THEN
            sigmoid_f := 2044;
        ELSIF x = 12432 THEN
            sigmoid_f := 2044;
        ELSIF x = 12433 THEN
            sigmoid_f := 2044;
        ELSIF x = 12434 THEN
            sigmoid_f := 2044;
        ELSIF x = 12435 THEN
            sigmoid_f := 2044;
        ELSIF x = 12436 THEN
            sigmoid_f := 2044;
        ELSIF x = 12437 THEN
            sigmoid_f := 2044;
        ELSIF x = 12438 THEN
            sigmoid_f := 2044;
        ELSIF x = 12439 THEN
            sigmoid_f := 2044;
        ELSIF x = 12440 THEN
            sigmoid_f := 2044;
        ELSIF x = 12441 THEN
            sigmoid_f := 2044;
        ELSIF x = 12442 THEN
            sigmoid_f := 2044;
        ELSIF x = 12443 THEN
            sigmoid_f := 2044;
        ELSIF x = 12444 THEN
            sigmoid_f := 2044;
        ELSIF x = 12445 THEN
            sigmoid_f := 2044;
        ELSIF x = 12446 THEN
            sigmoid_f := 2044;
        ELSIF x = 12447 THEN
            sigmoid_f := 2044;
        ELSIF x = 12448 THEN
            sigmoid_f := 2044;
        ELSIF x = 12449 THEN
            sigmoid_f := 2044;
        ELSIF x = 12450 THEN
            sigmoid_f := 2044;
        ELSIF x = 12451 THEN
            sigmoid_f := 2044;
        ELSIF x = 12452 THEN
            sigmoid_f := 2044;
        ELSIF x = 12453 THEN
            sigmoid_f := 2044;
        ELSIF x = 12454 THEN
            sigmoid_f := 2044;
        ELSIF x = 12455 THEN
            sigmoid_f := 2044;
        ELSIF x = 12456 THEN
            sigmoid_f := 2044;
        ELSIF x = 12457 THEN
            sigmoid_f := 2044;
        ELSIF x = 12458 THEN
            sigmoid_f := 2044;
        ELSIF x = 12459 THEN
            sigmoid_f := 2044;
        ELSIF x = 12460 THEN
            sigmoid_f := 2044;
        ELSIF x = 12461 THEN
            sigmoid_f := 2044;
        ELSIF x = 12462 THEN
            sigmoid_f := 2044;
        ELSIF x = 12463 THEN
            sigmoid_f := 2044;
        ELSIF x = 12464 THEN
            sigmoid_f := 2044;
        ELSIF x = 12465 THEN
            sigmoid_f := 2044;
        ELSIF x = 12466 THEN
            sigmoid_f := 2044;
        ELSIF x = 12467 THEN
            sigmoid_f := 2044;
        ELSIF x = 12468 THEN
            sigmoid_f := 2044;
        ELSIF x = 12469 THEN
            sigmoid_f := 2044;
        ELSIF x = 12470 THEN
            sigmoid_f := 2044;
        ELSIF x = 12471 THEN
            sigmoid_f := 2044;
        ELSIF x = 12472 THEN
            sigmoid_f := 2044;
        ELSIF x = 12473 THEN
            sigmoid_f := 2044;
        ELSIF x = 12474 THEN
            sigmoid_f := 2044;
        ELSIF x = 12475 THEN
            sigmoid_f := 2044;
        ELSIF x = 12476 THEN
            sigmoid_f := 2044;
        ELSIF x = 12477 THEN
            sigmoid_f := 2044;
        ELSIF x = 12478 THEN
            sigmoid_f := 2044;
        ELSIF x = 12479 THEN
            sigmoid_f := 2044;
        ELSIF x = 12480 THEN
            sigmoid_f := 2044;
        ELSIF x = 12481 THEN
            sigmoid_f := 2044;
        ELSIF x = 12482 THEN
            sigmoid_f := 2044;
        ELSIF x = 12483 THEN
            sigmoid_f := 2044;
        ELSIF x = 12484 THEN
            sigmoid_f := 2044;
        ELSIF x = 12485 THEN
            sigmoid_f := 2044;
        ELSIF x = 12486 THEN
            sigmoid_f := 2044;
        ELSIF x = 12487 THEN
            sigmoid_f := 2044;
        ELSIF x = 12488 THEN
            sigmoid_f := 2044;
        ELSIF x = 12489 THEN
            sigmoid_f := 2044;
        ELSIF x = 12490 THEN
            sigmoid_f := 2044;
        ELSIF x = 12491 THEN
            sigmoid_f := 2044;
        ELSIF x = 12492 THEN
            sigmoid_f := 2044;
        ELSIF x = 12493 THEN
            sigmoid_f := 2044;
        ELSIF x = 12494 THEN
            sigmoid_f := 2044;
        ELSIF x = 12495 THEN
            sigmoid_f := 2044;
        ELSIF x = 12496 THEN
            sigmoid_f := 2044;
        ELSIF x = 12497 THEN
            sigmoid_f := 2044;
        ELSIF x = 12498 THEN
            sigmoid_f := 2044;
        ELSIF x = 12499 THEN
            sigmoid_f := 2044;
        ELSIF x = 12500 THEN
            sigmoid_f := 2044;
        ELSIF x = 12501 THEN
            sigmoid_f := 2044;
        ELSIF x = 12502 THEN
            sigmoid_f := 2044;
        ELSIF x = 12503 THEN
            sigmoid_f := 2044;
        ELSIF x = 12504 THEN
            sigmoid_f := 2044;
        ELSIF x = 12505 THEN
            sigmoid_f := 2044;
        ELSIF x = 12506 THEN
            sigmoid_f := 2044;
        ELSIF x = 12507 THEN
            sigmoid_f := 2044;
        ELSIF x = 12508 THEN
            sigmoid_f := 2044;
        ELSIF x = 12509 THEN
            sigmoid_f := 2044;
        ELSIF x = 12510 THEN
            sigmoid_f := 2044;
        ELSIF x = 12511 THEN
            sigmoid_f := 2044;
        ELSIF x = 12512 THEN
            sigmoid_f := 2044;
        ELSIF x = 12513 THEN
            sigmoid_f := 2044;
        ELSIF x = 12514 THEN
            sigmoid_f := 2044;
        ELSIF x = 12515 THEN
            sigmoid_f := 2044;
        ELSIF x = 12516 THEN
            sigmoid_f := 2044;
        ELSIF x = 12517 THEN
            sigmoid_f := 2044;
        ELSIF x = 12518 THEN
            sigmoid_f := 2044;
        ELSIF x = 12519 THEN
            sigmoid_f := 2044;
        ELSIF x = 12520 THEN
            sigmoid_f := 2044;
        ELSIF x = 12521 THEN
            sigmoid_f := 2044;
        ELSIF x = 12522 THEN
            sigmoid_f := 2044;
        ELSIF x = 12523 THEN
            sigmoid_f := 2044;
        ELSIF x = 12524 THEN
            sigmoid_f := 2044;
        ELSIF x = 12525 THEN
            sigmoid_f := 2044;
        ELSIF x = 12526 THEN
            sigmoid_f := 2044;
        ELSIF x = 12527 THEN
            sigmoid_f := 2044;
        ELSIF x = 12528 THEN
            sigmoid_f := 2044;
        ELSIF x = 12529 THEN
            sigmoid_f := 2044;
        ELSIF x = 12530 THEN
            sigmoid_f := 2044;
        ELSIF x = 12531 THEN
            sigmoid_f := 2044;
        ELSIF x = 12532 THEN
            sigmoid_f := 2044;
        ELSIF x = 12533 THEN
            sigmoid_f := 2044;
        ELSIF x = 12534 THEN
            sigmoid_f := 2044;
        ELSIF x = 12535 THEN
            sigmoid_f := 2044;
        ELSIF x = 12536 THEN
            sigmoid_f := 2044;
        ELSIF x = 12537 THEN
            sigmoid_f := 2044;
        ELSIF x = 12538 THEN
            sigmoid_f := 2044;
        ELSIF x = 12539 THEN
            sigmoid_f := 2044;
        ELSIF x = 12540 THEN
            sigmoid_f := 2044;
        ELSIF x = 12541 THEN
            sigmoid_f := 2044;
        ELSIF x = 12542 THEN
            sigmoid_f := 2044;
        ELSIF x = 12543 THEN
            sigmoid_f := 2044;
        ELSIF x = 12544 THEN
            sigmoid_f := 2044;
        ELSIF x = 12545 THEN
            sigmoid_f := 2044;
        ELSIF x = 12546 THEN
            sigmoid_f := 2044;
        ELSIF x = 12547 THEN
            sigmoid_f := 2044;
        ELSIF x = 12548 THEN
            sigmoid_f := 2044;
        ELSIF x = 12549 THEN
            sigmoid_f := 2044;
        ELSIF x = 12550 THEN
            sigmoid_f := 2044;
        ELSIF x = 12551 THEN
            sigmoid_f := 2044;
        ELSIF x = 12552 THEN
            sigmoid_f := 2044;
        ELSIF x = 12553 THEN
            sigmoid_f := 2044;
        ELSIF x = 12554 THEN
            sigmoid_f := 2044;
        ELSIF x = 12555 THEN
            sigmoid_f := 2044;
        ELSIF x = 12556 THEN
            sigmoid_f := 2044;
        ELSIF x = 12557 THEN
            sigmoid_f := 2044;
        ELSIF x = 12558 THEN
            sigmoid_f := 2044;
        ELSIF x = 12559 THEN
            sigmoid_f := 2044;
        ELSIF x = 12560 THEN
            sigmoid_f := 2044;
        ELSIF x = 12561 THEN
            sigmoid_f := 2044;
        ELSIF x = 12562 THEN
            sigmoid_f := 2044;
        ELSIF x = 12563 THEN
            sigmoid_f := 2044;
        ELSIF x = 12564 THEN
            sigmoid_f := 2044;
        ELSIF x = 12565 THEN
            sigmoid_f := 2044;
        ELSIF x = 12566 THEN
            sigmoid_f := 2044;
        ELSIF x = 12567 THEN
            sigmoid_f := 2044;
        ELSIF x = 12568 THEN
            sigmoid_f := 2044;
        ELSIF x = 12569 THEN
            sigmoid_f := 2044;
        ELSIF x = 12570 THEN
            sigmoid_f := 2044;
        ELSIF x = 12571 THEN
            sigmoid_f := 2044;
        ELSIF x = 12572 THEN
            sigmoid_f := 2044;
        ELSIF x = 12573 THEN
            sigmoid_f := 2044;
        ELSIF x = 12574 THEN
            sigmoid_f := 2044;
        ELSIF x = 12575 THEN
            sigmoid_f := 2044;
        ELSIF x = 12576 THEN
            sigmoid_f := 2044;
        ELSIF x = 12577 THEN
            sigmoid_f := 2044;
        ELSIF x = 12578 THEN
            sigmoid_f := 2044;
        ELSIF x = 12579 THEN
            sigmoid_f := 2044;
        ELSIF x = 12580 THEN
            sigmoid_f := 2044;
        ELSIF x = 12581 THEN
            sigmoid_f := 2044;
        ELSIF x = 12582 THEN
            sigmoid_f := 2044;
        ELSIF x = 12583 THEN
            sigmoid_f := 2044;
        ELSIF x = 12584 THEN
            sigmoid_f := 2044;
        ELSIF x = 12585 THEN
            sigmoid_f := 2044;
        ELSIF x = 12586 THEN
            sigmoid_f := 2044;
        ELSIF x = 12587 THEN
            sigmoid_f := 2044;
        ELSIF x = 12588 THEN
            sigmoid_f := 2044;
        ELSIF x = 12589 THEN
            sigmoid_f := 2044;
        ELSIF x = 12590 THEN
            sigmoid_f := 2044;
        ELSIF x = 12591 THEN
            sigmoid_f := 2044;
        ELSIF x = 12592 THEN
            sigmoid_f := 2044;
        ELSIF x = 12593 THEN
            sigmoid_f := 2044;
        ELSIF x = 12594 THEN
            sigmoid_f := 2044;
        ELSIF x = 12595 THEN
            sigmoid_f := 2044;
        ELSIF x = 12596 THEN
            sigmoid_f := 2044;
        ELSIF x = 12597 THEN
            sigmoid_f := 2044;
        ELSIF x = 12598 THEN
            sigmoid_f := 2044;
        ELSIF x = 12599 THEN
            sigmoid_f := 2044;
        ELSIF x = 12600 THEN
            sigmoid_f := 2044;
        ELSIF x = 12601 THEN
            sigmoid_f := 2044;
        ELSIF x = 12602 THEN
            sigmoid_f := 2044;
        ELSIF x = 12603 THEN
            sigmoid_f := 2044;
        ELSIF x = 12604 THEN
            sigmoid_f := 2044;
        ELSIF x = 12605 THEN
            sigmoid_f := 2044;
        ELSIF x = 12606 THEN
            sigmoid_f := 2044;
        ELSIF x = 12607 THEN
            sigmoid_f := 2044;
        ELSIF x = 12608 THEN
            sigmoid_f := 2044;
        ELSIF x = 12609 THEN
            sigmoid_f := 2044;
        ELSIF x = 12610 THEN
            sigmoid_f := 2044;
        ELSIF x = 12611 THEN
            sigmoid_f := 2044;
        ELSIF x = 12612 THEN
            sigmoid_f := 2044;
        ELSIF x = 12613 THEN
            sigmoid_f := 2044;
        ELSIF x = 12614 THEN
            sigmoid_f := 2044;
        ELSIF x = 12615 THEN
            sigmoid_f := 2044;
        ELSIF x = 12616 THEN
            sigmoid_f := 2044;
        ELSIF x = 12617 THEN
            sigmoid_f := 2044;
        ELSIF x = 12618 THEN
            sigmoid_f := 2044;
        ELSIF x = 12619 THEN
            sigmoid_f := 2044;
        ELSIF x = 12620 THEN
            sigmoid_f := 2044;
        ELSIF x = 12621 THEN
            sigmoid_f := 2044;
        ELSIF x = 12622 THEN
            sigmoid_f := 2044;
        ELSIF x = 12623 THEN
            sigmoid_f := 2044;
        ELSIF x = 12624 THEN
            sigmoid_f := 2044;
        ELSIF x = 12625 THEN
            sigmoid_f := 2044;
        ELSIF x = 12626 THEN
            sigmoid_f := 2044;
        ELSIF x = 12627 THEN
            sigmoid_f := 2044;
        ELSIF x = 12628 THEN
            sigmoid_f := 2044;
        ELSIF x = 12629 THEN
            sigmoid_f := 2044;
        ELSIF x = 12630 THEN
            sigmoid_f := 2044;
        ELSIF x = 12631 THEN
            sigmoid_f := 2044;
        ELSIF x = 12632 THEN
            sigmoid_f := 2044;
        ELSIF x = 12633 THEN
            sigmoid_f := 2044;
        ELSIF x = 12634 THEN
            sigmoid_f := 2044;
        ELSIF x = 12635 THEN
            sigmoid_f := 2044;
        ELSIF x = 12636 THEN
            sigmoid_f := 2044;
        ELSIF x = 12637 THEN
            sigmoid_f := 2044;
        ELSIF x = 12638 THEN
            sigmoid_f := 2044;
        ELSIF x = 12639 THEN
            sigmoid_f := 2044;
        ELSIF x = 12640 THEN
            sigmoid_f := 2044;
        ELSIF x = 12641 THEN
            sigmoid_f := 2044;
        ELSIF x = 12642 THEN
            sigmoid_f := 2044;
        ELSIF x = 12643 THEN
            sigmoid_f := 2044;
        ELSIF x = 12644 THEN
            sigmoid_f := 2044;
        ELSIF x = 12645 THEN
            sigmoid_f := 2044;
        ELSIF x = 12646 THEN
            sigmoid_f := 2044;
        ELSIF x = 12647 THEN
            sigmoid_f := 2044;
        ELSIF x = 12648 THEN
            sigmoid_f := 2044;
        ELSIF x = 12649 THEN
            sigmoid_f := 2044;
        ELSIF x = 12650 THEN
            sigmoid_f := 2044;
        ELSIF x = 12651 THEN
            sigmoid_f := 2044;
        ELSIF x = 12652 THEN
            sigmoid_f := 2044;
        ELSIF x = 12653 THEN
            sigmoid_f := 2044;
        ELSIF x = 12654 THEN
            sigmoid_f := 2044;
        ELSIF x = 12655 THEN
            sigmoid_f := 2044;
        ELSIF x = 12656 THEN
            sigmoid_f := 2044;
        ELSIF x = 12657 THEN
            sigmoid_f := 2044;
        ELSIF x = 12658 THEN
            sigmoid_f := 2044;
        ELSIF x = 12659 THEN
            sigmoid_f := 2044;
        ELSIF x = 12660 THEN
            sigmoid_f := 2044;
        ELSIF x = 12661 THEN
            sigmoid_f := 2044;
        ELSIF x = 12662 THEN
            sigmoid_f := 2044;
        ELSIF x = 12663 THEN
            sigmoid_f := 2044;
        ELSIF x = 12664 THEN
            sigmoid_f := 2044;
        ELSIF x = 12665 THEN
            sigmoid_f := 2044;
        ELSIF x = 12666 THEN
            sigmoid_f := 2044;
        ELSIF x = 12667 THEN
            sigmoid_f := 2044;
        ELSIF x = 12668 THEN
            sigmoid_f := 2044;
        ELSIF x = 12669 THEN
            sigmoid_f := 2044;
        ELSIF x = 12670 THEN
            sigmoid_f := 2044;
        ELSIF x = 12671 THEN
            sigmoid_f := 2044;
        ELSIF x = 12672 THEN
            sigmoid_f := 2044;
        ELSIF x = 12673 THEN
            sigmoid_f := 2044;
        ELSIF x = 12674 THEN
            sigmoid_f := 2044;
        ELSIF x = 12675 THEN
            sigmoid_f := 2044;
        ELSIF x = 12676 THEN
            sigmoid_f := 2044;
        ELSIF x = 12677 THEN
            sigmoid_f := 2044;
        ELSIF x = 12678 THEN
            sigmoid_f := 2044;
        ELSIF x = 12679 THEN
            sigmoid_f := 2044;
        ELSIF x = 12680 THEN
            sigmoid_f := 2044;
        ELSIF x = 12681 THEN
            sigmoid_f := 2044;
        ELSIF x = 12682 THEN
            sigmoid_f := 2044;
        ELSIF x = 12683 THEN
            sigmoid_f := 2044;
        ELSIF x = 12684 THEN
            sigmoid_f := 2044;
        ELSIF x = 12685 THEN
            sigmoid_f := 2044;
        ELSIF x = 12686 THEN
            sigmoid_f := 2044;
        ELSIF x = 12687 THEN
            sigmoid_f := 2044;
        ELSIF x = 12688 THEN
            sigmoid_f := 2044;
        ELSIF x = 12689 THEN
            sigmoid_f := 2044;
        ELSIF x = 12690 THEN
            sigmoid_f := 2044;
        ELSIF x = 12691 THEN
            sigmoid_f := 2044;
        ELSIF x = 12692 THEN
            sigmoid_f := 2044;
        ELSIF x = 12693 THEN
            sigmoid_f := 2044;
        ELSIF x = 12694 THEN
            sigmoid_f := 2044;
        ELSIF x = 12695 THEN
            sigmoid_f := 2044;
        ELSIF x = 12696 THEN
            sigmoid_f := 2044;
        ELSIF x = 12697 THEN
            sigmoid_f := 2044;
        ELSIF x = 12698 THEN
            sigmoid_f := 2044;
        ELSIF x = 12699 THEN
            sigmoid_f := 2044;
        ELSIF x = 12700 THEN
            sigmoid_f := 2044;
        ELSIF x = 12701 THEN
            sigmoid_f := 2044;
        ELSIF x = 12702 THEN
            sigmoid_f := 2044;
        ELSIF x = 12703 THEN
            sigmoid_f := 2044;
        ELSIF x = 12704 THEN
            sigmoid_f := 2044;
        ELSIF x = 12705 THEN
            sigmoid_f := 2044;
        ELSIF x = 12706 THEN
            sigmoid_f := 2044;
        ELSIF x = 12707 THEN
            sigmoid_f := 2044;
        ELSIF x = 12708 THEN
            sigmoid_f := 2044;
        ELSIF x = 12709 THEN
            sigmoid_f := 2044;
        ELSIF x = 12710 THEN
            sigmoid_f := 2044;
        ELSIF x = 12711 THEN
            sigmoid_f := 2044;
        ELSIF x = 12712 THEN
            sigmoid_f := 2044;
        ELSIF x = 12713 THEN
            sigmoid_f := 2044;
        ELSIF x = 12714 THEN
            sigmoid_f := 2044;
        ELSIF x = 12715 THEN
            sigmoid_f := 2044;
        ELSIF x = 12716 THEN
            sigmoid_f := 2044;
        ELSIF x = 12717 THEN
            sigmoid_f := 2044;
        ELSIF x = 12718 THEN
            sigmoid_f := 2044;
        ELSIF x = 12719 THEN
            sigmoid_f := 2044;
        ELSIF x = 12720 THEN
            sigmoid_f := 2044;
        ELSIF x = 12721 THEN
            sigmoid_f := 2044;
        ELSIF x = 12722 THEN
            sigmoid_f := 2044;
        ELSIF x = 12723 THEN
            sigmoid_f := 2044;
        ELSIF x = 12724 THEN
            sigmoid_f := 2044;
        ELSIF x = 12725 THEN
            sigmoid_f := 2044;
        ELSIF x = 12726 THEN
            sigmoid_f := 2044;
        ELSIF x = 12727 THEN
            sigmoid_f := 2044;
        ELSIF x = 12728 THEN
            sigmoid_f := 2044;
        ELSIF x = 12729 THEN
            sigmoid_f := 2044;
        ELSIF x = 12730 THEN
            sigmoid_f := 2044;
        ELSIF x = 12731 THEN
            sigmoid_f := 2044;
        ELSIF x = 12732 THEN
            sigmoid_f := 2044;
        ELSIF x = 12733 THEN
            sigmoid_f := 2044;
        ELSIF x = 12734 THEN
            sigmoid_f := 2044;
        ELSIF x = 12735 THEN
            sigmoid_f := 2044;
        ELSIF x = 12736 THEN
            sigmoid_f := 2044;
        ELSIF x = 12737 THEN
            sigmoid_f := 2044;
        ELSIF x = 12738 THEN
            sigmoid_f := 2044;
        ELSIF x = 12739 THEN
            sigmoid_f := 2044;
        ELSIF x = 12740 THEN
            sigmoid_f := 2044;
        ELSIF x = 12741 THEN
            sigmoid_f := 2044;
        ELSIF x = 12742 THEN
            sigmoid_f := 2044;
        ELSIF x = 12743 THEN
            sigmoid_f := 2044;
        ELSIF x = 12744 THEN
            sigmoid_f := 2044;
        ELSIF x = 12745 THEN
            sigmoid_f := 2044;
        ELSIF x = 12746 THEN
            sigmoid_f := 2044;
        ELSIF x = 12747 THEN
            sigmoid_f := 2044;
        ELSIF x = 12748 THEN
            sigmoid_f := 2044;
        ELSIF x = 12749 THEN
            sigmoid_f := 2044;
        ELSIF x = 12750 THEN
            sigmoid_f := 2044;
        ELSIF x = 12751 THEN
            sigmoid_f := 2044;
        ELSIF x = 12752 THEN
            sigmoid_f := 2044;
        ELSIF x = 12753 THEN
            sigmoid_f := 2044;
        ELSIF x = 12754 THEN
            sigmoid_f := 2044;
        ELSIF x = 12755 THEN
            sigmoid_f := 2044;
        ELSIF x = 12756 THEN
            sigmoid_f := 2044;
        ELSIF x = 12757 THEN
            sigmoid_f := 2044;
        ELSIF x = 12758 THEN
            sigmoid_f := 2044;
        ELSIF x = 12759 THEN
            sigmoid_f := 2044;
        ELSIF x = 12760 THEN
            sigmoid_f := 2044;
        ELSIF x = 12761 THEN
            sigmoid_f := 2044;
        ELSIF x = 12762 THEN
            sigmoid_f := 2044;
        ELSIF x = 12763 THEN
            sigmoid_f := 2044;
        ELSIF x = 12764 THEN
            sigmoid_f := 2044;
        ELSIF x = 12765 THEN
            sigmoid_f := 2044;
        ELSIF x = 12766 THEN
            sigmoid_f := 2044;
        ELSIF x = 12767 THEN
            sigmoid_f := 2044;
        ELSIF x = 12768 THEN
            sigmoid_f := 2044;
        ELSIF x = 12769 THEN
            sigmoid_f := 2044;
        ELSIF x = 12770 THEN
            sigmoid_f := 2044;
        ELSIF x = 12771 THEN
            sigmoid_f := 2044;
        ELSIF x = 12772 THEN
            sigmoid_f := 2044;
        ELSIF x = 12773 THEN
            sigmoid_f := 2044;
        ELSIF x = 12774 THEN
            sigmoid_f := 2044;
        ELSIF x = 12775 THEN
            sigmoid_f := 2044;
        ELSIF x = 12776 THEN
            sigmoid_f := 2044;
        ELSIF x = 12777 THEN
            sigmoid_f := 2044;
        ELSIF x = 12778 THEN
            sigmoid_f := 2044;
        ELSIF x = 12779 THEN
            sigmoid_f := 2044;
        ELSIF x = 12780 THEN
            sigmoid_f := 2044;
        ELSIF x = 12781 THEN
            sigmoid_f := 2044;
        ELSIF x = 12782 THEN
            sigmoid_f := 2044;
        ELSIF x = 12783 THEN
            sigmoid_f := 2044;
        ELSIF x = 12784 THEN
            sigmoid_f := 2044;
        ELSIF x = 12785 THEN
            sigmoid_f := 2044;
        ELSIF x = 12786 THEN
            sigmoid_f := 2044;
        ELSIF x = 12787 THEN
            sigmoid_f := 2044;
        ELSIF x = 12788 THEN
            sigmoid_f := 2044;
        ELSIF x = 12789 THEN
            sigmoid_f := 2044;
        ELSIF x = 12790 THEN
            sigmoid_f := 2044;
        ELSIF x = 12791 THEN
            sigmoid_f := 2044;
        ELSIF x = 12792 THEN
            sigmoid_f := 2044;
        ELSIF x = 12793 THEN
            sigmoid_f := 2044;
        ELSIF x = 12794 THEN
            sigmoid_f := 2044;
        ELSIF x = 12795 THEN
            sigmoid_f := 2044;
        ELSIF x = 12796 THEN
            sigmoid_f := 2044;
        ELSIF x = 12797 THEN
            sigmoid_f := 2044;
        ELSIF x = 12798 THEN
            sigmoid_f := 2044;
        ELSIF x = 12799 THEN
            sigmoid_f := 2044;
        ELSIF x = 12800 THEN
            sigmoid_f := 2045;
        ELSIF x = 12801 THEN
            sigmoid_f := 2045;
        ELSIF x = 12802 THEN
            sigmoid_f := 2045;
        ELSIF x = 12803 THEN
            sigmoid_f := 2045;
        ELSIF x = 12804 THEN
            sigmoid_f := 2045;
        ELSIF x = 12805 THEN
            sigmoid_f := 2045;
        ELSIF x = 12806 THEN
            sigmoid_f := 2045;
        ELSIF x = 12807 THEN
            sigmoid_f := 2045;
        ELSIF x = 12808 THEN
            sigmoid_f := 2045;
        ELSIF x = 12809 THEN
            sigmoid_f := 2045;
        ELSIF x = 12810 THEN
            sigmoid_f := 2045;
        ELSIF x = 12811 THEN
            sigmoid_f := 2045;
        ELSIF x = 12812 THEN
            sigmoid_f := 2045;
        ELSIF x = 12813 THEN
            sigmoid_f := 2045;
        ELSIF x = 12814 THEN
            sigmoid_f := 2045;
        ELSIF x = 12815 THEN
            sigmoid_f := 2045;
        ELSIF x = 12816 THEN
            sigmoid_f := 2045;
        ELSIF x = 12817 THEN
            sigmoid_f := 2045;
        ELSIF x = 12818 THEN
            sigmoid_f := 2045;
        ELSIF x = 12819 THEN
            sigmoid_f := 2045;
        ELSIF x = 12820 THEN
            sigmoid_f := 2045;
        ELSIF x = 12821 THEN
            sigmoid_f := 2045;
        ELSIF x = 12822 THEN
            sigmoid_f := 2045;
        ELSIF x = 12823 THEN
            sigmoid_f := 2045;
        ELSIF x = 12824 THEN
            sigmoid_f := 2045;
        ELSIF x = 12825 THEN
            sigmoid_f := 2045;
        ELSIF x = 12826 THEN
            sigmoid_f := 2045;
        ELSIF x = 12827 THEN
            sigmoid_f := 2045;
        ELSIF x = 12828 THEN
            sigmoid_f := 2045;
        ELSIF x = 12829 THEN
            sigmoid_f := 2045;
        ELSIF x = 12830 THEN
            sigmoid_f := 2045;
        ELSIF x = 12831 THEN
            sigmoid_f := 2045;
        ELSIF x = 12832 THEN
            sigmoid_f := 2045;
        ELSIF x = 12833 THEN
            sigmoid_f := 2045;
        ELSIF x = 12834 THEN
            sigmoid_f := 2045;
        ELSIF x = 12835 THEN
            sigmoid_f := 2045;
        ELSIF x = 12836 THEN
            sigmoid_f := 2045;
        ELSIF x = 12837 THEN
            sigmoid_f := 2045;
        ELSIF x = 12838 THEN
            sigmoid_f := 2045;
        ELSIF x = 12839 THEN
            sigmoid_f := 2045;
        ELSIF x = 12840 THEN
            sigmoid_f := 2045;
        ELSIF x = 12841 THEN
            sigmoid_f := 2045;
        ELSIF x = 12842 THEN
            sigmoid_f := 2045;
        ELSIF x = 12843 THEN
            sigmoid_f := 2045;
        ELSIF x = 12844 THEN
            sigmoid_f := 2045;
        ELSIF x = 12845 THEN
            sigmoid_f := 2045;
        ELSIF x = 12846 THEN
            sigmoid_f := 2045;
        ELSIF x = 12847 THEN
            sigmoid_f := 2045;
        ELSIF x = 12848 THEN
            sigmoid_f := 2045;
        ELSIF x = 12849 THEN
            sigmoid_f := 2045;
        ELSIF x = 12850 THEN
            sigmoid_f := 2045;
        ELSIF x = 12851 THEN
            sigmoid_f := 2045;
        ELSIF x = 12852 THEN
            sigmoid_f := 2045;
        ELSIF x = 12853 THEN
            sigmoid_f := 2045;
        ELSIF x = 12854 THEN
            sigmoid_f := 2045;
        ELSIF x = 12855 THEN
            sigmoid_f := 2045;
        ELSIF x = 12856 THEN
            sigmoid_f := 2045;
        ELSIF x = 12857 THEN
            sigmoid_f := 2045;
        ELSIF x = 12858 THEN
            sigmoid_f := 2045;
        ELSIF x = 12859 THEN
            sigmoid_f := 2045;
        ELSIF x = 12860 THEN
            sigmoid_f := 2045;
        ELSIF x = 12861 THEN
            sigmoid_f := 2045;
        ELSIF x = 12862 THEN
            sigmoid_f := 2045;
        ELSIF x = 12863 THEN
            sigmoid_f := 2045;
        ELSIF x = 12864 THEN
            sigmoid_f := 2045;
        ELSIF x = 12865 THEN
            sigmoid_f := 2045;
        ELSIF x = 12866 THEN
            sigmoid_f := 2045;
        ELSIF x = 12867 THEN
            sigmoid_f := 2045;
        ELSIF x = 12868 THEN
            sigmoid_f := 2045;
        ELSIF x = 12869 THEN
            sigmoid_f := 2045;
        ELSIF x = 12870 THEN
            sigmoid_f := 2045;
        ELSIF x = 12871 THEN
            sigmoid_f := 2045;
        ELSIF x = 12872 THEN
            sigmoid_f := 2045;
        ELSIF x = 12873 THEN
            sigmoid_f := 2045;
        ELSIF x = 12874 THEN
            sigmoid_f := 2045;
        ELSIF x = 12875 THEN
            sigmoid_f := 2045;
        ELSIF x = 12876 THEN
            sigmoid_f := 2045;
        ELSIF x = 12877 THEN
            sigmoid_f := 2045;
        ELSIF x = 12878 THEN
            sigmoid_f := 2045;
        ELSIF x = 12879 THEN
            sigmoid_f := 2045;
        ELSIF x = 12880 THEN
            sigmoid_f := 2045;
        ELSIF x = 12881 THEN
            sigmoid_f := 2045;
        ELSIF x = 12882 THEN
            sigmoid_f := 2045;
        ELSIF x = 12883 THEN
            sigmoid_f := 2045;
        ELSIF x = 12884 THEN
            sigmoid_f := 2045;
        ELSIF x = 12885 THEN
            sigmoid_f := 2045;
        ELSIF x = 12886 THEN
            sigmoid_f := 2045;
        ELSIF x = 12887 THEN
            sigmoid_f := 2045;
        ELSIF x = 12888 THEN
            sigmoid_f := 2045;
        ELSIF x = 12889 THEN
            sigmoid_f := 2045;
        ELSIF x = 12890 THEN
            sigmoid_f := 2045;
        ELSIF x = 12891 THEN
            sigmoid_f := 2045;
        ELSIF x = 12892 THEN
            sigmoid_f := 2045;
        ELSIF x = 12893 THEN
            sigmoid_f := 2045;
        ELSIF x = 12894 THEN
            sigmoid_f := 2045;
        ELSIF x = 12895 THEN
            sigmoid_f := 2045;
        ELSIF x = 12896 THEN
            sigmoid_f := 2045;
        ELSIF x = 12897 THEN
            sigmoid_f := 2045;
        ELSIF x = 12898 THEN
            sigmoid_f := 2045;
        ELSIF x = 12899 THEN
            sigmoid_f := 2045;
        ELSIF x = 12900 THEN
            sigmoid_f := 2045;
        ELSIF x = 12901 THEN
            sigmoid_f := 2045;
        ELSIF x = 12902 THEN
            sigmoid_f := 2045;
        ELSIF x = 12903 THEN
            sigmoid_f := 2045;
        ELSIF x = 12904 THEN
            sigmoid_f := 2045;
        ELSIF x = 12905 THEN
            sigmoid_f := 2045;
        ELSIF x = 12906 THEN
            sigmoid_f := 2045;
        ELSIF x = 12907 THEN
            sigmoid_f := 2045;
        ELSIF x = 12908 THEN
            sigmoid_f := 2045;
        ELSIF x = 12909 THEN
            sigmoid_f := 2045;
        ELSIF x = 12910 THEN
            sigmoid_f := 2045;
        ELSIF x = 12911 THEN
            sigmoid_f := 2045;
        ELSIF x = 12912 THEN
            sigmoid_f := 2045;
        ELSIF x = 12913 THEN
            sigmoid_f := 2045;
        ELSIF x = 12914 THEN
            sigmoid_f := 2045;
        ELSIF x = 12915 THEN
            sigmoid_f := 2045;
        ELSIF x = 12916 THEN
            sigmoid_f := 2045;
        ELSIF x = 12917 THEN
            sigmoid_f := 2045;
        ELSIF x = 12918 THEN
            sigmoid_f := 2045;
        ELSIF x = 12919 THEN
            sigmoid_f := 2045;
        ELSIF x = 12920 THEN
            sigmoid_f := 2045;
        ELSIF x = 12921 THEN
            sigmoid_f := 2045;
        ELSIF x = 12922 THEN
            sigmoid_f := 2045;
        ELSIF x = 12923 THEN
            sigmoid_f := 2045;
        ELSIF x = 12924 THEN
            sigmoid_f := 2045;
        ELSIF x = 12925 THEN
            sigmoid_f := 2045;
        ELSIF x = 12926 THEN
            sigmoid_f := 2045;
        ELSIF x = 12927 THEN
            sigmoid_f := 2045;
        ELSIF x = 12928 THEN
            sigmoid_f := 2045;
        ELSIF x = 12929 THEN
            sigmoid_f := 2045;
        ELSIF x = 12930 THEN
            sigmoid_f := 2045;
        ELSIF x = 12931 THEN
            sigmoid_f := 2045;
        ELSIF x = 12932 THEN
            sigmoid_f := 2045;
        ELSIF x = 12933 THEN
            sigmoid_f := 2045;
        ELSIF x = 12934 THEN
            sigmoid_f := 2045;
        ELSIF x = 12935 THEN
            sigmoid_f := 2045;
        ELSIF x = 12936 THEN
            sigmoid_f := 2045;
        ELSIF x = 12937 THEN
            sigmoid_f := 2045;
        ELSIF x = 12938 THEN
            sigmoid_f := 2045;
        ELSIF x = 12939 THEN
            sigmoid_f := 2045;
        ELSIF x = 12940 THEN
            sigmoid_f := 2045;
        ELSIF x = 12941 THEN
            sigmoid_f := 2045;
        ELSIF x = 12942 THEN
            sigmoid_f := 2045;
        ELSIF x = 12943 THEN
            sigmoid_f := 2045;
        ELSIF x = 12944 THEN
            sigmoid_f := 2045;
        ELSIF x = 12945 THEN
            sigmoid_f := 2045;
        ELSIF x = 12946 THEN
            sigmoid_f := 2045;
        ELSIF x = 12947 THEN
            sigmoid_f := 2045;
        ELSIF x = 12948 THEN
            sigmoid_f := 2045;
        ELSIF x = 12949 THEN
            sigmoid_f := 2045;
        ELSIF x = 12950 THEN
            sigmoid_f := 2045;
        ELSIF x = 12951 THEN
            sigmoid_f := 2045;
        ELSIF x = 12952 THEN
            sigmoid_f := 2045;
        ELSIF x = 12953 THEN
            sigmoid_f := 2045;
        ELSIF x = 12954 THEN
            sigmoid_f := 2045;
        ELSIF x = 12955 THEN
            sigmoid_f := 2045;
        ELSIF x = 12956 THEN
            sigmoid_f := 2045;
        ELSIF x = 12957 THEN
            sigmoid_f := 2045;
        ELSIF x = 12958 THEN
            sigmoid_f := 2045;
        ELSIF x = 12959 THEN
            sigmoid_f := 2045;
        ELSIF x = 12960 THEN
            sigmoid_f := 2045;
        ELSIF x = 12961 THEN
            sigmoid_f := 2045;
        ELSIF x = 12962 THEN
            sigmoid_f := 2045;
        ELSIF x = 12963 THEN
            sigmoid_f := 2045;
        ELSIF x = 12964 THEN
            sigmoid_f := 2045;
        ELSIF x = 12965 THEN
            sigmoid_f := 2045;
        ELSIF x = 12966 THEN
            sigmoid_f := 2045;
        ELSIF x = 12967 THEN
            sigmoid_f := 2045;
        ELSIF x = 12968 THEN
            sigmoid_f := 2045;
        ELSIF x = 12969 THEN
            sigmoid_f := 2045;
        ELSIF x = 12970 THEN
            sigmoid_f := 2045;
        ELSIF x = 12971 THEN
            sigmoid_f := 2045;
        ELSIF x = 12972 THEN
            sigmoid_f := 2045;
        ELSIF x = 12973 THEN
            sigmoid_f := 2045;
        ELSIF x = 12974 THEN
            sigmoid_f := 2045;
        ELSIF x = 12975 THEN
            sigmoid_f := 2045;
        ELSIF x = 12976 THEN
            sigmoid_f := 2045;
        ELSIF x = 12977 THEN
            sigmoid_f := 2045;
        ELSIF x = 12978 THEN
            sigmoid_f := 2045;
        ELSIF x = 12979 THEN
            sigmoid_f := 2045;
        ELSIF x = 12980 THEN
            sigmoid_f := 2045;
        ELSIF x = 12981 THEN
            sigmoid_f := 2045;
        ELSIF x = 12982 THEN
            sigmoid_f := 2045;
        ELSIF x = 12983 THEN
            sigmoid_f := 2045;
        ELSIF x = 12984 THEN
            sigmoid_f := 2045;
        ELSIF x = 12985 THEN
            sigmoid_f := 2045;
        ELSIF x = 12986 THEN
            sigmoid_f := 2045;
        ELSIF x = 12987 THEN
            sigmoid_f := 2045;
        ELSIF x = 12988 THEN
            sigmoid_f := 2045;
        ELSIF x = 12989 THEN
            sigmoid_f := 2045;
        ELSIF x = 12990 THEN
            sigmoid_f := 2045;
        ELSIF x = 12991 THEN
            sigmoid_f := 2045;
        ELSIF x = 12992 THEN
            sigmoid_f := 2045;
        ELSIF x = 12993 THEN
            sigmoid_f := 2045;
        ELSIF x = 12994 THEN
            sigmoid_f := 2045;
        ELSIF x = 12995 THEN
            sigmoid_f := 2045;
        ELSIF x = 12996 THEN
            sigmoid_f := 2045;
        ELSIF x = 12997 THEN
            sigmoid_f := 2045;
        ELSIF x = 12998 THEN
            sigmoid_f := 2045;
        ELSIF x = 12999 THEN
            sigmoid_f := 2045;
        ELSIF x = 13000 THEN
            sigmoid_f := 2045;
        ELSIF x = 13001 THEN
            sigmoid_f := 2045;
        ELSIF x = 13002 THEN
            sigmoid_f := 2045;
        ELSIF x = 13003 THEN
            sigmoid_f := 2045;
        ELSIF x = 13004 THEN
            sigmoid_f := 2045;
        ELSIF x = 13005 THEN
            sigmoid_f := 2045;
        ELSIF x = 13006 THEN
            sigmoid_f := 2045;
        ELSIF x = 13007 THEN
            sigmoid_f := 2045;
        ELSIF x = 13008 THEN
            sigmoid_f := 2045;
        ELSIF x = 13009 THEN
            sigmoid_f := 2045;
        ELSIF x = 13010 THEN
            sigmoid_f := 2045;
        ELSIF x = 13011 THEN
            sigmoid_f := 2045;
        ELSIF x = 13012 THEN
            sigmoid_f := 2045;
        ELSIF x = 13013 THEN
            sigmoid_f := 2045;
        ELSIF x = 13014 THEN
            sigmoid_f := 2045;
        ELSIF x = 13015 THEN
            sigmoid_f := 2045;
        ELSIF x = 13016 THEN
            sigmoid_f := 2045;
        ELSIF x = 13017 THEN
            sigmoid_f := 2045;
        ELSIF x = 13018 THEN
            sigmoid_f := 2045;
        ELSIF x = 13019 THEN
            sigmoid_f := 2045;
        ELSIF x = 13020 THEN
            sigmoid_f := 2045;
        ELSIF x = 13021 THEN
            sigmoid_f := 2045;
        ELSIF x = 13022 THEN
            sigmoid_f := 2045;
        ELSIF x = 13023 THEN
            sigmoid_f := 2045;
        ELSIF x = 13024 THEN
            sigmoid_f := 2045;
        ELSIF x = 13025 THEN
            sigmoid_f := 2045;
        ELSIF x = 13026 THEN
            sigmoid_f := 2045;
        ELSIF x = 13027 THEN
            sigmoid_f := 2045;
        ELSIF x = 13028 THEN
            sigmoid_f := 2045;
        ELSIF x = 13029 THEN
            sigmoid_f := 2045;
        ELSIF x = 13030 THEN
            sigmoid_f := 2045;
        ELSIF x = 13031 THEN
            sigmoid_f := 2045;
        ELSIF x = 13032 THEN
            sigmoid_f := 2045;
        ELSIF x = 13033 THEN
            sigmoid_f := 2045;
        ELSIF x = 13034 THEN
            sigmoid_f := 2045;
        ELSIF x = 13035 THEN
            sigmoid_f := 2045;
        ELSIF x = 13036 THEN
            sigmoid_f := 2045;
        ELSIF x = 13037 THEN
            sigmoid_f := 2045;
        ELSIF x = 13038 THEN
            sigmoid_f := 2045;
        ELSIF x = 13039 THEN
            sigmoid_f := 2045;
        ELSIF x = 13040 THEN
            sigmoid_f := 2045;
        ELSIF x = 13041 THEN
            sigmoid_f := 2045;
        ELSIF x = 13042 THEN
            sigmoid_f := 2045;
        ELSIF x = 13043 THEN
            sigmoid_f := 2045;
        ELSIF x = 13044 THEN
            sigmoid_f := 2045;
        ELSIF x = 13045 THEN
            sigmoid_f := 2045;
        ELSIF x = 13046 THEN
            sigmoid_f := 2045;
        ELSIF x = 13047 THEN
            sigmoid_f := 2045;
        ELSIF x = 13048 THEN
            sigmoid_f := 2045;
        ELSIF x = 13049 THEN
            sigmoid_f := 2045;
        ELSIF x = 13050 THEN
            sigmoid_f := 2045;
        ELSIF x = 13051 THEN
            sigmoid_f := 2045;
        ELSIF x = 13052 THEN
            sigmoid_f := 2045;
        ELSIF x = 13053 THEN
            sigmoid_f := 2045;
        ELSIF x = 13054 THEN
            sigmoid_f := 2045;
        ELSIF x = 13055 THEN
            sigmoid_f := 2045;
        ELSIF x = 13056 THEN
            sigmoid_f := 2045;
        ELSIF x = 13057 THEN
            sigmoid_f := 2045;
        ELSIF x = 13058 THEN
            sigmoid_f := 2045;
        ELSIF x = 13059 THEN
            sigmoid_f := 2045;
        ELSIF x = 13060 THEN
            sigmoid_f := 2045;
        ELSIF x = 13061 THEN
            sigmoid_f := 2045;
        ELSIF x = 13062 THEN
            sigmoid_f := 2045;
        ELSIF x = 13063 THEN
            sigmoid_f := 2045;
        ELSIF x = 13064 THEN
            sigmoid_f := 2045;
        ELSIF x = 13065 THEN
            sigmoid_f := 2045;
        ELSIF x = 13066 THEN
            sigmoid_f := 2045;
        ELSIF x = 13067 THEN
            sigmoid_f := 2045;
        ELSIF x = 13068 THEN
            sigmoid_f := 2045;
        ELSIF x = 13069 THEN
            sigmoid_f := 2045;
        ELSIF x = 13070 THEN
            sigmoid_f := 2045;
        ELSIF x = 13071 THEN
            sigmoid_f := 2045;
        ELSIF x = 13072 THEN
            sigmoid_f := 2045;
        ELSIF x = 13073 THEN
            sigmoid_f := 2045;
        ELSIF x = 13074 THEN
            sigmoid_f := 2045;
        ELSIF x = 13075 THEN
            sigmoid_f := 2045;
        ELSIF x = 13076 THEN
            sigmoid_f := 2045;
        ELSIF x = 13077 THEN
            sigmoid_f := 2045;
        ELSIF x = 13078 THEN
            sigmoid_f := 2045;
        ELSIF x = 13079 THEN
            sigmoid_f := 2045;
        ELSIF x = 13080 THEN
            sigmoid_f := 2045;
        ELSIF x = 13081 THEN
            sigmoid_f := 2045;
        ELSIF x = 13082 THEN
            sigmoid_f := 2045;
        ELSIF x = 13083 THEN
            sigmoid_f := 2045;
        ELSIF x = 13084 THEN
            sigmoid_f := 2045;
        ELSIF x = 13085 THEN
            sigmoid_f := 2045;
        ELSIF x = 13086 THEN
            sigmoid_f := 2045;
        ELSIF x = 13087 THEN
            sigmoid_f := 2045;
        ELSIF x = 13088 THEN
            sigmoid_f := 2045;
        ELSIF x = 13089 THEN
            sigmoid_f := 2045;
        ELSIF x = 13090 THEN
            sigmoid_f := 2045;
        ELSIF x = 13091 THEN
            sigmoid_f := 2045;
        ELSIF x = 13092 THEN
            sigmoid_f := 2045;
        ELSIF x = 13093 THEN
            sigmoid_f := 2045;
        ELSIF x = 13094 THEN
            sigmoid_f := 2045;
        ELSIF x = 13095 THEN
            sigmoid_f := 2045;
        ELSIF x = 13096 THEN
            sigmoid_f := 2045;
        ELSIF x = 13097 THEN
            sigmoid_f := 2045;
        ELSIF x = 13098 THEN
            sigmoid_f := 2045;
        ELSIF x = 13099 THEN
            sigmoid_f := 2045;
        ELSIF x = 13100 THEN
            sigmoid_f := 2045;
        ELSIF x = 13101 THEN
            sigmoid_f := 2045;
        ELSIF x = 13102 THEN
            sigmoid_f := 2045;
        ELSIF x = 13103 THEN
            sigmoid_f := 2045;
        ELSIF x = 13104 THEN
            sigmoid_f := 2045;
        ELSIF x = 13105 THEN
            sigmoid_f := 2045;
        ELSIF x = 13106 THEN
            sigmoid_f := 2045;
        ELSIF x = 13107 THEN
            sigmoid_f := 2045;
        ELSIF x = 13108 THEN
            sigmoid_f := 2045;
        ELSIF x = 13109 THEN
            sigmoid_f := 2045;
        ELSIF x = 13110 THEN
            sigmoid_f := 2045;
        ELSIF x = 13111 THEN
            sigmoid_f := 2045;
        ELSIF x = 13112 THEN
            sigmoid_f := 2045;
        ELSIF x = 13113 THEN
            sigmoid_f := 2045;
        ELSIF x = 13114 THEN
            sigmoid_f := 2045;
        ELSIF x = 13115 THEN
            sigmoid_f := 2045;
        ELSIF x = 13116 THEN
            sigmoid_f := 2045;
        ELSIF x = 13117 THEN
            sigmoid_f := 2045;
        ELSIF x = 13118 THEN
            sigmoid_f := 2045;
        ELSIF x = 13119 THEN
            sigmoid_f := 2045;
        ELSIF x = 13120 THEN
            sigmoid_f := 2045;
        ELSIF x = 13121 THEN
            sigmoid_f := 2045;
        ELSIF x = 13122 THEN
            sigmoid_f := 2045;
        ELSIF x = 13123 THEN
            sigmoid_f := 2045;
        ELSIF x = 13124 THEN
            sigmoid_f := 2045;
        ELSIF x = 13125 THEN
            sigmoid_f := 2045;
        ELSIF x = 13126 THEN
            sigmoid_f := 2045;
        ELSIF x = 13127 THEN
            sigmoid_f := 2045;
        ELSIF x = 13128 THEN
            sigmoid_f := 2045;
        ELSIF x = 13129 THEN
            sigmoid_f := 2045;
        ELSIF x = 13130 THEN
            sigmoid_f := 2045;
        ELSIF x = 13131 THEN
            sigmoid_f := 2045;
        ELSIF x = 13132 THEN
            sigmoid_f := 2045;
        ELSIF x = 13133 THEN
            sigmoid_f := 2045;
        ELSIF x = 13134 THEN
            sigmoid_f := 2045;
        ELSIF x = 13135 THEN
            sigmoid_f := 2045;
        ELSIF x = 13136 THEN
            sigmoid_f := 2045;
        ELSIF x = 13137 THEN
            sigmoid_f := 2045;
        ELSIF x = 13138 THEN
            sigmoid_f := 2045;
        ELSIF x = 13139 THEN
            sigmoid_f := 2045;
        ELSIF x = 13140 THEN
            sigmoid_f := 2045;
        ELSIF x = 13141 THEN
            sigmoid_f := 2045;
        ELSIF x = 13142 THEN
            sigmoid_f := 2045;
        ELSIF x = 13143 THEN
            sigmoid_f := 2045;
        ELSIF x = 13144 THEN
            sigmoid_f := 2045;
        ELSIF x = 13145 THEN
            sigmoid_f := 2045;
        ELSIF x = 13146 THEN
            sigmoid_f := 2045;
        ELSIF x = 13147 THEN
            sigmoid_f := 2045;
        ELSIF x = 13148 THEN
            sigmoid_f := 2045;
        ELSIF x = 13149 THEN
            sigmoid_f := 2045;
        ELSIF x = 13150 THEN
            sigmoid_f := 2045;
        ELSIF x = 13151 THEN
            sigmoid_f := 2045;
        ELSIF x = 13152 THEN
            sigmoid_f := 2045;
        ELSIF x = 13153 THEN
            sigmoid_f := 2045;
        ELSIF x = 13154 THEN
            sigmoid_f := 2045;
        ELSIF x = 13155 THEN
            sigmoid_f := 2045;
        ELSIF x = 13156 THEN
            sigmoid_f := 2045;
        ELSIF x = 13157 THEN
            sigmoid_f := 2045;
        ELSIF x = 13158 THEN
            sigmoid_f := 2045;
        ELSIF x = 13159 THEN
            sigmoid_f := 2045;
        ELSIF x = 13160 THEN
            sigmoid_f := 2045;
        ELSIF x = 13161 THEN
            sigmoid_f := 2045;
        ELSIF x = 13162 THEN
            sigmoid_f := 2045;
        ELSIF x = 13163 THEN
            sigmoid_f := 2045;
        ELSIF x = 13164 THEN
            sigmoid_f := 2045;
        ELSIF x = 13165 THEN
            sigmoid_f := 2045;
        ELSIF x = 13166 THEN
            sigmoid_f := 2045;
        ELSIF x = 13167 THEN
            sigmoid_f := 2045;
        ELSIF x = 13168 THEN
            sigmoid_f := 2045;
        ELSIF x = 13169 THEN
            sigmoid_f := 2045;
        ELSIF x = 13170 THEN
            sigmoid_f := 2045;
        ELSIF x = 13171 THEN
            sigmoid_f := 2045;
        ELSIF x = 13172 THEN
            sigmoid_f := 2045;
        ELSIF x = 13173 THEN
            sigmoid_f := 2045;
        ELSIF x = 13174 THEN
            sigmoid_f := 2045;
        ELSIF x = 13175 THEN
            sigmoid_f := 2045;
        ELSIF x = 13176 THEN
            sigmoid_f := 2045;
        ELSIF x = 13177 THEN
            sigmoid_f := 2045;
        ELSIF x = 13178 THEN
            sigmoid_f := 2045;
        ELSIF x = 13179 THEN
            sigmoid_f := 2045;
        ELSIF x = 13180 THEN
            sigmoid_f := 2045;
        ELSIF x = 13181 THEN
            sigmoid_f := 2045;
        ELSIF x = 13182 THEN
            sigmoid_f := 2045;
        ELSIF x = 13183 THEN
            sigmoid_f := 2045;
        ELSIF x = 13184 THEN
            sigmoid_f := 2045;
        ELSIF x = 13185 THEN
            sigmoid_f := 2045;
        ELSIF x = 13186 THEN
            sigmoid_f := 2045;
        ELSIF x = 13187 THEN
            sigmoid_f := 2045;
        ELSIF x = 13188 THEN
            sigmoid_f := 2045;
        ELSIF x = 13189 THEN
            sigmoid_f := 2045;
        ELSIF x = 13190 THEN
            sigmoid_f := 2045;
        ELSIF x = 13191 THEN
            sigmoid_f := 2045;
        ELSIF x = 13192 THEN
            sigmoid_f := 2045;
        ELSIF x = 13193 THEN
            sigmoid_f := 2045;
        ELSIF x = 13194 THEN
            sigmoid_f := 2045;
        ELSIF x = 13195 THEN
            sigmoid_f := 2045;
        ELSIF x = 13196 THEN
            sigmoid_f := 2045;
        ELSIF x = 13197 THEN
            sigmoid_f := 2045;
        ELSIF x = 13198 THEN
            sigmoid_f := 2045;
        ELSIF x = 13199 THEN
            sigmoid_f := 2045;
        ELSIF x = 13200 THEN
            sigmoid_f := 2045;
        ELSIF x = 13201 THEN
            sigmoid_f := 2045;
        ELSIF x = 13202 THEN
            sigmoid_f := 2045;
        ELSIF x = 13203 THEN
            sigmoid_f := 2045;
        ELSIF x = 13204 THEN
            sigmoid_f := 2045;
        ELSIF x = 13205 THEN
            sigmoid_f := 2045;
        ELSIF x = 13206 THEN
            sigmoid_f := 2045;
        ELSIF x = 13207 THEN
            sigmoid_f := 2045;
        ELSIF x = 13208 THEN
            sigmoid_f := 2045;
        ELSIF x = 13209 THEN
            sigmoid_f := 2045;
        ELSIF x = 13210 THEN
            sigmoid_f := 2045;
        ELSIF x = 13211 THEN
            sigmoid_f := 2045;
        ELSIF x = 13212 THEN
            sigmoid_f := 2045;
        ELSIF x = 13213 THEN
            sigmoid_f := 2045;
        ELSIF x = 13214 THEN
            sigmoid_f := 2045;
        ELSIF x = 13215 THEN
            sigmoid_f := 2045;
        ELSIF x = 13216 THEN
            sigmoid_f := 2045;
        ELSIF x = 13217 THEN
            sigmoid_f := 2045;
        ELSIF x = 13218 THEN
            sigmoid_f := 2045;
        ELSIF x = 13219 THEN
            sigmoid_f := 2045;
        ELSIF x = 13220 THEN
            sigmoid_f := 2045;
        ELSIF x = 13221 THEN
            sigmoid_f := 2045;
        ELSIF x = 13222 THEN
            sigmoid_f := 2045;
        ELSIF x = 13223 THEN
            sigmoid_f := 2045;
        ELSIF x = 13224 THEN
            sigmoid_f := 2045;
        ELSIF x = 13225 THEN
            sigmoid_f := 2045;
        ELSIF x = 13226 THEN
            sigmoid_f := 2045;
        ELSIF x = 13227 THEN
            sigmoid_f := 2045;
        ELSIF x = 13228 THEN
            sigmoid_f := 2045;
        ELSIF x = 13229 THEN
            sigmoid_f := 2045;
        ELSIF x = 13230 THEN
            sigmoid_f := 2045;
        ELSIF x = 13231 THEN
            sigmoid_f := 2045;
        ELSIF x = 13232 THEN
            sigmoid_f := 2045;
        ELSIF x = 13233 THEN
            sigmoid_f := 2045;
        ELSIF x = 13234 THEN
            sigmoid_f := 2045;
        ELSIF x = 13235 THEN
            sigmoid_f := 2045;
        ELSIF x = 13236 THEN
            sigmoid_f := 2045;
        ELSIF x = 13237 THEN
            sigmoid_f := 2045;
        ELSIF x = 13238 THEN
            sigmoid_f := 2045;
        ELSIF x = 13239 THEN
            sigmoid_f := 2045;
        ELSIF x = 13240 THEN
            sigmoid_f := 2045;
        ELSIF x = 13241 THEN
            sigmoid_f := 2045;
        ELSIF x = 13242 THEN
            sigmoid_f := 2045;
        ELSIF x = 13243 THEN
            sigmoid_f := 2045;
        ELSIF x = 13244 THEN
            sigmoid_f := 2045;
        ELSIF x = 13245 THEN
            sigmoid_f := 2045;
        ELSIF x = 13246 THEN
            sigmoid_f := 2045;
        ELSIF x = 13247 THEN
            sigmoid_f := 2045;
        ELSIF x = 13248 THEN
            sigmoid_f := 2045;
        ELSIF x = 13249 THEN
            sigmoid_f := 2045;
        ELSIF x = 13250 THEN
            sigmoid_f := 2045;
        ELSIF x = 13251 THEN
            sigmoid_f := 2045;
        ELSIF x = 13252 THEN
            sigmoid_f := 2045;
        ELSIF x = 13253 THEN
            sigmoid_f := 2045;
        ELSIF x = 13254 THEN
            sigmoid_f := 2045;
        ELSIF x = 13255 THEN
            sigmoid_f := 2045;
        ELSIF x = 13256 THEN
            sigmoid_f := 2045;
        ELSIF x = 13257 THEN
            sigmoid_f := 2045;
        ELSIF x = 13258 THEN
            sigmoid_f := 2045;
        ELSIF x = 13259 THEN
            sigmoid_f := 2045;
        ELSIF x = 13260 THEN
            sigmoid_f := 2045;
        ELSIF x = 13261 THEN
            sigmoid_f := 2045;
        ELSIF x = 13262 THEN
            sigmoid_f := 2045;
        ELSIF x = 13263 THEN
            sigmoid_f := 2045;
        ELSIF x = 13264 THEN
            sigmoid_f := 2045;
        ELSIF x = 13265 THEN
            sigmoid_f := 2045;
        ELSIF x = 13266 THEN
            sigmoid_f := 2045;
        ELSIF x = 13267 THEN
            sigmoid_f := 2045;
        ELSIF x = 13268 THEN
            sigmoid_f := 2045;
        ELSIF x = 13269 THEN
            sigmoid_f := 2045;
        ELSIF x = 13270 THEN
            sigmoid_f := 2045;
        ELSIF x = 13271 THEN
            sigmoid_f := 2045;
        ELSIF x = 13272 THEN
            sigmoid_f := 2045;
        ELSIF x = 13273 THEN
            sigmoid_f := 2045;
        ELSIF x = 13274 THEN
            sigmoid_f := 2045;
        ELSIF x = 13275 THEN
            sigmoid_f := 2045;
        ELSIF x = 13276 THEN
            sigmoid_f := 2045;
        ELSIF x = 13277 THEN
            sigmoid_f := 2045;
        ELSIF x = 13278 THEN
            sigmoid_f := 2045;
        ELSIF x = 13279 THEN
            sigmoid_f := 2045;
        ELSIF x = 13280 THEN
            sigmoid_f := 2045;
        ELSIF x = 13281 THEN
            sigmoid_f := 2045;
        ELSIF x = 13282 THEN
            sigmoid_f := 2045;
        ELSIF x = 13283 THEN
            sigmoid_f := 2045;
        ELSIF x = 13284 THEN
            sigmoid_f := 2045;
        ELSIF x = 13285 THEN
            sigmoid_f := 2045;
        ELSIF x = 13286 THEN
            sigmoid_f := 2045;
        ELSIF x = 13287 THEN
            sigmoid_f := 2045;
        ELSIF x = 13288 THEN
            sigmoid_f := 2045;
        ELSIF x = 13289 THEN
            sigmoid_f := 2045;
        ELSIF x = 13290 THEN
            sigmoid_f := 2045;
        ELSIF x = 13291 THEN
            sigmoid_f := 2045;
        ELSIF x = 13292 THEN
            sigmoid_f := 2045;
        ELSIF x = 13293 THEN
            sigmoid_f := 2045;
        ELSIF x = 13294 THEN
            sigmoid_f := 2045;
        ELSIF x = 13295 THEN
            sigmoid_f := 2045;
        ELSIF x = 13296 THEN
            sigmoid_f := 2045;
        ELSIF x = 13297 THEN
            sigmoid_f := 2045;
        ELSIF x = 13298 THEN
            sigmoid_f := 2045;
        ELSIF x = 13299 THEN
            sigmoid_f := 2045;
        ELSIF x = 13300 THEN
            sigmoid_f := 2045;
        ELSIF x = 13301 THEN
            sigmoid_f := 2045;
        ELSIF x = 13302 THEN
            sigmoid_f := 2045;
        ELSIF x = 13303 THEN
            sigmoid_f := 2045;
        ELSIF x = 13304 THEN
            sigmoid_f := 2045;
        ELSIF x = 13305 THEN
            sigmoid_f := 2045;
        ELSIF x = 13306 THEN
            sigmoid_f := 2045;
        ELSIF x = 13307 THEN
            sigmoid_f := 2045;
        ELSIF x = 13308 THEN
            sigmoid_f := 2045;
        ELSIF x = 13309 THEN
            sigmoid_f := 2045;
        ELSIF x = 13310 THEN
            sigmoid_f := 2045;
        ELSIF x = 13311 THEN
            sigmoid_f := 2045;
        ELSIF x = 13312 THEN
            sigmoid_f := 2045;
        ELSIF x = 13313 THEN
            sigmoid_f := 2045;
        ELSIF x = 13314 THEN
            sigmoid_f := 2045;
        ELSIF x = 13315 THEN
            sigmoid_f := 2045;
        ELSIF x = 13316 THEN
            sigmoid_f := 2045;
        ELSIF x = 13317 THEN
            sigmoid_f := 2045;
        ELSIF x = 13318 THEN
            sigmoid_f := 2045;
        ELSIF x = 13319 THEN
            sigmoid_f := 2045;
        ELSIF x = 13320 THEN
            sigmoid_f := 2045;
        ELSIF x = 13321 THEN
            sigmoid_f := 2045;
        ELSIF x = 13322 THEN
            sigmoid_f := 2045;
        ELSIF x = 13323 THEN
            sigmoid_f := 2045;
        ELSIF x = 13324 THEN
            sigmoid_f := 2045;
        ELSIF x = 13325 THEN
            sigmoid_f := 2045;
        ELSIF x = 13326 THEN
            sigmoid_f := 2045;
        ELSIF x = 13327 THEN
            sigmoid_f := 2045;
        ELSIF x = 13328 THEN
            sigmoid_f := 2045;
        ELSIF x = 13329 THEN
            sigmoid_f := 2045;
        ELSIF x = 13330 THEN
            sigmoid_f := 2045;
        ELSIF x = 13331 THEN
            sigmoid_f := 2045;
        ELSIF x = 13332 THEN
            sigmoid_f := 2045;
        ELSIF x = 13333 THEN
            sigmoid_f := 2045;
        ELSIF x = 13334 THEN
            sigmoid_f := 2045;
        ELSIF x = 13335 THEN
            sigmoid_f := 2045;
        ELSIF x = 13336 THEN
            sigmoid_f := 2045;
        ELSIF x = 13337 THEN
            sigmoid_f := 2045;
        ELSIF x = 13338 THEN
            sigmoid_f := 2045;
        ELSIF x = 13339 THEN
            sigmoid_f := 2045;
        ELSIF x = 13340 THEN
            sigmoid_f := 2045;
        ELSIF x = 13341 THEN
            sigmoid_f := 2045;
        ELSIF x = 13342 THEN
            sigmoid_f := 2045;
        ELSIF x = 13343 THEN
            sigmoid_f := 2045;
        ELSIF x = 13344 THEN
            sigmoid_f := 2045;
        ELSIF x = 13345 THEN
            sigmoid_f := 2045;
        ELSIF x = 13346 THEN
            sigmoid_f := 2045;
        ELSIF x = 13347 THEN
            sigmoid_f := 2045;
        ELSIF x = 13348 THEN
            sigmoid_f := 2045;
        ELSIF x = 13349 THEN
            sigmoid_f := 2045;
        ELSIF x = 13350 THEN
            sigmoid_f := 2045;
        ELSIF x = 13351 THEN
            sigmoid_f := 2045;
        ELSIF x = 13352 THEN
            sigmoid_f := 2045;
        ELSIF x = 13353 THEN
            sigmoid_f := 2045;
        ELSIF x = 13354 THEN
            sigmoid_f := 2045;
        ELSIF x = 13355 THEN
            sigmoid_f := 2045;
        ELSIF x = 13356 THEN
            sigmoid_f := 2045;
        ELSIF x = 13357 THEN
            sigmoid_f := 2045;
        ELSIF x = 13358 THEN
            sigmoid_f := 2045;
        ELSIF x = 13359 THEN
            sigmoid_f := 2045;
        ELSIF x = 13360 THEN
            sigmoid_f := 2045;
        ELSIF x = 13361 THEN
            sigmoid_f := 2045;
        ELSIF x = 13362 THEN
            sigmoid_f := 2045;
        ELSIF x = 13363 THEN
            sigmoid_f := 2045;
        ELSIF x = 13364 THEN
            sigmoid_f := 2045;
        ELSIF x = 13365 THEN
            sigmoid_f := 2045;
        ELSIF x = 13366 THEN
            sigmoid_f := 2045;
        ELSIF x = 13367 THEN
            sigmoid_f := 2045;
        ELSIF x = 13368 THEN
            sigmoid_f := 2045;
        ELSIF x = 13369 THEN
            sigmoid_f := 2045;
        ELSIF x = 13370 THEN
            sigmoid_f := 2045;
        ELSIF x = 13371 THEN
            sigmoid_f := 2045;
        ELSIF x = 13372 THEN
            sigmoid_f := 2045;
        ELSIF x = 13373 THEN
            sigmoid_f := 2045;
        ELSIF x = 13374 THEN
            sigmoid_f := 2045;
        ELSIF x = 13375 THEN
            sigmoid_f := 2045;
        ELSIF x = 13376 THEN
            sigmoid_f := 2045;
        ELSIF x = 13377 THEN
            sigmoid_f := 2045;
        ELSIF x = 13378 THEN
            sigmoid_f := 2045;
        ELSIF x = 13379 THEN
            sigmoid_f := 2045;
        ELSIF x = 13380 THEN
            sigmoid_f := 2045;
        ELSIF x = 13381 THEN
            sigmoid_f := 2045;
        ELSIF x = 13382 THEN
            sigmoid_f := 2045;
        ELSIF x = 13383 THEN
            sigmoid_f := 2045;
        ELSIF x = 13384 THEN
            sigmoid_f := 2045;
        ELSIF x = 13385 THEN
            sigmoid_f := 2045;
        ELSIF x = 13386 THEN
            sigmoid_f := 2045;
        ELSIF x = 13387 THEN
            sigmoid_f := 2045;
        ELSIF x = 13388 THEN
            sigmoid_f := 2045;
        ELSIF x = 13389 THEN
            sigmoid_f := 2045;
        ELSIF x = 13390 THEN
            sigmoid_f := 2045;
        ELSIF x = 13391 THEN
            sigmoid_f := 2045;
        ELSIF x = 13392 THEN
            sigmoid_f := 2045;
        ELSIF x = 13393 THEN
            sigmoid_f := 2045;
        ELSIF x = 13394 THEN
            sigmoid_f := 2045;
        ELSIF x = 13395 THEN
            sigmoid_f := 2045;
        ELSIF x = 13396 THEN
            sigmoid_f := 2045;
        ELSIF x = 13397 THEN
            sigmoid_f := 2045;
        ELSIF x = 13398 THEN
            sigmoid_f := 2045;
        ELSIF x = 13399 THEN
            sigmoid_f := 2045;
        ELSIF x = 13400 THEN
            sigmoid_f := 2045;
        ELSIF x = 13401 THEN
            sigmoid_f := 2045;
        ELSIF x = 13402 THEN
            sigmoid_f := 2045;
        ELSIF x = 13403 THEN
            sigmoid_f := 2045;
        ELSIF x = 13404 THEN
            sigmoid_f := 2045;
        ELSIF x = 13405 THEN
            sigmoid_f := 2045;
        ELSIF x = 13406 THEN
            sigmoid_f := 2045;
        ELSIF x = 13407 THEN
            sigmoid_f := 2045;
        ELSIF x = 13408 THEN
            sigmoid_f := 2045;
        ELSIF x = 13409 THEN
            sigmoid_f := 2045;
        ELSIF x = 13410 THEN
            sigmoid_f := 2045;
        ELSIF x = 13411 THEN
            sigmoid_f := 2045;
        ELSIF x = 13412 THEN
            sigmoid_f := 2045;
        ELSIF x = 13413 THEN
            sigmoid_f := 2045;
        ELSIF x = 13414 THEN
            sigmoid_f := 2045;
        ELSIF x = 13415 THEN
            sigmoid_f := 2045;
        ELSIF x = 13416 THEN
            sigmoid_f := 2045;
        ELSIF x = 13417 THEN
            sigmoid_f := 2045;
        ELSIF x = 13418 THEN
            sigmoid_f := 2045;
        ELSIF x = 13419 THEN
            sigmoid_f := 2045;
        ELSIF x = 13420 THEN
            sigmoid_f := 2045;
        ELSIF x = 13421 THEN
            sigmoid_f := 2045;
        ELSIF x = 13422 THEN
            sigmoid_f := 2045;
        ELSIF x = 13423 THEN
            sigmoid_f := 2045;
        ELSIF x = 13424 THEN
            sigmoid_f := 2045;
        ELSIF x = 13425 THEN
            sigmoid_f := 2045;
        ELSIF x = 13426 THEN
            sigmoid_f := 2045;
        ELSIF x = 13427 THEN
            sigmoid_f := 2045;
        ELSIF x = 13428 THEN
            sigmoid_f := 2045;
        ELSIF x = 13429 THEN
            sigmoid_f := 2045;
        ELSIF x = 13430 THEN
            sigmoid_f := 2045;
        ELSIF x = 13431 THEN
            sigmoid_f := 2045;
        ELSIF x = 13432 THEN
            sigmoid_f := 2045;
        ELSIF x = 13433 THEN
            sigmoid_f := 2045;
        ELSIF x = 13434 THEN
            sigmoid_f := 2045;
        ELSIF x = 13435 THEN
            sigmoid_f := 2045;
        ELSIF x = 13436 THEN
            sigmoid_f := 2045;
        ELSIF x = 13437 THEN
            sigmoid_f := 2045;
        ELSIF x = 13438 THEN
            sigmoid_f := 2045;
        ELSIF x = 13439 THEN
            sigmoid_f := 2045;
        ELSIF x = 13440 THEN
            sigmoid_f := 2045;
        ELSIF x = 13441 THEN
            sigmoid_f := 2045;
        ELSIF x = 13442 THEN
            sigmoid_f := 2045;
        ELSIF x = 13443 THEN
            sigmoid_f := 2045;
        ELSIF x = 13444 THEN
            sigmoid_f := 2045;
        ELSIF x = 13445 THEN
            sigmoid_f := 2045;
        ELSIF x = 13446 THEN
            sigmoid_f := 2045;
        ELSIF x = 13447 THEN
            sigmoid_f := 2045;
        ELSIF x = 13448 THEN
            sigmoid_f := 2045;
        ELSIF x = 13449 THEN
            sigmoid_f := 2045;
        ELSIF x = 13450 THEN
            sigmoid_f := 2045;
        ELSIF x = 13451 THEN
            sigmoid_f := 2045;
        ELSIF x = 13452 THEN
            sigmoid_f := 2045;
        ELSIF x = 13453 THEN
            sigmoid_f := 2045;
        ELSIF x = 13454 THEN
            sigmoid_f := 2045;
        ELSIF x = 13455 THEN
            sigmoid_f := 2045;
        ELSIF x = 13456 THEN
            sigmoid_f := 2045;
        ELSIF x = 13457 THEN
            sigmoid_f := 2045;
        ELSIF x = 13458 THEN
            sigmoid_f := 2045;
        ELSIF x = 13459 THEN
            sigmoid_f := 2045;
        ELSIF x = 13460 THEN
            sigmoid_f := 2045;
        ELSIF x = 13461 THEN
            sigmoid_f := 2045;
        ELSIF x = 13462 THEN
            sigmoid_f := 2045;
        ELSIF x = 13463 THEN
            sigmoid_f := 2045;
        ELSIF x = 13464 THEN
            sigmoid_f := 2045;
        ELSIF x = 13465 THEN
            sigmoid_f := 2045;
        ELSIF x = 13466 THEN
            sigmoid_f := 2045;
        ELSIF x = 13467 THEN
            sigmoid_f := 2045;
        ELSIF x = 13468 THEN
            sigmoid_f := 2045;
        ELSIF x = 13469 THEN
            sigmoid_f := 2045;
        ELSIF x = 13470 THEN
            sigmoid_f := 2045;
        ELSIF x = 13471 THEN
            sigmoid_f := 2045;
        ELSIF x = 13472 THEN
            sigmoid_f := 2045;
        ELSIF x = 13473 THEN
            sigmoid_f := 2045;
        ELSIF x = 13474 THEN
            sigmoid_f := 2045;
        ELSIF x = 13475 THEN
            sigmoid_f := 2045;
        ELSIF x = 13476 THEN
            sigmoid_f := 2045;
        ELSIF x = 13477 THEN
            sigmoid_f := 2045;
        ELSIF x = 13478 THEN
            sigmoid_f := 2045;
        ELSIF x = 13479 THEN
            sigmoid_f := 2045;
        ELSIF x = 13480 THEN
            sigmoid_f := 2045;
        ELSIF x = 13481 THEN
            sigmoid_f := 2045;
        ELSIF x = 13482 THEN
            sigmoid_f := 2045;
        ELSIF x = 13483 THEN
            sigmoid_f := 2045;
        ELSIF x = 13484 THEN
            sigmoid_f := 2045;
        ELSIF x = 13485 THEN
            sigmoid_f := 2045;
        ELSIF x = 13486 THEN
            sigmoid_f := 2045;
        ELSIF x = 13487 THEN
            sigmoid_f := 2045;
        ELSIF x = 13488 THEN
            sigmoid_f := 2045;
        ELSIF x = 13489 THEN
            sigmoid_f := 2045;
        ELSIF x = 13490 THEN
            sigmoid_f := 2045;
        ELSIF x = 13491 THEN
            sigmoid_f := 2045;
        ELSIF x = 13492 THEN
            sigmoid_f := 2045;
        ELSIF x = 13493 THEN
            sigmoid_f := 2045;
        ELSIF x = 13494 THEN
            sigmoid_f := 2045;
        ELSIF x = 13495 THEN
            sigmoid_f := 2045;
        ELSIF x = 13496 THEN
            sigmoid_f := 2045;
        ELSIF x = 13497 THEN
            sigmoid_f := 2045;
        ELSIF x = 13498 THEN
            sigmoid_f := 2045;
        ELSIF x = 13499 THEN
            sigmoid_f := 2045;
        ELSIF x = 13500 THEN
            sigmoid_f := 2045;
        ELSIF x = 13501 THEN
            sigmoid_f := 2045;
        ELSIF x = 13502 THEN
            sigmoid_f := 2045;
        ELSIF x = 13503 THEN
            sigmoid_f := 2045;
        ELSIF x = 13504 THEN
            sigmoid_f := 2045;
        ELSIF x = 13505 THEN
            sigmoid_f := 2045;
        ELSIF x = 13506 THEN
            sigmoid_f := 2045;
        ELSIF x = 13507 THEN
            sigmoid_f := 2045;
        ELSIF x = 13508 THEN
            sigmoid_f := 2045;
        ELSIF x = 13509 THEN
            sigmoid_f := 2045;
        ELSIF x = 13510 THEN
            sigmoid_f := 2045;
        ELSIF x = 13511 THEN
            sigmoid_f := 2045;
        ELSIF x = 13512 THEN
            sigmoid_f := 2045;
        ELSIF x = 13513 THEN
            sigmoid_f := 2045;
        ELSIF x = 13514 THEN
            sigmoid_f := 2045;
        ELSIF x = 13515 THEN
            sigmoid_f := 2045;
        ELSIF x = 13516 THEN
            sigmoid_f := 2045;
        ELSIF x = 13517 THEN
            sigmoid_f := 2045;
        ELSIF x = 13518 THEN
            sigmoid_f := 2045;
        ELSIF x = 13519 THEN
            sigmoid_f := 2045;
        ELSIF x = 13520 THEN
            sigmoid_f := 2045;
        ELSIF x = 13521 THEN
            sigmoid_f := 2045;
        ELSIF x = 13522 THEN
            sigmoid_f := 2045;
        ELSIF x = 13523 THEN
            sigmoid_f := 2045;
        ELSIF x = 13524 THEN
            sigmoid_f := 2045;
        ELSIF x = 13525 THEN
            sigmoid_f := 2045;
        ELSIF x = 13526 THEN
            sigmoid_f := 2045;
        ELSIF x = 13527 THEN
            sigmoid_f := 2045;
        ELSIF x = 13528 THEN
            sigmoid_f := 2045;
        ELSIF x = 13529 THEN
            sigmoid_f := 2045;
        ELSIF x = 13530 THEN
            sigmoid_f := 2045;
        ELSIF x = 13531 THEN
            sigmoid_f := 2045;
        ELSIF x = 13532 THEN
            sigmoid_f := 2045;
        ELSIF x = 13533 THEN
            sigmoid_f := 2045;
        ELSIF x = 13534 THEN
            sigmoid_f := 2045;
        ELSIF x = 13535 THEN
            sigmoid_f := 2045;
        ELSIF x = 13536 THEN
            sigmoid_f := 2045;
        ELSIF x = 13537 THEN
            sigmoid_f := 2045;
        ELSIF x = 13538 THEN
            sigmoid_f := 2045;
        ELSIF x = 13539 THEN
            sigmoid_f := 2045;
        ELSIF x = 13540 THEN
            sigmoid_f := 2045;
        ELSIF x = 13541 THEN
            sigmoid_f := 2045;
        ELSIF x = 13542 THEN
            sigmoid_f := 2045;
        ELSIF x = 13543 THEN
            sigmoid_f := 2045;
        ELSIF x = 13544 THEN
            sigmoid_f := 2045;
        ELSIF x = 13545 THEN
            sigmoid_f := 2045;
        ELSIF x = 13546 THEN
            sigmoid_f := 2045;
        ELSIF x = 13547 THEN
            sigmoid_f := 2045;
        ELSIF x = 13548 THEN
            sigmoid_f := 2045;
        ELSIF x = 13549 THEN
            sigmoid_f := 2045;
        ELSIF x = 13550 THEN
            sigmoid_f := 2045;
        ELSIF x = 13551 THEN
            sigmoid_f := 2045;
        ELSIF x = 13552 THEN
            sigmoid_f := 2045;
        ELSIF x = 13553 THEN
            sigmoid_f := 2045;
        ELSIF x = 13554 THEN
            sigmoid_f := 2045;
        ELSIF x = 13555 THEN
            sigmoid_f := 2045;
        ELSIF x = 13556 THEN
            sigmoid_f := 2045;
        ELSIF x = 13557 THEN
            sigmoid_f := 2045;
        ELSIF x = 13558 THEN
            sigmoid_f := 2045;
        ELSIF x = 13559 THEN
            sigmoid_f := 2045;
        ELSIF x = 13560 THEN
            sigmoid_f := 2045;
        ELSIF x = 13561 THEN
            sigmoid_f := 2045;
        ELSIF x = 13562 THEN
            sigmoid_f := 2045;
        ELSIF x = 13563 THEN
            sigmoid_f := 2045;
        ELSIF x = 13564 THEN
            sigmoid_f := 2045;
        ELSIF x = 13565 THEN
            sigmoid_f := 2045;
        ELSIF x = 13566 THEN
            sigmoid_f := 2045;
        ELSIF x = 13567 THEN
            sigmoid_f := 2045;
        ELSIF x = 13568 THEN
            sigmoid_f := 2045;
        ELSIF x = 13569 THEN
            sigmoid_f := 2045;
        ELSIF x = 13570 THEN
            sigmoid_f := 2045;
        ELSIF x = 13571 THEN
            sigmoid_f := 2045;
        ELSIF x = 13572 THEN
            sigmoid_f := 2045;
        ELSIF x = 13573 THEN
            sigmoid_f := 2045;
        ELSIF x = 13574 THEN
            sigmoid_f := 2045;
        ELSIF x = 13575 THEN
            sigmoid_f := 2045;
        ELSIF x = 13576 THEN
            sigmoid_f := 2045;
        ELSIF x = 13577 THEN
            sigmoid_f := 2045;
        ELSIF x = 13578 THEN
            sigmoid_f := 2045;
        ELSIF x = 13579 THEN
            sigmoid_f := 2045;
        ELSIF x = 13580 THEN
            sigmoid_f := 2045;
        ELSIF x = 13581 THEN
            sigmoid_f := 2045;
        ELSIF x = 13582 THEN
            sigmoid_f := 2045;
        ELSIF x = 13583 THEN
            sigmoid_f := 2045;
        ELSIF x = 13584 THEN
            sigmoid_f := 2045;
        ELSIF x = 13585 THEN
            sigmoid_f := 2045;
        ELSIF x = 13586 THEN
            sigmoid_f := 2045;
        ELSIF x = 13587 THEN
            sigmoid_f := 2045;
        ELSIF x = 13588 THEN
            sigmoid_f := 2045;
        ELSIF x = 13589 THEN
            sigmoid_f := 2045;
        ELSIF x = 13590 THEN
            sigmoid_f := 2045;
        ELSIF x = 13591 THEN
            sigmoid_f := 2045;
        ELSIF x = 13592 THEN
            sigmoid_f := 2045;
        ELSIF x = 13593 THEN
            sigmoid_f := 2045;
        ELSIF x = 13594 THEN
            sigmoid_f := 2045;
        ELSIF x = 13595 THEN
            sigmoid_f := 2045;
        ELSIF x = 13596 THEN
            sigmoid_f := 2045;
        ELSIF x = 13597 THEN
            sigmoid_f := 2045;
        ELSIF x = 13598 THEN
            sigmoid_f := 2045;
        ELSIF x = 13599 THEN
            sigmoid_f := 2045;
        ELSIF x = 13600 THEN
            sigmoid_f := 2045;
        ELSIF x = 13601 THEN
            sigmoid_f := 2045;
        ELSIF x = 13602 THEN
            sigmoid_f := 2045;
        ELSIF x = 13603 THEN
            sigmoid_f := 2045;
        ELSIF x = 13604 THEN
            sigmoid_f := 2045;
        ELSIF x = 13605 THEN
            sigmoid_f := 2045;
        ELSIF x = 13606 THEN
            sigmoid_f := 2045;
        ELSIF x = 13607 THEN
            sigmoid_f := 2045;
        ELSIF x = 13608 THEN
            sigmoid_f := 2045;
        ELSIF x = 13609 THEN
            sigmoid_f := 2045;
        ELSIF x = 13610 THEN
            sigmoid_f := 2045;
        ELSIF x = 13611 THEN
            sigmoid_f := 2045;
        ELSIF x = 13612 THEN
            sigmoid_f := 2045;
        ELSIF x = 13613 THEN
            sigmoid_f := 2045;
        ELSIF x = 13614 THEN
            sigmoid_f := 2045;
        ELSIF x = 13615 THEN
            sigmoid_f := 2045;
        ELSIF x = 13616 THEN
            sigmoid_f := 2045;
        ELSIF x = 13617 THEN
            sigmoid_f := 2045;
        ELSIF x = 13618 THEN
            sigmoid_f := 2045;
        ELSIF x = 13619 THEN
            sigmoid_f := 2045;
        ELSIF x = 13620 THEN
            sigmoid_f := 2045;
        ELSIF x = 13621 THEN
            sigmoid_f := 2045;
        ELSIF x = 13622 THEN
            sigmoid_f := 2045;
        ELSIF x = 13623 THEN
            sigmoid_f := 2045;
        ELSIF x = 13624 THEN
            sigmoid_f := 2045;
        ELSIF x = 13625 THEN
            sigmoid_f := 2045;
        ELSIF x = 13626 THEN
            sigmoid_f := 2045;
        ELSIF x = 13627 THEN
            sigmoid_f := 2045;
        ELSIF x = 13628 THEN
            sigmoid_f := 2045;
        ELSIF x = 13629 THEN
            sigmoid_f := 2045;
        ELSIF x = 13630 THEN
            sigmoid_f := 2045;
        ELSIF x = 13631 THEN
            sigmoid_f := 2045;
        ELSIF x = 13632 THEN
            sigmoid_f := 2045;
        ELSIF x = 13633 THEN
            sigmoid_f := 2045;
        ELSIF x = 13634 THEN
            sigmoid_f := 2045;
        ELSIF x = 13635 THEN
            sigmoid_f := 2045;
        ELSIF x = 13636 THEN
            sigmoid_f := 2045;
        ELSIF x = 13637 THEN
            sigmoid_f := 2045;
        ELSIF x = 13638 THEN
            sigmoid_f := 2045;
        ELSIF x = 13639 THEN
            sigmoid_f := 2045;
        ELSIF x = 13640 THEN
            sigmoid_f := 2045;
        ELSIF x = 13641 THEN
            sigmoid_f := 2045;
        ELSIF x = 13642 THEN
            sigmoid_f := 2045;
        ELSIF x = 13643 THEN
            sigmoid_f := 2045;
        ELSIF x = 13644 THEN
            sigmoid_f := 2045;
        ELSIF x = 13645 THEN
            sigmoid_f := 2045;
        ELSIF x = 13646 THEN
            sigmoid_f := 2045;
        ELSIF x = 13647 THEN
            sigmoid_f := 2045;
        ELSIF x = 13648 THEN
            sigmoid_f := 2045;
        ELSIF x = 13649 THEN
            sigmoid_f := 2045;
        ELSIF x = 13650 THEN
            sigmoid_f := 2045;
        ELSIF x = 13651 THEN
            sigmoid_f := 2045;
        ELSIF x = 13652 THEN
            sigmoid_f := 2045;
        ELSIF x = 13653 THEN
            sigmoid_f := 2045;
        ELSIF x = 13654 THEN
            sigmoid_f := 2045;
        ELSIF x = 13655 THEN
            sigmoid_f := 2045;
        ELSIF x = 13656 THEN
            sigmoid_f := 2045;
        ELSIF x = 13657 THEN
            sigmoid_f := 2045;
        ELSIF x = 13658 THEN
            sigmoid_f := 2045;
        ELSIF x = 13659 THEN
            sigmoid_f := 2045;
        ELSIF x = 13660 THEN
            sigmoid_f := 2045;
        ELSIF x = 13661 THEN
            sigmoid_f := 2045;
        ELSIF x = 13662 THEN
            sigmoid_f := 2045;
        ELSIF x = 13663 THEN
            sigmoid_f := 2045;
        ELSIF x = 13664 THEN
            sigmoid_f := 2045;
        ELSIF x = 13665 THEN
            sigmoid_f := 2045;
        ELSIF x = 13666 THEN
            sigmoid_f := 2045;
        ELSIF x = 13667 THEN
            sigmoid_f := 2045;
        ELSIF x = 13668 THEN
            sigmoid_f := 2045;
        ELSIF x = 13669 THEN
            sigmoid_f := 2045;
        ELSIF x = 13670 THEN
            sigmoid_f := 2045;
        ELSIF x = 13671 THEN
            sigmoid_f := 2045;
        ELSIF x = 13672 THEN
            sigmoid_f := 2045;
        ELSIF x = 13673 THEN
            sigmoid_f := 2045;
        ELSIF x = 13674 THEN
            sigmoid_f := 2045;
        ELSIF x = 13675 THEN
            sigmoid_f := 2045;
        ELSIF x = 13676 THEN
            sigmoid_f := 2045;
        ELSIF x = 13677 THEN
            sigmoid_f := 2045;
        ELSIF x = 13678 THEN
            sigmoid_f := 2045;
        ELSIF x = 13679 THEN
            sigmoid_f := 2045;
        ELSIF x = 13680 THEN
            sigmoid_f := 2045;
        ELSIF x = 13681 THEN
            sigmoid_f := 2045;
        ELSIF x = 13682 THEN
            sigmoid_f := 2045;
        ELSIF x = 13683 THEN
            sigmoid_f := 2045;
        ELSIF x = 13684 THEN
            sigmoid_f := 2045;
        ELSIF x = 13685 THEN
            sigmoid_f := 2045;
        ELSIF x = 13686 THEN
            sigmoid_f := 2045;
        ELSIF x = 13687 THEN
            sigmoid_f := 2045;
        ELSIF x = 13688 THEN
            sigmoid_f := 2045;
        ELSIF x = 13689 THEN
            sigmoid_f := 2045;
        ELSIF x = 13690 THEN
            sigmoid_f := 2045;
        ELSIF x = 13691 THEN
            sigmoid_f := 2045;
        ELSIF x = 13692 THEN
            sigmoid_f := 2045;
        ELSIF x = 13693 THEN
            sigmoid_f := 2045;
        ELSIF x = 13694 THEN
            sigmoid_f := 2045;
        ELSIF x = 13695 THEN
            sigmoid_f := 2045;
        ELSIF x = 13696 THEN
            sigmoid_f := 2045;
        ELSIF x = 13697 THEN
            sigmoid_f := 2045;
        ELSIF x = 13698 THEN
            sigmoid_f := 2045;
        ELSIF x = 13699 THEN
            sigmoid_f := 2045;
        ELSIF x = 13700 THEN
            sigmoid_f := 2045;
        ELSIF x = 13701 THEN
            sigmoid_f := 2045;
        ELSIF x = 13702 THEN
            sigmoid_f := 2045;
        ELSIF x = 13703 THEN
            sigmoid_f := 2045;
        ELSIF x = 13704 THEN
            sigmoid_f := 2045;
        ELSIF x = 13705 THEN
            sigmoid_f := 2045;
        ELSIF x = 13706 THEN
            sigmoid_f := 2045;
        ELSIF x = 13707 THEN
            sigmoid_f := 2045;
        ELSIF x = 13708 THEN
            sigmoid_f := 2045;
        ELSIF x = 13709 THEN
            sigmoid_f := 2045;
        ELSIF x = 13710 THEN
            sigmoid_f := 2045;
        ELSIF x = 13711 THEN
            sigmoid_f := 2045;
        ELSIF x = 13712 THEN
            sigmoid_f := 2045;
        ELSIF x = 13713 THEN
            sigmoid_f := 2045;
        ELSIF x = 13714 THEN
            sigmoid_f := 2045;
        ELSIF x = 13715 THEN
            sigmoid_f := 2045;
        ELSIF x = 13716 THEN
            sigmoid_f := 2045;
        ELSIF x = 13717 THEN
            sigmoid_f := 2045;
        ELSIF x = 13718 THEN
            sigmoid_f := 2045;
        ELSIF x = 13719 THEN
            sigmoid_f := 2045;
        ELSIF x = 13720 THEN
            sigmoid_f := 2045;
        ELSIF x = 13721 THEN
            sigmoid_f := 2045;
        ELSIF x = 13722 THEN
            sigmoid_f := 2045;
        ELSIF x = 13723 THEN
            sigmoid_f := 2045;
        ELSIF x = 13724 THEN
            sigmoid_f := 2045;
        ELSIF x = 13725 THEN
            sigmoid_f := 2045;
        ELSIF x = 13726 THEN
            sigmoid_f := 2045;
        ELSIF x = 13727 THEN
            sigmoid_f := 2045;
        ELSIF x = 13728 THEN
            sigmoid_f := 2045;
        ELSIF x = 13729 THEN
            sigmoid_f := 2045;
        ELSIF x = 13730 THEN
            sigmoid_f := 2045;
        ELSIF x = 13731 THEN
            sigmoid_f := 2045;
        ELSIF x = 13732 THEN
            sigmoid_f := 2045;
        ELSIF x = 13733 THEN
            sigmoid_f := 2045;
        ELSIF x = 13734 THEN
            sigmoid_f := 2045;
        ELSIF x = 13735 THEN
            sigmoid_f := 2045;
        ELSIF x = 13736 THEN
            sigmoid_f := 2045;
        ELSIF x = 13737 THEN
            sigmoid_f := 2045;
        ELSIF x = 13738 THEN
            sigmoid_f := 2045;
        ELSIF x = 13739 THEN
            sigmoid_f := 2045;
        ELSIF x = 13740 THEN
            sigmoid_f := 2045;
        ELSIF x = 13741 THEN
            sigmoid_f := 2045;
        ELSIF x = 13742 THEN
            sigmoid_f := 2045;
        ELSIF x = 13743 THEN
            sigmoid_f := 2045;
        ELSIF x = 13744 THEN
            sigmoid_f := 2045;
        ELSIF x = 13745 THEN
            sigmoid_f := 2045;
        ELSIF x = 13746 THEN
            sigmoid_f := 2045;
        ELSIF x = 13747 THEN
            sigmoid_f := 2045;
        ELSIF x = 13748 THEN
            sigmoid_f := 2045;
        ELSIF x = 13749 THEN
            sigmoid_f := 2045;
        ELSIF x = 13750 THEN
            sigmoid_f := 2045;
        ELSIF x = 13751 THEN
            sigmoid_f := 2045;
        ELSIF x = 13752 THEN
            sigmoid_f := 2045;
        ELSIF x = 13753 THEN
            sigmoid_f := 2045;
        ELSIF x = 13754 THEN
            sigmoid_f := 2045;
        ELSIF x = 13755 THEN
            sigmoid_f := 2045;
        ELSIF x = 13756 THEN
            sigmoid_f := 2045;
        ELSIF x = 13757 THEN
            sigmoid_f := 2045;
        ELSIF x = 13758 THEN
            sigmoid_f := 2045;
        ELSIF x = 13759 THEN
            sigmoid_f := 2045;
        ELSIF x = 13760 THEN
            sigmoid_f := 2045;
        ELSIF x = 13761 THEN
            sigmoid_f := 2045;
        ELSIF x = 13762 THEN
            sigmoid_f := 2045;
        ELSIF x = 13763 THEN
            sigmoid_f := 2045;
        ELSIF x = 13764 THEN
            sigmoid_f := 2045;
        ELSIF x = 13765 THEN
            sigmoid_f := 2045;
        ELSIF x = 13766 THEN
            sigmoid_f := 2045;
        ELSIF x = 13767 THEN
            sigmoid_f := 2045;
        ELSIF x = 13768 THEN
            sigmoid_f := 2045;
        ELSIF x = 13769 THEN
            sigmoid_f := 2045;
        ELSIF x = 13770 THEN
            sigmoid_f := 2045;
        ELSIF x = 13771 THEN
            sigmoid_f := 2045;
        ELSIF x = 13772 THEN
            sigmoid_f := 2045;
        ELSIF x = 13773 THEN
            sigmoid_f := 2045;
        ELSIF x = 13774 THEN
            sigmoid_f := 2045;
        ELSIF x = 13775 THEN
            sigmoid_f := 2045;
        ELSIF x = 13776 THEN
            sigmoid_f := 2045;
        ELSIF x = 13777 THEN
            sigmoid_f := 2045;
        ELSIF x = 13778 THEN
            sigmoid_f := 2045;
        ELSIF x = 13779 THEN
            sigmoid_f := 2045;
        ELSIF x = 13780 THEN
            sigmoid_f := 2045;
        ELSIF x = 13781 THEN
            sigmoid_f := 2045;
        ELSIF x = 13782 THEN
            sigmoid_f := 2045;
        ELSIF x = 13783 THEN
            sigmoid_f := 2045;
        ELSIF x = 13784 THEN
            sigmoid_f := 2045;
        ELSIF x = 13785 THEN
            sigmoid_f := 2045;
        ELSIF x = 13786 THEN
            sigmoid_f := 2045;
        ELSIF x = 13787 THEN
            sigmoid_f := 2045;
        ELSIF x = 13788 THEN
            sigmoid_f := 2045;
        ELSIF x = 13789 THEN
            sigmoid_f := 2045;
        ELSIF x = 13790 THEN
            sigmoid_f := 2045;
        ELSIF x = 13791 THEN
            sigmoid_f := 2045;
        ELSIF x = 13792 THEN
            sigmoid_f := 2045;
        ELSIF x = 13793 THEN
            sigmoid_f := 2045;
        ELSIF x = 13794 THEN
            sigmoid_f := 2045;
        ELSIF x = 13795 THEN
            sigmoid_f := 2045;
        ELSIF x = 13796 THEN
            sigmoid_f := 2045;
        ELSIF x = 13797 THEN
            sigmoid_f := 2045;
        ELSIF x = 13798 THEN
            sigmoid_f := 2045;
        ELSIF x = 13799 THEN
            sigmoid_f := 2045;
        ELSIF x = 13800 THEN
            sigmoid_f := 2045;
        ELSIF x = 13801 THEN
            sigmoid_f := 2045;
        ELSIF x = 13802 THEN
            sigmoid_f := 2045;
        ELSIF x = 13803 THEN
            sigmoid_f := 2045;
        ELSIF x = 13804 THEN
            sigmoid_f := 2045;
        ELSIF x = 13805 THEN
            sigmoid_f := 2045;
        ELSIF x = 13806 THEN
            sigmoid_f := 2045;
        ELSIF x = 13807 THEN
            sigmoid_f := 2045;
        ELSIF x = 13808 THEN
            sigmoid_f := 2045;
        ELSIF x = 13809 THEN
            sigmoid_f := 2045;
        ELSIF x = 13810 THEN
            sigmoid_f := 2045;
        ELSIF x = 13811 THEN
            sigmoid_f := 2045;
        ELSIF x = 13812 THEN
            sigmoid_f := 2045;
        ELSIF x = 13813 THEN
            sigmoid_f := 2045;
        ELSIF x = 13814 THEN
            sigmoid_f := 2045;
        ELSIF x = 13815 THEN
            sigmoid_f := 2045;
        ELSIF x = 13816 THEN
            sigmoid_f := 2045;
        ELSIF x = 13817 THEN
            sigmoid_f := 2045;
        ELSIF x = 13818 THEN
            sigmoid_f := 2045;
        ELSIF x = 13819 THEN
            sigmoid_f := 2045;
        ELSIF x = 13820 THEN
            sigmoid_f := 2045;
        ELSIF x = 13821 THEN
            sigmoid_f := 2045;
        ELSIF x = 13822 THEN
            sigmoid_f := 2045;
        ELSIF x = 13823 THEN
            sigmoid_f := 2045;
        ELSIF x = 13824 THEN
            sigmoid_f := 2046;
        ELSIF x = 13825 THEN
            sigmoid_f := 2046;
        ELSIF x = 13826 THEN
            sigmoid_f := 2046;
        ELSIF x = 13827 THEN
            sigmoid_f := 2046;
        ELSIF x = 13828 THEN
            sigmoid_f := 2046;
        ELSIF x = 13829 THEN
            sigmoid_f := 2046;
        ELSIF x = 13830 THEN
            sigmoid_f := 2046;
        ELSIF x = 13831 THEN
            sigmoid_f := 2046;
        ELSIF x = 13832 THEN
            sigmoid_f := 2046;
        ELSIF x = 13833 THEN
            sigmoid_f := 2046;
        ELSIF x = 13834 THEN
            sigmoid_f := 2046;
        ELSIF x = 13835 THEN
            sigmoid_f := 2046;
        ELSIF x = 13836 THEN
            sigmoid_f := 2046;
        ELSIF x = 13837 THEN
            sigmoid_f := 2046;
        ELSIF x = 13838 THEN
            sigmoid_f := 2046;
        ELSIF x = 13839 THEN
            sigmoid_f := 2046;
        ELSIF x = 13840 THEN
            sigmoid_f := 2046;
        ELSIF x = 13841 THEN
            sigmoid_f := 2046;
        ELSIF x = 13842 THEN
            sigmoid_f := 2046;
        ELSIF x = 13843 THEN
            sigmoid_f := 2046;
        ELSIF x = 13844 THEN
            sigmoid_f := 2046;
        ELSIF x = 13845 THEN
            sigmoid_f := 2046;
        ELSIF x = 13846 THEN
            sigmoid_f := 2046;
        ELSIF x = 13847 THEN
            sigmoid_f := 2046;
        ELSIF x = 13848 THEN
            sigmoid_f := 2046;
        ELSIF x = 13849 THEN
            sigmoid_f := 2046;
        ELSIF x = 13850 THEN
            sigmoid_f := 2046;
        ELSIF x = 13851 THEN
            sigmoid_f := 2046;
        ELSIF x = 13852 THEN
            sigmoid_f := 2046;
        ELSIF x = 13853 THEN
            sigmoid_f := 2046;
        ELSIF x = 13854 THEN
            sigmoid_f := 2046;
        ELSIF x = 13855 THEN
            sigmoid_f := 2046;
        ELSIF x = 13856 THEN
            sigmoid_f := 2046;
        ELSIF x = 13857 THEN
            sigmoid_f := 2046;
        ELSIF x = 13858 THEN
            sigmoid_f := 2046;
        ELSIF x = 13859 THEN
            sigmoid_f := 2046;
        ELSIF x = 13860 THEN
            sigmoid_f := 2046;
        ELSIF x = 13861 THEN
            sigmoid_f := 2046;
        ELSIF x = 13862 THEN
            sigmoid_f := 2046;
        ELSIF x = 13863 THEN
            sigmoid_f := 2046;
        ELSIF x = 13864 THEN
            sigmoid_f := 2046;
        ELSIF x = 13865 THEN
            sigmoid_f := 2046;
        ELSIF x = 13866 THEN
            sigmoid_f := 2046;
        ELSIF x = 13867 THEN
            sigmoid_f := 2046;
        ELSIF x = 13868 THEN
            sigmoid_f := 2046;
        ELSIF x = 13869 THEN
            sigmoid_f := 2046;
        ELSIF x = 13870 THEN
            sigmoid_f := 2046;
        ELSIF x = 13871 THEN
            sigmoid_f := 2046;
        ELSIF x = 13872 THEN
            sigmoid_f := 2046;
        ELSIF x = 13873 THEN
            sigmoid_f := 2046;
        ELSIF x = 13874 THEN
            sigmoid_f := 2046;
        ELSIF x = 13875 THEN
            sigmoid_f := 2046;
        ELSIF x = 13876 THEN
            sigmoid_f := 2046;
        ELSIF x = 13877 THEN
            sigmoid_f := 2046;
        ELSIF x = 13878 THEN
            sigmoid_f := 2046;
        ELSIF x = 13879 THEN
            sigmoid_f := 2046;
        ELSIF x = 13880 THEN
            sigmoid_f := 2046;
        ELSIF x = 13881 THEN
            sigmoid_f := 2046;
        ELSIF x = 13882 THEN
            sigmoid_f := 2046;
        ELSIF x = 13883 THEN
            sigmoid_f := 2046;
        ELSIF x = 13884 THEN
            sigmoid_f := 2046;
        ELSIF x = 13885 THEN
            sigmoid_f := 2046;
        ELSIF x = 13886 THEN
            sigmoid_f := 2046;
        ELSIF x = 13887 THEN
            sigmoid_f := 2046;
        ELSIF x = 13888 THEN
            sigmoid_f := 2046;
        ELSIF x = 13889 THEN
            sigmoid_f := 2046;
        ELSIF x = 13890 THEN
            sigmoid_f := 2046;
        ELSIF x = 13891 THEN
            sigmoid_f := 2046;
        ELSIF x = 13892 THEN
            sigmoid_f := 2046;
        ELSIF x = 13893 THEN
            sigmoid_f := 2046;
        ELSIF x = 13894 THEN
            sigmoid_f := 2046;
        ELSIF x = 13895 THEN
            sigmoid_f := 2046;
        ELSIF x = 13896 THEN
            sigmoid_f := 2046;
        ELSIF x = 13897 THEN
            sigmoid_f := 2046;
        ELSIF x = 13898 THEN
            sigmoid_f := 2046;
        ELSIF x = 13899 THEN
            sigmoid_f := 2046;
        ELSIF x = 13900 THEN
            sigmoid_f := 2046;
        ELSIF x = 13901 THEN
            sigmoid_f := 2046;
        ELSIF x = 13902 THEN
            sigmoid_f := 2046;
        ELSIF x = 13903 THEN
            sigmoid_f := 2046;
        ELSIF x = 13904 THEN
            sigmoid_f := 2046;
        ELSIF x = 13905 THEN
            sigmoid_f := 2046;
        ELSIF x = 13906 THEN
            sigmoid_f := 2046;
        ELSIF x = 13907 THEN
            sigmoid_f := 2046;
        ELSIF x = 13908 THEN
            sigmoid_f := 2046;
        ELSIF x = 13909 THEN
            sigmoid_f := 2046;
        ELSIF x = 13910 THEN
            sigmoid_f := 2046;
        ELSIF x = 13911 THEN
            sigmoid_f := 2046;
        ELSIF x = 13912 THEN
            sigmoid_f := 2046;
        ELSIF x = 13913 THEN
            sigmoid_f := 2046;
        ELSIF x = 13914 THEN
            sigmoid_f := 2046;
        ELSIF x = 13915 THEN
            sigmoid_f := 2046;
        ELSIF x = 13916 THEN
            sigmoid_f := 2046;
        ELSIF x = 13917 THEN
            sigmoid_f := 2046;
        ELSIF x = 13918 THEN
            sigmoid_f := 2046;
        ELSIF x = 13919 THEN
            sigmoid_f := 2046;
        ELSIF x = 13920 THEN
            sigmoid_f := 2046;
        ELSIF x = 13921 THEN
            sigmoid_f := 2046;
        ELSIF x = 13922 THEN
            sigmoid_f := 2046;
        ELSIF x = 13923 THEN
            sigmoid_f := 2046;
        ELSIF x = 13924 THEN
            sigmoid_f := 2046;
        ELSIF x = 13925 THEN
            sigmoid_f := 2046;
        ELSIF x = 13926 THEN
            sigmoid_f := 2046;
        ELSIF x = 13927 THEN
            sigmoid_f := 2046;
        ELSIF x = 13928 THEN
            sigmoid_f := 2046;
        ELSIF x = 13929 THEN
            sigmoid_f := 2046;
        ELSIF x = 13930 THEN
            sigmoid_f := 2046;
        ELSIF x = 13931 THEN
            sigmoid_f := 2046;
        ELSIF x = 13932 THEN
            sigmoid_f := 2046;
        ELSIF x = 13933 THEN
            sigmoid_f := 2046;
        ELSIF x = 13934 THEN
            sigmoid_f := 2046;
        ELSIF x = 13935 THEN
            sigmoid_f := 2046;
        ELSIF x = 13936 THEN
            sigmoid_f := 2046;
        ELSIF x = 13937 THEN
            sigmoid_f := 2046;
        ELSIF x = 13938 THEN
            sigmoid_f := 2046;
        ELSIF x = 13939 THEN
            sigmoid_f := 2046;
        ELSIF x = 13940 THEN
            sigmoid_f := 2046;
        ELSIF x = 13941 THEN
            sigmoid_f := 2046;
        ELSIF x = 13942 THEN
            sigmoid_f := 2046;
        ELSIF x = 13943 THEN
            sigmoid_f := 2046;
        ELSIF x = 13944 THEN
            sigmoid_f := 2046;
        ELSIF x = 13945 THEN
            sigmoid_f := 2046;
        ELSIF x = 13946 THEN
            sigmoid_f := 2046;
        ELSIF x = 13947 THEN
            sigmoid_f := 2046;
        ELSIF x = 13948 THEN
            sigmoid_f := 2046;
        ELSIF x = 13949 THEN
            sigmoid_f := 2046;
        ELSIF x = 13950 THEN
            sigmoid_f := 2046;
        ELSIF x = 13951 THEN
            sigmoid_f := 2046;
        ELSIF x = 13952 THEN
            sigmoid_f := 2046;
        ELSIF x = 13953 THEN
            sigmoid_f := 2046;
        ELSIF x = 13954 THEN
            sigmoid_f := 2046;
        ELSIF x = 13955 THEN
            sigmoid_f := 2046;
        ELSIF x = 13956 THEN
            sigmoid_f := 2046;
        ELSIF x = 13957 THEN
            sigmoid_f := 2046;
        ELSIF x = 13958 THEN
            sigmoid_f := 2046;
        ELSIF x = 13959 THEN
            sigmoid_f := 2046;
        ELSIF x = 13960 THEN
            sigmoid_f := 2046;
        ELSIF x = 13961 THEN
            sigmoid_f := 2046;
        ELSIF x = 13962 THEN
            sigmoid_f := 2046;
        ELSIF x = 13963 THEN
            sigmoid_f := 2046;
        ELSIF x = 13964 THEN
            sigmoid_f := 2046;
        ELSIF x = 13965 THEN
            sigmoid_f := 2046;
        ELSIF x = 13966 THEN
            sigmoid_f := 2046;
        ELSIF x = 13967 THEN
            sigmoid_f := 2046;
        ELSIF x = 13968 THEN
            sigmoid_f := 2046;
        ELSIF x = 13969 THEN
            sigmoid_f := 2046;
        ELSIF x = 13970 THEN
            sigmoid_f := 2046;
        ELSIF x = 13971 THEN
            sigmoid_f := 2046;
        ELSIF x = 13972 THEN
            sigmoid_f := 2046;
        ELSIF x = 13973 THEN
            sigmoid_f := 2046;
        ELSIF x = 13974 THEN
            sigmoid_f := 2046;
        ELSIF x = 13975 THEN
            sigmoid_f := 2046;
        ELSIF x = 13976 THEN
            sigmoid_f := 2046;
        ELSIF x = 13977 THEN
            sigmoid_f := 2046;
        ELSIF x = 13978 THEN
            sigmoid_f := 2046;
        ELSIF x = 13979 THEN
            sigmoid_f := 2046;
        ELSIF x = 13980 THEN
            sigmoid_f := 2046;
        ELSIF x = 13981 THEN
            sigmoid_f := 2046;
        ELSIF x = 13982 THEN
            sigmoid_f := 2046;
        ELSIF x = 13983 THEN
            sigmoid_f := 2046;
        ELSIF x = 13984 THEN
            sigmoid_f := 2046;
        ELSIF x = 13985 THEN
            sigmoid_f := 2046;
        ELSIF x = 13986 THEN
            sigmoid_f := 2046;
        ELSIF x = 13987 THEN
            sigmoid_f := 2046;
        ELSIF x = 13988 THEN
            sigmoid_f := 2046;
        ELSIF x = 13989 THEN
            sigmoid_f := 2046;
        ELSIF x = 13990 THEN
            sigmoid_f := 2046;
        ELSIF x = 13991 THEN
            sigmoid_f := 2046;
        ELSIF x = 13992 THEN
            sigmoid_f := 2046;
        ELSIF x = 13993 THEN
            sigmoid_f := 2046;
        ELSIF x = 13994 THEN
            sigmoid_f := 2046;
        ELSIF x = 13995 THEN
            sigmoid_f := 2046;
        ELSIF x = 13996 THEN
            sigmoid_f := 2046;
        ELSIF x = 13997 THEN
            sigmoid_f := 2046;
        ELSIF x = 13998 THEN
            sigmoid_f := 2046;
        ELSIF x = 13999 THEN
            sigmoid_f := 2046;
        ELSIF x = 14000 THEN
            sigmoid_f := 2046;
        ELSIF x = 14001 THEN
            sigmoid_f := 2046;
        ELSIF x = 14002 THEN
            sigmoid_f := 2046;
        ELSIF x = 14003 THEN
            sigmoid_f := 2046;
        ELSIF x = 14004 THEN
            sigmoid_f := 2046;
        ELSIF x = 14005 THEN
            sigmoid_f := 2046;
        ELSIF x = 14006 THEN
            sigmoid_f := 2046;
        ELSIF x = 14007 THEN
            sigmoid_f := 2046;
        ELSIF x = 14008 THEN
            sigmoid_f := 2046;
        ELSIF x = 14009 THEN
            sigmoid_f := 2046;
        ELSIF x = 14010 THEN
            sigmoid_f := 2046;
        ELSIF x = 14011 THEN
            sigmoid_f := 2046;
        ELSIF x = 14012 THEN
            sigmoid_f := 2046;
        ELSIF x = 14013 THEN
            sigmoid_f := 2046;
        ELSIF x = 14014 THEN
            sigmoid_f := 2046;
        ELSIF x = 14015 THEN
            sigmoid_f := 2046;
        ELSIF x = 14016 THEN
            sigmoid_f := 2046;
        ELSIF x = 14017 THEN
            sigmoid_f := 2046;
        ELSIF x = 14018 THEN
            sigmoid_f := 2046;
        ELSIF x = 14019 THEN
            sigmoid_f := 2046;
        ELSIF x = 14020 THEN
            sigmoid_f := 2046;
        ELSIF x = 14021 THEN
            sigmoid_f := 2046;
        ELSIF x = 14022 THEN
            sigmoid_f := 2046;
        ELSIF x = 14023 THEN
            sigmoid_f := 2046;
        ELSIF x = 14024 THEN
            sigmoid_f := 2046;
        ELSIF x = 14025 THEN
            sigmoid_f := 2046;
        ELSIF x = 14026 THEN
            sigmoid_f := 2046;
        ELSIF x = 14027 THEN
            sigmoid_f := 2046;
        ELSIF x = 14028 THEN
            sigmoid_f := 2046;
        ELSIF x = 14029 THEN
            sigmoid_f := 2046;
        ELSIF x = 14030 THEN
            sigmoid_f := 2046;
        ELSIF x = 14031 THEN
            sigmoid_f := 2046;
        ELSIF x = 14032 THEN
            sigmoid_f := 2046;
        ELSIF x = 14033 THEN
            sigmoid_f := 2046;
        ELSIF x = 14034 THEN
            sigmoid_f := 2046;
        ELSIF x = 14035 THEN
            sigmoid_f := 2046;
        ELSIF x = 14036 THEN
            sigmoid_f := 2046;
        ELSIF x = 14037 THEN
            sigmoid_f := 2046;
        ELSIF x = 14038 THEN
            sigmoid_f := 2046;
        ELSIF x = 14039 THEN
            sigmoid_f := 2046;
        ELSIF x = 14040 THEN
            sigmoid_f := 2046;
        ELSIF x = 14041 THEN
            sigmoid_f := 2046;
        ELSIF x = 14042 THEN
            sigmoid_f := 2046;
        ELSIF x = 14043 THEN
            sigmoid_f := 2046;
        ELSIF x = 14044 THEN
            sigmoid_f := 2046;
        ELSIF x = 14045 THEN
            sigmoid_f := 2046;
        ELSIF x = 14046 THEN
            sigmoid_f := 2046;
        ELSIF x = 14047 THEN
            sigmoid_f := 2046;
        ELSIF x = 14048 THEN
            sigmoid_f := 2046;
        ELSIF x = 14049 THEN
            sigmoid_f := 2046;
        ELSIF x = 14050 THEN
            sigmoid_f := 2046;
        ELSIF x = 14051 THEN
            sigmoid_f := 2046;
        ELSIF x = 14052 THEN
            sigmoid_f := 2046;
        ELSIF x = 14053 THEN
            sigmoid_f := 2046;
        ELSIF x = 14054 THEN
            sigmoid_f := 2046;
        ELSIF x = 14055 THEN
            sigmoid_f := 2046;
        ELSIF x = 14056 THEN
            sigmoid_f := 2046;
        ELSIF x = 14057 THEN
            sigmoid_f := 2046;
        ELSIF x = 14058 THEN
            sigmoid_f := 2046;
        ELSIF x = 14059 THEN
            sigmoid_f := 2046;
        ELSIF x = 14060 THEN
            sigmoid_f := 2046;
        ELSIF x = 14061 THEN
            sigmoid_f := 2046;
        ELSIF x = 14062 THEN
            sigmoid_f := 2046;
        ELSIF x = 14063 THEN
            sigmoid_f := 2046;
        ELSIF x = 14064 THEN
            sigmoid_f := 2046;
        ELSIF x = 14065 THEN
            sigmoid_f := 2046;
        ELSIF x = 14066 THEN
            sigmoid_f := 2046;
        ELSIF x = 14067 THEN
            sigmoid_f := 2046;
        ELSIF x = 14068 THEN
            sigmoid_f := 2046;
        ELSIF x = 14069 THEN
            sigmoid_f := 2046;
        ELSIF x = 14070 THEN
            sigmoid_f := 2046;
        ELSIF x = 14071 THEN
            sigmoid_f := 2046;
        ELSIF x = 14072 THEN
            sigmoid_f := 2046;
        ELSIF x = 14073 THEN
            sigmoid_f := 2046;
        ELSIF x = 14074 THEN
            sigmoid_f := 2046;
        ELSIF x = 14075 THEN
            sigmoid_f := 2046;
        ELSIF x = 14076 THEN
            sigmoid_f := 2046;
        ELSIF x = 14077 THEN
            sigmoid_f := 2046;
        ELSIF x = 14078 THEN
            sigmoid_f := 2046;
        ELSIF x = 14079 THEN
            sigmoid_f := 2046;
        ELSIF x = 14080 THEN
            sigmoid_f := 2046;
        ELSIF x = 14081 THEN
            sigmoid_f := 2046;
        ELSIF x = 14082 THEN
            sigmoid_f := 2046;
        ELSIF x = 14083 THEN
            sigmoid_f := 2046;
        ELSIF x = 14084 THEN
            sigmoid_f := 2046;
        ELSIF x = 14085 THEN
            sigmoid_f := 2046;
        ELSIF x = 14086 THEN
            sigmoid_f := 2046;
        ELSIF x = 14087 THEN
            sigmoid_f := 2046;
        ELSIF x = 14088 THEN
            sigmoid_f := 2046;
        ELSIF x = 14089 THEN
            sigmoid_f := 2046;
        ELSIF x = 14090 THEN
            sigmoid_f := 2046;
        ELSIF x = 14091 THEN
            sigmoid_f := 2046;
        ELSIF x = 14092 THEN
            sigmoid_f := 2046;
        ELSIF x = 14093 THEN
            sigmoid_f := 2046;
        ELSIF x = 14094 THEN
            sigmoid_f := 2046;
        ELSIF x = 14095 THEN
            sigmoid_f := 2046;
        ELSIF x = 14096 THEN
            sigmoid_f := 2046;
        ELSIF x = 14097 THEN
            sigmoid_f := 2046;
        ELSIF x = 14098 THEN
            sigmoid_f := 2046;
        ELSIF x = 14099 THEN
            sigmoid_f := 2046;
        ELSIF x = 14100 THEN
            sigmoid_f := 2046;
        ELSIF x = 14101 THEN
            sigmoid_f := 2046;
        ELSIF x = 14102 THEN
            sigmoid_f := 2046;
        ELSIF x = 14103 THEN
            sigmoid_f := 2046;
        ELSIF x = 14104 THEN
            sigmoid_f := 2046;
        ELSIF x = 14105 THEN
            sigmoid_f := 2046;
        ELSIF x = 14106 THEN
            sigmoid_f := 2046;
        ELSIF x = 14107 THEN
            sigmoid_f := 2046;
        ELSIF x = 14108 THEN
            sigmoid_f := 2046;
        ELSIF x = 14109 THEN
            sigmoid_f := 2046;
        ELSIF x = 14110 THEN
            sigmoid_f := 2046;
        ELSIF x = 14111 THEN
            sigmoid_f := 2046;
        ELSIF x = 14112 THEN
            sigmoid_f := 2046;
        ELSIF x = 14113 THEN
            sigmoid_f := 2046;
        ELSIF x = 14114 THEN
            sigmoid_f := 2046;
        ELSIF x = 14115 THEN
            sigmoid_f := 2046;
        ELSIF x = 14116 THEN
            sigmoid_f := 2046;
        ELSIF x = 14117 THEN
            sigmoid_f := 2046;
        ELSIF x = 14118 THEN
            sigmoid_f := 2046;
        ELSIF x = 14119 THEN
            sigmoid_f := 2046;
        ELSIF x = 14120 THEN
            sigmoid_f := 2046;
        ELSIF x = 14121 THEN
            sigmoid_f := 2046;
        ELSIF x = 14122 THEN
            sigmoid_f := 2046;
        ELSIF x = 14123 THEN
            sigmoid_f := 2046;
        ELSIF x = 14124 THEN
            sigmoid_f := 2046;
        ELSIF x = 14125 THEN
            sigmoid_f := 2046;
        ELSIF x = 14126 THEN
            sigmoid_f := 2046;
        ELSIF x = 14127 THEN
            sigmoid_f := 2046;
        ELSIF x = 14128 THEN
            sigmoid_f := 2046;
        ELSIF x = 14129 THEN
            sigmoid_f := 2046;
        ELSIF x = 14130 THEN
            sigmoid_f := 2046;
        ELSIF x = 14131 THEN
            sigmoid_f := 2046;
        ELSIF x = 14132 THEN
            sigmoid_f := 2046;
        ELSIF x = 14133 THEN
            sigmoid_f := 2046;
        ELSIF x = 14134 THEN
            sigmoid_f := 2046;
        ELSIF x = 14135 THEN
            sigmoid_f := 2046;
        ELSIF x = 14136 THEN
            sigmoid_f := 2046;
        ELSIF x = 14137 THEN
            sigmoid_f := 2046;
        ELSIF x = 14138 THEN
            sigmoid_f := 2046;
        ELSIF x = 14139 THEN
            sigmoid_f := 2046;
        ELSIF x = 14140 THEN
            sigmoid_f := 2046;
        ELSIF x = 14141 THEN
            sigmoid_f := 2046;
        ELSIF x = 14142 THEN
            sigmoid_f := 2046;
        ELSIF x = 14143 THEN
            sigmoid_f := 2046;
        ELSIF x = 14144 THEN
            sigmoid_f := 2046;
        ELSIF x = 14145 THEN
            sigmoid_f := 2046;
        ELSIF x = 14146 THEN
            sigmoid_f := 2046;
        ELSIF x = 14147 THEN
            sigmoid_f := 2046;
        ELSIF x = 14148 THEN
            sigmoid_f := 2046;
        ELSIF x = 14149 THEN
            sigmoid_f := 2046;
        ELSIF x = 14150 THEN
            sigmoid_f := 2046;
        ELSIF x = 14151 THEN
            sigmoid_f := 2046;
        ELSIF x = 14152 THEN
            sigmoid_f := 2046;
        ELSIF x = 14153 THEN
            sigmoid_f := 2046;
        ELSIF x = 14154 THEN
            sigmoid_f := 2046;
        ELSIF x = 14155 THEN
            sigmoid_f := 2046;
        ELSIF x = 14156 THEN
            sigmoid_f := 2046;
        ELSIF x = 14157 THEN
            sigmoid_f := 2046;
        ELSIF x = 14158 THEN
            sigmoid_f := 2046;
        ELSIF x = 14159 THEN
            sigmoid_f := 2046;
        ELSIF x = 14160 THEN
            sigmoid_f := 2046;
        ELSIF x = 14161 THEN
            sigmoid_f := 2046;
        ELSIF x = 14162 THEN
            sigmoid_f := 2046;
        ELSIF x = 14163 THEN
            sigmoid_f := 2046;
        ELSIF x = 14164 THEN
            sigmoid_f := 2046;
        ELSIF x = 14165 THEN
            sigmoid_f := 2046;
        ELSIF x = 14166 THEN
            sigmoid_f := 2046;
        ELSIF x = 14167 THEN
            sigmoid_f := 2046;
        ELSIF x = 14168 THEN
            sigmoid_f := 2046;
        ELSIF x = 14169 THEN
            sigmoid_f := 2046;
        ELSIF x = 14170 THEN
            sigmoid_f := 2046;
        ELSIF x = 14171 THEN
            sigmoid_f := 2046;
        ELSIF x = 14172 THEN
            sigmoid_f := 2046;
        ELSIF x = 14173 THEN
            sigmoid_f := 2046;
        ELSIF x = 14174 THEN
            sigmoid_f := 2046;
        ELSIF x = 14175 THEN
            sigmoid_f := 2046;
        ELSIF x = 14176 THEN
            sigmoid_f := 2046;
        ELSIF x = 14177 THEN
            sigmoid_f := 2046;
        ELSIF x = 14178 THEN
            sigmoid_f := 2046;
        ELSIF x = 14179 THEN
            sigmoid_f := 2046;
        ELSIF x = 14180 THEN
            sigmoid_f := 2046;
        ELSIF x = 14181 THEN
            sigmoid_f := 2046;
        ELSIF x = 14182 THEN
            sigmoid_f := 2046;
        ELSIF x = 14183 THEN
            sigmoid_f := 2046;
        ELSIF x = 14184 THEN
            sigmoid_f := 2046;
        ELSIF x = 14185 THEN
            sigmoid_f := 2046;
        ELSIF x = 14186 THEN
            sigmoid_f := 2046;
        ELSIF x = 14187 THEN
            sigmoid_f := 2046;
        ELSIF x = 14188 THEN
            sigmoid_f := 2046;
        ELSIF x = 14189 THEN
            sigmoid_f := 2046;
        ELSIF x = 14190 THEN
            sigmoid_f := 2046;
        ELSIF x = 14191 THEN
            sigmoid_f := 2046;
        ELSIF x = 14192 THEN
            sigmoid_f := 2046;
        ELSIF x = 14193 THEN
            sigmoid_f := 2046;
        ELSIF x = 14194 THEN
            sigmoid_f := 2046;
        ELSIF x = 14195 THEN
            sigmoid_f := 2046;
        ELSIF x = 14196 THEN
            sigmoid_f := 2046;
        ELSIF x = 14197 THEN
            sigmoid_f := 2046;
        ELSIF x = 14198 THEN
            sigmoid_f := 2046;
        ELSIF x = 14199 THEN
            sigmoid_f := 2046;
        ELSIF x = 14200 THEN
            sigmoid_f := 2046;
        ELSIF x = 14201 THEN
            sigmoid_f := 2046;
        ELSIF x = 14202 THEN
            sigmoid_f := 2046;
        ELSIF x = 14203 THEN
            sigmoid_f := 2046;
        ELSIF x = 14204 THEN
            sigmoid_f := 2046;
        ELSIF x = 14205 THEN
            sigmoid_f := 2046;
        ELSIF x = 14206 THEN
            sigmoid_f := 2046;
        ELSIF x = 14207 THEN
            sigmoid_f := 2046;
        ELSIF x = 14208 THEN
            sigmoid_f := 2046;
        ELSIF x = 14209 THEN
            sigmoid_f := 2046;
        ELSIF x = 14210 THEN
            sigmoid_f := 2046;
        ELSIF x = 14211 THEN
            sigmoid_f := 2046;
        ELSIF x = 14212 THEN
            sigmoid_f := 2046;
        ELSIF x = 14213 THEN
            sigmoid_f := 2046;
        ELSIF x = 14214 THEN
            sigmoid_f := 2046;
        ELSIF x = 14215 THEN
            sigmoid_f := 2046;
        ELSIF x = 14216 THEN
            sigmoid_f := 2046;
        ELSIF x = 14217 THEN
            sigmoid_f := 2046;
        ELSIF x = 14218 THEN
            sigmoid_f := 2046;
        ELSIF x = 14219 THEN
            sigmoid_f := 2046;
        ELSIF x = 14220 THEN
            sigmoid_f := 2046;
        ELSIF x = 14221 THEN
            sigmoid_f := 2046;
        ELSIF x = 14222 THEN
            sigmoid_f := 2046;
        ELSIF x = 14223 THEN
            sigmoid_f := 2046;
        ELSIF x = 14224 THEN
            sigmoid_f := 2046;
        ELSIF x = 14225 THEN
            sigmoid_f := 2046;
        ELSIF x = 14226 THEN
            sigmoid_f := 2046;
        ELSIF x = 14227 THEN
            sigmoid_f := 2046;
        ELSIF x = 14228 THEN
            sigmoid_f := 2046;
        ELSIF x = 14229 THEN
            sigmoid_f := 2046;
        ELSIF x = 14230 THEN
            sigmoid_f := 2046;
        ELSIF x = 14231 THEN
            sigmoid_f := 2046;
        ELSIF x = 14232 THEN
            sigmoid_f := 2046;
        ELSIF x = 14233 THEN
            sigmoid_f := 2046;
        ELSIF x = 14234 THEN
            sigmoid_f := 2046;
        ELSIF x = 14235 THEN
            sigmoid_f := 2046;
        ELSIF x = 14236 THEN
            sigmoid_f := 2046;
        ELSIF x = 14237 THEN
            sigmoid_f := 2046;
        ELSIF x = 14238 THEN
            sigmoid_f := 2046;
        ELSIF x = 14239 THEN
            sigmoid_f := 2046;
        ELSIF x = 14240 THEN
            sigmoid_f := 2046;
        ELSIF x = 14241 THEN
            sigmoid_f := 2046;
        ELSIF x = 14242 THEN
            sigmoid_f := 2046;
        ELSIF x = 14243 THEN
            sigmoid_f := 2046;
        ELSIF x = 14244 THEN
            sigmoid_f := 2046;
        ELSIF x = 14245 THEN
            sigmoid_f := 2046;
        ELSIF x = 14246 THEN
            sigmoid_f := 2046;
        ELSIF x = 14247 THEN
            sigmoid_f := 2046;
        ELSIF x = 14248 THEN
            sigmoid_f := 2046;
        ELSIF x = 14249 THEN
            sigmoid_f := 2046;
        ELSIF x = 14250 THEN
            sigmoid_f := 2046;
        ELSIF x = 14251 THEN
            sigmoid_f := 2046;
        ELSIF x = 14252 THEN
            sigmoid_f := 2046;
        ELSIF x = 14253 THEN
            sigmoid_f := 2046;
        ELSIF x = 14254 THEN
            sigmoid_f := 2046;
        ELSIF x = 14255 THEN
            sigmoid_f := 2046;
        ELSIF x = 14256 THEN
            sigmoid_f := 2046;
        ELSIF x = 14257 THEN
            sigmoid_f := 2046;
        ELSIF x = 14258 THEN
            sigmoid_f := 2046;
        ELSIF x = 14259 THEN
            sigmoid_f := 2046;
        ELSIF x = 14260 THEN
            sigmoid_f := 2046;
        ELSIF x = 14261 THEN
            sigmoid_f := 2046;
        ELSIF x = 14262 THEN
            sigmoid_f := 2046;
        ELSIF x = 14263 THEN
            sigmoid_f := 2046;
        ELSIF x = 14264 THEN
            sigmoid_f := 2046;
        ELSIF x = 14265 THEN
            sigmoid_f := 2046;
        ELSIF x = 14266 THEN
            sigmoid_f := 2046;
        ELSIF x = 14267 THEN
            sigmoid_f := 2046;
        ELSIF x = 14268 THEN
            sigmoid_f := 2046;
        ELSIF x = 14269 THEN
            sigmoid_f := 2046;
        ELSIF x = 14270 THEN
            sigmoid_f := 2046;
        ELSIF x = 14271 THEN
            sigmoid_f := 2046;
        ELSIF x = 14272 THEN
            sigmoid_f := 2046;
        ELSIF x = 14273 THEN
            sigmoid_f := 2046;
        ELSIF x = 14274 THEN
            sigmoid_f := 2046;
        ELSIF x = 14275 THEN
            sigmoid_f := 2046;
        ELSIF x = 14276 THEN
            sigmoid_f := 2046;
        ELSIF x = 14277 THEN
            sigmoid_f := 2046;
        ELSIF x = 14278 THEN
            sigmoid_f := 2046;
        ELSIF x = 14279 THEN
            sigmoid_f := 2046;
        ELSIF x = 14280 THEN
            sigmoid_f := 2046;
        ELSIF x = 14281 THEN
            sigmoid_f := 2046;
        ELSIF x = 14282 THEN
            sigmoid_f := 2046;
        ELSIF x = 14283 THEN
            sigmoid_f := 2046;
        ELSIF x = 14284 THEN
            sigmoid_f := 2046;
        ELSIF x = 14285 THEN
            sigmoid_f := 2046;
        ELSIF x = 14286 THEN
            sigmoid_f := 2046;
        ELSIF x = 14287 THEN
            sigmoid_f := 2046;
        ELSIF x = 14288 THEN
            sigmoid_f := 2046;
        ELSIF x = 14289 THEN
            sigmoid_f := 2046;
        ELSIF x = 14290 THEN
            sigmoid_f := 2046;
        ELSIF x = 14291 THEN
            sigmoid_f := 2046;
        ELSIF x = 14292 THEN
            sigmoid_f := 2046;
        ELSIF x = 14293 THEN
            sigmoid_f := 2046;
        ELSIF x = 14294 THEN
            sigmoid_f := 2046;
        ELSIF x = 14295 THEN
            sigmoid_f := 2046;
        ELSIF x = 14296 THEN
            sigmoid_f := 2046;
        ELSIF x = 14297 THEN
            sigmoid_f := 2046;
        ELSIF x = 14298 THEN
            sigmoid_f := 2046;
        ELSIF x = 14299 THEN
            sigmoid_f := 2046;
        ELSIF x = 14300 THEN
            sigmoid_f := 2046;
        ELSIF x = 14301 THEN
            sigmoid_f := 2046;
        ELSIF x = 14302 THEN
            sigmoid_f := 2046;
        ELSIF x = 14303 THEN
            sigmoid_f := 2046;
        ELSIF x = 14304 THEN
            sigmoid_f := 2046;
        ELSIF x = 14305 THEN
            sigmoid_f := 2046;
        ELSIF x = 14306 THEN
            sigmoid_f := 2046;
        ELSIF x = 14307 THEN
            sigmoid_f := 2046;
        ELSIF x = 14308 THEN
            sigmoid_f := 2046;
        ELSIF x = 14309 THEN
            sigmoid_f := 2046;
        ELSIF x = 14310 THEN
            sigmoid_f := 2046;
        ELSIF x = 14311 THEN
            sigmoid_f := 2046;
        ELSIF x = 14312 THEN
            sigmoid_f := 2046;
        ELSIF x = 14313 THEN
            sigmoid_f := 2046;
        ELSIF x = 14314 THEN
            sigmoid_f := 2046;
        ELSIF x = 14315 THEN
            sigmoid_f := 2046;
        ELSIF x = 14316 THEN
            sigmoid_f := 2046;
        ELSIF x = 14317 THEN
            sigmoid_f := 2046;
        ELSIF x = 14318 THEN
            sigmoid_f := 2046;
        ELSIF x = 14319 THEN
            sigmoid_f := 2046;
        ELSIF x = 14320 THEN
            sigmoid_f := 2046;
        ELSIF x = 14321 THEN
            sigmoid_f := 2046;
        ELSIF x = 14322 THEN
            sigmoid_f := 2046;
        ELSIF x = 14323 THEN
            sigmoid_f := 2046;
        ELSIF x = 14324 THEN
            sigmoid_f := 2046;
        ELSIF x = 14325 THEN
            sigmoid_f := 2046;
        ELSIF x = 14326 THEN
            sigmoid_f := 2046;
        ELSIF x = 14327 THEN
            sigmoid_f := 2046;
        ELSIF x = 14328 THEN
            sigmoid_f := 2046;
        ELSIF x = 14329 THEN
            sigmoid_f := 2046;
        ELSIF x = 14330 THEN
            sigmoid_f := 2046;
        ELSIF x = 14331 THEN
            sigmoid_f := 2046;
        ELSIF x = 14332 THEN
            sigmoid_f := 2046;
        ELSIF x = 14333 THEN
            sigmoid_f := 2046;
        ELSIF x = 14334 THEN
            sigmoid_f := 2046;
        ELSIF x = 14335 THEN
            sigmoid_f := 2046;
        ELSIF x = 14336 THEN
            sigmoid_f := 2046;
        ELSIF x = 14337 THEN
            sigmoid_f := 2046;
        ELSIF x = 14338 THEN
            sigmoid_f := 2046;
        ELSIF x = 14339 THEN
            sigmoid_f := 2046;
        ELSIF x = 14340 THEN
            sigmoid_f := 2046;
        ELSIF x = 14341 THEN
            sigmoid_f := 2046;
        ELSIF x = 14342 THEN
            sigmoid_f := 2046;
        ELSIF x = 14343 THEN
            sigmoid_f := 2046;
        ELSIF x = 14344 THEN
            sigmoid_f := 2046;
        ELSIF x = 14345 THEN
            sigmoid_f := 2046;
        ELSIF x = 14346 THEN
            sigmoid_f := 2046;
        ELSIF x = 14347 THEN
            sigmoid_f := 2046;
        ELSIF x = 14348 THEN
            sigmoid_f := 2046;
        ELSIF x = 14349 THEN
            sigmoid_f := 2046;
        ELSIF x = 14350 THEN
            sigmoid_f := 2046;
        ELSIF x = 14351 THEN
            sigmoid_f := 2046;
        ELSIF x = 14352 THEN
            sigmoid_f := 2046;
        ELSIF x = 14353 THEN
            sigmoid_f := 2046;
        ELSIF x = 14354 THEN
            sigmoid_f := 2046;
        ELSIF x = 14355 THEN
            sigmoid_f := 2046;
        ELSIF x = 14356 THEN
            sigmoid_f := 2046;
        ELSIF x = 14357 THEN
            sigmoid_f := 2046;
        ELSIF x = 14358 THEN
            sigmoid_f := 2046;
        ELSIF x = 14359 THEN
            sigmoid_f := 2046;
        ELSIF x = 14360 THEN
            sigmoid_f := 2046;
        ELSIF x = 14361 THEN
            sigmoid_f := 2046;
        ELSIF x = 14362 THEN
            sigmoid_f := 2046;
        ELSIF x = 14363 THEN
            sigmoid_f := 2046;
        ELSIF x = 14364 THEN
            sigmoid_f := 2046;
        ELSIF x = 14365 THEN
            sigmoid_f := 2046;
        ELSIF x = 14366 THEN
            sigmoid_f := 2046;
        ELSIF x = 14367 THEN
            sigmoid_f := 2046;
        ELSIF x = 14368 THEN
            sigmoid_f := 2046;
        ELSIF x = 14369 THEN
            sigmoid_f := 2046;
        ELSIF x = 14370 THEN
            sigmoid_f := 2046;
        ELSIF x = 14371 THEN
            sigmoid_f := 2046;
        ELSIF x = 14372 THEN
            sigmoid_f := 2046;
        ELSIF x = 14373 THEN
            sigmoid_f := 2046;
        ELSIF x = 14374 THEN
            sigmoid_f := 2046;
        ELSIF x = 14375 THEN
            sigmoid_f := 2046;
        ELSIF x = 14376 THEN
            sigmoid_f := 2046;
        ELSIF x = 14377 THEN
            sigmoid_f := 2046;
        ELSIF x = 14378 THEN
            sigmoid_f := 2046;
        ELSIF x = 14379 THEN
            sigmoid_f := 2046;
        ELSIF x = 14380 THEN
            sigmoid_f := 2046;
        ELSIF x = 14381 THEN
            sigmoid_f := 2046;
        ELSIF x = 14382 THEN
            sigmoid_f := 2046;
        ELSIF x = 14383 THEN
            sigmoid_f := 2046;
        ELSIF x = 14384 THEN
            sigmoid_f := 2046;
        ELSIF x = 14385 THEN
            sigmoid_f := 2046;
        ELSIF x = 14386 THEN
            sigmoid_f := 2046;
        ELSIF x = 14387 THEN
            sigmoid_f := 2046;
        ELSIF x = 14388 THEN
            sigmoid_f := 2046;
        ELSIF x = 14389 THEN
            sigmoid_f := 2046;
        ELSIF x = 14390 THEN
            sigmoid_f := 2046;
        ELSIF x = 14391 THEN
            sigmoid_f := 2046;
        ELSIF x = 14392 THEN
            sigmoid_f := 2046;
        ELSIF x = 14393 THEN
            sigmoid_f := 2046;
        ELSIF x = 14394 THEN
            sigmoid_f := 2046;
        ELSIF x = 14395 THEN
            sigmoid_f := 2046;
        ELSIF x = 14396 THEN
            sigmoid_f := 2046;
        ELSIF x = 14397 THEN
            sigmoid_f := 2046;
        ELSIF x = 14398 THEN
            sigmoid_f := 2046;
        ELSIF x = 14399 THEN
            sigmoid_f := 2046;
        ELSIF x = 14400 THEN
            sigmoid_f := 2046;
        ELSIF x = 14401 THEN
            sigmoid_f := 2046;
        ELSIF x = 14402 THEN
            sigmoid_f := 2046;
        ELSIF x = 14403 THEN
            sigmoid_f := 2046;
        ELSIF x = 14404 THEN
            sigmoid_f := 2046;
        ELSIF x = 14405 THEN
            sigmoid_f := 2046;
        ELSIF x = 14406 THEN
            sigmoid_f := 2046;
        ELSIF x = 14407 THEN
            sigmoid_f := 2046;
        ELSIF x = 14408 THEN
            sigmoid_f := 2046;
        ELSIF x = 14409 THEN
            sigmoid_f := 2046;
        ELSIF x = 14410 THEN
            sigmoid_f := 2046;
        ELSIF x = 14411 THEN
            sigmoid_f := 2046;
        ELSIF x = 14412 THEN
            sigmoid_f := 2046;
        ELSIF x = 14413 THEN
            sigmoid_f := 2046;
        ELSIF x = 14414 THEN
            sigmoid_f := 2046;
        ELSIF x = 14415 THEN
            sigmoid_f := 2046;
        ELSIF x = 14416 THEN
            sigmoid_f := 2046;
        ELSIF x = 14417 THEN
            sigmoid_f := 2046;
        ELSIF x = 14418 THEN
            sigmoid_f := 2046;
        ELSIF x = 14419 THEN
            sigmoid_f := 2046;
        ELSIF x = 14420 THEN
            sigmoid_f := 2046;
        ELSIF x = 14421 THEN
            sigmoid_f := 2046;
        ELSIF x = 14422 THEN
            sigmoid_f := 2046;
        ELSIF x = 14423 THEN
            sigmoid_f := 2046;
        ELSIF x = 14424 THEN
            sigmoid_f := 2046;
        ELSIF x = 14425 THEN
            sigmoid_f := 2046;
        ELSIF x = 14426 THEN
            sigmoid_f := 2046;
        ELSIF x = 14427 THEN
            sigmoid_f := 2046;
        ELSIF x = 14428 THEN
            sigmoid_f := 2046;
        ELSIF x = 14429 THEN
            sigmoid_f := 2046;
        ELSIF x = 14430 THEN
            sigmoid_f := 2046;
        ELSIF x = 14431 THEN
            sigmoid_f := 2046;
        ELSIF x = 14432 THEN
            sigmoid_f := 2046;
        ELSIF x = 14433 THEN
            sigmoid_f := 2046;
        ELSIF x = 14434 THEN
            sigmoid_f := 2046;
        ELSIF x = 14435 THEN
            sigmoid_f := 2046;
        ELSIF x = 14436 THEN
            sigmoid_f := 2046;
        ELSIF x = 14437 THEN
            sigmoid_f := 2046;
        ELSIF x = 14438 THEN
            sigmoid_f := 2046;
        ELSIF x = 14439 THEN
            sigmoid_f := 2046;
        ELSIF x = 14440 THEN
            sigmoid_f := 2046;
        ELSIF x = 14441 THEN
            sigmoid_f := 2046;
        ELSIF x = 14442 THEN
            sigmoid_f := 2046;
        ELSIF x = 14443 THEN
            sigmoid_f := 2046;
        ELSIF x = 14444 THEN
            sigmoid_f := 2046;
        ELSIF x = 14445 THEN
            sigmoid_f := 2046;
        ELSIF x = 14446 THEN
            sigmoid_f := 2046;
        ELSIF x = 14447 THEN
            sigmoid_f := 2046;
        ELSIF x = 14448 THEN
            sigmoid_f := 2046;
        ELSIF x = 14449 THEN
            sigmoid_f := 2046;
        ELSIF x = 14450 THEN
            sigmoid_f := 2046;
        ELSIF x = 14451 THEN
            sigmoid_f := 2046;
        ELSIF x = 14452 THEN
            sigmoid_f := 2046;
        ELSIF x = 14453 THEN
            sigmoid_f := 2046;
        ELSIF x = 14454 THEN
            sigmoid_f := 2046;
        ELSIF x = 14455 THEN
            sigmoid_f := 2046;
        ELSIF x = 14456 THEN
            sigmoid_f := 2046;
        ELSIF x = 14457 THEN
            sigmoid_f := 2046;
        ELSIF x = 14458 THEN
            sigmoid_f := 2046;
        ELSIF x = 14459 THEN
            sigmoid_f := 2046;
        ELSIF x = 14460 THEN
            sigmoid_f := 2046;
        ELSIF x = 14461 THEN
            sigmoid_f := 2046;
        ELSIF x = 14462 THEN
            sigmoid_f := 2046;
        ELSIF x = 14463 THEN
            sigmoid_f := 2046;
        ELSIF x = 14464 THEN
            sigmoid_f := 2046;
        ELSIF x = 14465 THEN
            sigmoid_f := 2046;
        ELSIF x = 14466 THEN
            sigmoid_f := 2046;
        ELSIF x = 14467 THEN
            sigmoid_f := 2046;
        ELSIF x = 14468 THEN
            sigmoid_f := 2046;
        ELSIF x = 14469 THEN
            sigmoid_f := 2046;
        ELSIF x = 14470 THEN
            sigmoid_f := 2046;
        ELSIF x = 14471 THEN
            sigmoid_f := 2046;
        ELSIF x = 14472 THEN
            sigmoid_f := 2046;
        ELSIF x = 14473 THEN
            sigmoid_f := 2046;
        ELSIF x = 14474 THEN
            sigmoid_f := 2046;
        ELSIF x = 14475 THEN
            sigmoid_f := 2046;
        ELSIF x = 14476 THEN
            sigmoid_f := 2046;
        ELSIF x = 14477 THEN
            sigmoid_f := 2046;
        ELSIF x = 14478 THEN
            sigmoid_f := 2046;
        ELSIF x = 14479 THEN
            sigmoid_f := 2046;
        ELSIF x = 14480 THEN
            sigmoid_f := 2046;
        ELSIF x = 14481 THEN
            sigmoid_f := 2046;
        ELSIF x = 14482 THEN
            sigmoid_f := 2046;
        ELSIF x = 14483 THEN
            sigmoid_f := 2046;
        ELSIF x = 14484 THEN
            sigmoid_f := 2046;
        ELSIF x = 14485 THEN
            sigmoid_f := 2046;
        ELSIF x = 14486 THEN
            sigmoid_f := 2046;
        ELSIF x = 14487 THEN
            sigmoid_f := 2046;
        ELSIF x = 14488 THEN
            sigmoid_f := 2046;
        ELSIF x = 14489 THEN
            sigmoid_f := 2046;
        ELSIF x = 14490 THEN
            sigmoid_f := 2046;
        ELSIF x = 14491 THEN
            sigmoid_f := 2046;
        ELSIF x = 14492 THEN
            sigmoid_f := 2046;
        ELSIF x = 14493 THEN
            sigmoid_f := 2046;
        ELSIF x = 14494 THEN
            sigmoid_f := 2046;
        ELSIF x = 14495 THEN
            sigmoid_f := 2046;
        ELSIF x = 14496 THEN
            sigmoid_f := 2046;
        ELSIF x = 14497 THEN
            sigmoid_f := 2046;
        ELSIF x = 14498 THEN
            sigmoid_f := 2046;
        ELSIF x = 14499 THEN
            sigmoid_f := 2046;
        ELSIF x = 14500 THEN
            sigmoid_f := 2046;
        ELSIF x = 14501 THEN
            sigmoid_f := 2046;
        ELSIF x = 14502 THEN
            sigmoid_f := 2046;
        ELSIF x = 14503 THEN
            sigmoid_f := 2046;
        ELSIF x = 14504 THEN
            sigmoid_f := 2046;
        ELSIF x = 14505 THEN
            sigmoid_f := 2046;
        ELSIF x = 14506 THEN
            sigmoid_f := 2046;
        ELSIF x = 14507 THEN
            sigmoid_f := 2046;
        ELSIF x = 14508 THEN
            sigmoid_f := 2046;
        ELSIF x = 14509 THEN
            sigmoid_f := 2046;
        ELSIF x = 14510 THEN
            sigmoid_f := 2046;
        ELSIF x = 14511 THEN
            sigmoid_f := 2046;
        ELSIF x = 14512 THEN
            sigmoid_f := 2046;
        ELSIF x = 14513 THEN
            sigmoid_f := 2046;
        ELSIF x = 14514 THEN
            sigmoid_f := 2046;
        ELSIF x = 14515 THEN
            sigmoid_f := 2046;
        ELSIF x = 14516 THEN
            sigmoid_f := 2046;
        ELSIF x = 14517 THEN
            sigmoid_f := 2046;
        ELSIF x = 14518 THEN
            sigmoid_f := 2046;
        ELSIF x = 14519 THEN
            sigmoid_f := 2046;
        ELSIF x = 14520 THEN
            sigmoid_f := 2046;
        ELSIF x = 14521 THEN
            sigmoid_f := 2046;
        ELSIF x = 14522 THEN
            sigmoid_f := 2046;
        ELSIF x = 14523 THEN
            sigmoid_f := 2046;
        ELSIF x = 14524 THEN
            sigmoid_f := 2046;
        ELSIF x = 14525 THEN
            sigmoid_f := 2046;
        ELSIF x = 14526 THEN
            sigmoid_f := 2046;
        ELSIF x = 14527 THEN
            sigmoid_f := 2046;
        ELSIF x = 14528 THEN
            sigmoid_f := 2046;
        ELSIF x = 14529 THEN
            sigmoid_f := 2046;
        ELSIF x = 14530 THEN
            sigmoid_f := 2046;
        ELSIF x = 14531 THEN
            sigmoid_f := 2046;
        ELSIF x = 14532 THEN
            sigmoid_f := 2046;
        ELSIF x = 14533 THEN
            sigmoid_f := 2046;
        ELSIF x = 14534 THEN
            sigmoid_f := 2046;
        ELSIF x = 14535 THEN
            sigmoid_f := 2046;
        ELSIF x = 14536 THEN
            sigmoid_f := 2046;
        ELSIF x = 14537 THEN
            sigmoid_f := 2046;
        ELSIF x = 14538 THEN
            sigmoid_f := 2046;
        ELSIF x = 14539 THEN
            sigmoid_f := 2046;
        ELSIF x = 14540 THEN
            sigmoid_f := 2046;
        ELSIF x = 14541 THEN
            sigmoid_f := 2046;
        ELSIF x = 14542 THEN
            sigmoid_f := 2046;
        ELSIF x = 14543 THEN
            sigmoid_f := 2046;
        ELSIF x = 14544 THEN
            sigmoid_f := 2046;
        ELSIF x = 14545 THEN
            sigmoid_f := 2046;
        ELSIF x = 14546 THEN
            sigmoid_f := 2046;
        ELSIF x = 14547 THEN
            sigmoid_f := 2046;
        ELSIF x = 14548 THEN
            sigmoid_f := 2046;
        ELSIF x = 14549 THEN
            sigmoid_f := 2046;
        ELSIF x = 14550 THEN
            sigmoid_f := 2046;
        ELSIF x = 14551 THEN
            sigmoid_f := 2046;
        ELSIF x = 14552 THEN
            sigmoid_f := 2046;
        ELSIF x = 14553 THEN
            sigmoid_f := 2046;
        ELSIF x = 14554 THEN
            sigmoid_f := 2046;
        ELSIF x = 14555 THEN
            sigmoid_f := 2046;
        ELSIF x = 14556 THEN
            sigmoid_f := 2046;
        ELSIF x = 14557 THEN
            sigmoid_f := 2046;
        ELSIF x = 14558 THEN
            sigmoid_f := 2046;
        ELSIF x = 14559 THEN
            sigmoid_f := 2046;
        ELSIF x = 14560 THEN
            sigmoid_f := 2046;
        ELSIF x = 14561 THEN
            sigmoid_f := 2046;
        ELSIF x = 14562 THEN
            sigmoid_f := 2046;
        ELSIF x = 14563 THEN
            sigmoid_f := 2046;
        ELSIF x = 14564 THEN
            sigmoid_f := 2046;
        ELSIF x = 14565 THEN
            sigmoid_f := 2046;
        ELSIF x = 14566 THEN
            sigmoid_f := 2046;
        ELSIF x = 14567 THEN
            sigmoid_f := 2046;
        ELSIF x = 14568 THEN
            sigmoid_f := 2046;
        ELSIF x = 14569 THEN
            sigmoid_f := 2046;
        ELSIF x = 14570 THEN
            sigmoid_f := 2046;
        ELSIF x = 14571 THEN
            sigmoid_f := 2046;
        ELSIF x = 14572 THEN
            sigmoid_f := 2046;
        ELSIF x = 14573 THEN
            sigmoid_f := 2046;
        ELSIF x = 14574 THEN
            sigmoid_f := 2046;
        ELSIF x = 14575 THEN
            sigmoid_f := 2046;
        ELSIF x = 14576 THEN
            sigmoid_f := 2046;
        ELSIF x = 14577 THEN
            sigmoid_f := 2046;
        ELSIF x = 14578 THEN
            sigmoid_f := 2046;
        ELSIF x = 14579 THEN
            sigmoid_f := 2046;
        ELSIF x = 14580 THEN
            sigmoid_f := 2046;
        ELSIF x = 14581 THEN
            sigmoid_f := 2046;
        ELSIF x = 14582 THEN
            sigmoid_f := 2046;
        ELSIF x = 14583 THEN
            sigmoid_f := 2046;
        ELSIF x = 14584 THEN
            sigmoid_f := 2046;
        ELSIF x = 14585 THEN
            sigmoid_f := 2046;
        ELSIF x = 14586 THEN
            sigmoid_f := 2046;
        ELSIF x = 14587 THEN
            sigmoid_f := 2046;
        ELSIF x = 14588 THEN
            sigmoid_f := 2046;
        ELSIF x = 14589 THEN
            sigmoid_f := 2046;
        ELSIF x = 14590 THEN
            sigmoid_f := 2046;
        ELSIF x = 14591 THEN
            sigmoid_f := 2046;
        ELSIF x = 14592 THEN
            sigmoid_f := 2046;
        ELSIF x = 14593 THEN
            sigmoid_f := 2046;
        ELSIF x = 14594 THEN
            sigmoid_f := 2046;
        ELSIF x = 14595 THEN
            sigmoid_f := 2046;
        ELSIF x = 14596 THEN
            sigmoid_f := 2046;
        ELSIF x = 14597 THEN
            sigmoid_f := 2046;
        ELSIF x = 14598 THEN
            sigmoid_f := 2046;
        ELSIF x = 14599 THEN
            sigmoid_f := 2046;
        ELSIF x = 14600 THEN
            sigmoid_f := 2046;
        ELSIF x = 14601 THEN
            sigmoid_f := 2046;
        ELSIF x = 14602 THEN
            sigmoid_f := 2046;
        ELSIF x = 14603 THEN
            sigmoid_f := 2046;
        ELSIF x = 14604 THEN
            sigmoid_f := 2046;
        ELSIF x = 14605 THEN
            sigmoid_f := 2046;
        ELSIF x = 14606 THEN
            sigmoid_f := 2046;
        ELSIF x = 14607 THEN
            sigmoid_f := 2046;
        ELSIF x = 14608 THEN
            sigmoid_f := 2046;
        ELSIF x = 14609 THEN
            sigmoid_f := 2046;
        ELSIF x = 14610 THEN
            sigmoid_f := 2046;
        ELSIF x = 14611 THEN
            sigmoid_f := 2046;
        ELSIF x = 14612 THEN
            sigmoid_f := 2046;
        ELSIF x = 14613 THEN
            sigmoid_f := 2046;
        ELSIF x = 14614 THEN
            sigmoid_f := 2046;
        ELSIF x = 14615 THEN
            sigmoid_f := 2046;
        ELSIF x = 14616 THEN
            sigmoid_f := 2046;
        ELSIF x = 14617 THEN
            sigmoid_f := 2046;
        ELSIF x = 14618 THEN
            sigmoid_f := 2046;
        ELSIF x = 14619 THEN
            sigmoid_f := 2046;
        ELSIF x = 14620 THEN
            sigmoid_f := 2046;
        ELSIF x = 14621 THEN
            sigmoid_f := 2046;
        ELSIF x = 14622 THEN
            sigmoid_f := 2046;
        ELSIF x = 14623 THEN
            sigmoid_f := 2046;
        ELSIF x = 14624 THEN
            sigmoid_f := 2046;
        ELSIF x = 14625 THEN
            sigmoid_f := 2046;
        ELSIF x = 14626 THEN
            sigmoid_f := 2046;
        ELSIF x = 14627 THEN
            sigmoid_f := 2046;
        ELSIF x = 14628 THEN
            sigmoid_f := 2046;
        ELSIF x = 14629 THEN
            sigmoid_f := 2046;
        ELSIF x = 14630 THEN
            sigmoid_f := 2046;
        ELSIF x = 14631 THEN
            sigmoid_f := 2046;
        ELSIF x = 14632 THEN
            sigmoid_f := 2046;
        ELSIF x = 14633 THEN
            sigmoid_f := 2046;
        ELSIF x = 14634 THEN
            sigmoid_f := 2046;
        ELSIF x = 14635 THEN
            sigmoid_f := 2046;
        ELSIF x = 14636 THEN
            sigmoid_f := 2046;
        ELSIF x = 14637 THEN
            sigmoid_f := 2046;
        ELSIF x = 14638 THEN
            sigmoid_f := 2046;
        ELSIF x = 14639 THEN
            sigmoid_f := 2046;
        ELSIF x = 14640 THEN
            sigmoid_f := 2046;
        ELSIF x = 14641 THEN
            sigmoid_f := 2046;
        ELSIF x = 14642 THEN
            sigmoid_f := 2046;
        ELSIF x = 14643 THEN
            sigmoid_f := 2046;
        ELSIF x = 14644 THEN
            sigmoid_f := 2046;
        ELSIF x = 14645 THEN
            sigmoid_f := 2046;
        ELSIF x = 14646 THEN
            sigmoid_f := 2046;
        ELSIF x = 14647 THEN
            sigmoid_f := 2046;
        ELSIF x = 14648 THEN
            sigmoid_f := 2046;
        ELSIF x = 14649 THEN
            sigmoid_f := 2046;
        ELSIF x = 14650 THEN
            sigmoid_f := 2046;
        ELSIF x = 14651 THEN
            sigmoid_f := 2046;
        ELSIF x = 14652 THEN
            sigmoid_f := 2046;
        ELSIF x = 14653 THEN
            sigmoid_f := 2046;
        ELSIF x = 14654 THEN
            sigmoid_f := 2046;
        ELSIF x = 14655 THEN
            sigmoid_f := 2046;
        ELSIF x = 14656 THEN
            sigmoid_f := 2046;
        ELSIF x = 14657 THEN
            sigmoid_f := 2046;
        ELSIF x = 14658 THEN
            sigmoid_f := 2046;
        ELSIF x = 14659 THEN
            sigmoid_f := 2046;
        ELSIF x = 14660 THEN
            sigmoid_f := 2046;
        ELSIF x = 14661 THEN
            sigmoid_f := 2046;
        ELSIF x = 14662 THEN
            sigmoid_f := 2046;
        ELSIF x = 14663 THEN
            sigmoid_f := 2046;
        ELSIF x = 14664 THEN
            sigmoid_f := 2046;
        ELSIF x = 14665 THEN
            sigmoid_f := 2046;
        ELSIF x = 14666 THEN
            sigmoid_f := 2046;
        ELSIF x = 14667 THEN
            sigmoid_f := 2046;
        ELSIF x = 14668 THEN
            sigmoid_f := 2046;
        ELSIF x = 14669 THEN
            sigmoid_f := 2046;
        ELSIF x = 14670 THEN
            sigmoid_f := 2046;
        ELSIF x = 14671 THEN
            sigmoid_f := 2046;
        ELSIF x = 14672 THEN
            sigmoid_f := 2046;
        ELSIF x = 14673 THEN
            sigmoid_f := 2046;
        ELSIF x = 14674 THEN
            sigmoid_f := 2046;
        ELSIF x = 14675 THEN
            sigmoid_f := 2046;
        ELSIF x = 14676 THEN
            sigmoid_f := 2046;
        ELSIF x = 14677 THEN
            sigmoid_f := 2046;
        ELSIF x = 14678 THEN
            sigmoid_f := 2046;
        ELSIF x = 14679 THEN
            sigmoid_f := 2046;
        ELSIF x = 14680 THEN
            sigmoid_f := 2046;
        ELSIF x = 14681 THEN
            sigmoid_f := 2046;
        ELSIF x = 14682 THEN
            sigmoid_f := 2046;
        ELSIF x = 14683 THEN
            sigmoid_f := 2046;
        ELSIF x = 14684 THEN
            sigmoid_f := 2046;
        ELSIF x = 14685 THEN
            sigmoid_f := 2046;
        ELSIF x = 14686 THEN
            sigmoid_f := 2046;
        ELSIF x = 14687 THEN
            sigmoid_f := 2046;
        ELSIF x = 14688 THEN
            sigmoid_f := 2046;
        ELSIF x = 14689 THEN
            sigmoid_f := 2046;
        ELSIF x = 14690 THEN
            sigmoid_f := 2046;
        ELSIF x = 14691 THEN
            sigmoid_f := 2046;
        ELSIF x = 14692 THEN
            sigmoid_f := 2046;
        ELSIF x = 14693 THEN
            sigmoid_f := 2046;
        ELSIF x = 14694 THEN
            sigmoid_f := 2046;
        ELSIF x = 14695 THEN
            sigmoid_f := 2046;
        ELSIF x = 14696 THEN
            sigmoid_f := 2046;
        ELSIF x = 14697 THEN
            sigmoid_f := 2046;
        ELSIF x = 14698 THEN
            sigmoid_f := 2046;
        ELSIF x = 14699 THEN
            sigmoid_f := 2046;
        ELSIF x = 14700 THEN
            sigmoid_f := 2046;
        ELSIF x = 14701 THEN
            sigmoid_f := 2046;
        ELSIF x = 14702 THEN
            sigmoid_f := 2046;
        ELSIF x = 14703 THEN
            sigmoid_f := 2046;
        ELSIF x = 14704 THEN
            sigmoid_f := 2046;
        ELSIF x = 14705 THEN
            sigmoid_f := 2046;
        ELSIF x = 14706 THEN
            sigmoid_f := 2046;
        ELSIF x = 14707 THEN
            sigmoid_f := 2046;
        ELSIF x = 14708 THEN
            sigmoid_f := 2046;
        ELSIF x = 14709 THEN
            sigmoid_f := 2046;
        ELSIF x = 14710 THEN
            sigmoid_f := 2046;
        ELSIF x = 14711 THEN
            sigmoid_f := 2046;
        ELSIF x = 14712 THEN
            sigmoid_f := 2046;
        ELSIF x = 14713 THEN
            sigmoid_f := 2046;
        ELSIF x = 14714 THEN
            sigmoid_f := 2046;
        ELSIF x = 14715 THEN
            sigmoid_f := 2046;
        ELSIF x = 14716 THEN
            sigmoid_f := 2046;
        ELSIF x = 14717 THEN
            sigmoid_f := 2046;
        ELSIF x = 14718 THEN
            sigmoid_f := 2046;
        ELSIF x = 14719 THEN
            sigmoid_f := 2046;
        ELSIF x = 14720 THEN
            sigmoid_f := 2046;
        ELSIF x = 14721 THEN
            sigmoid_f := 2046;
        ELSIF x = 14722 THEN
            sigmoid_f := 2046;
        ELSIF x = 14723 THEN
            sigmoid_f := 2046;
        ELSIF x = 14724 THEN
            sigmoid_f := 2046;
        ELSIF x = 14725 THEN
            sigmoid_f := 2046;
        ELSIF x = 14726 THEN
            sigmoid_f := 2046;
        ELSIF x = 14727 THEN
            sigmoid_f := 2046;
        ELSIF x = 14728 THEN
            sigmoid_f := 2046;
        ELSIF x = 14729 THEN
            sigmoid_f := 2046;
        ELSIF x = 14730 THEN
            sigmoid_f := 2046;
        ELSIF x = 14731 THEN
            sigmoid_f := 2046;
        ELSIF x = 14732 THEN
            sigmoid_f := 2046;
        ELSIF x = 14733 THEN
            sigmoid_f := 2046;
        ELSIF x = 14734 THEN
            sigmoid_f := 2046;
        ELSIF x = 14735 THEN
            sigmoid_f := 2046;
        ELSIF x = 14736 THEN
            sigmoid_f := 2046;
        ELSIF x = 14737 THEN
            sigmoid_f := 2046;
        ELSIF x = 14738 THEN
            sigmoid_f := 2046;
        ELSIF x = 14739 THEN
            sigmoid_f := 2046;
        ELSIF x = 14740 THEN
            sigmoid_f := 2046;
        ELSIF x = 14741 THEN
            sigmoid_f := 2046;
        ELSIF x = 14742 THEN
            sigmoid_f := 2046;
        ELSIF x = 14743 THEN
            sigmoid_f := 2046;
        ELSIF x = 14744 THEN
            sigmoid_f := 2046;
        ELSIF x = 14745 THEN
            sigmoid_f := 2046;
        ELSIF x = 14746 THEN
            sigmoid_f := 2046;
        ELSIF x = 14747 THEN
            sigmoid_f := 2046;
        ELSIF x = 14748 THEN
            sigmoid_f := 2046;
        ELSIF x = 14749 THEN
            sigmoid_f := 2046;
        ELSIF x = 14750 THEN
            sigmoid_f := 2046;
        ELSIF x = 14751 THEN
            sigmoid_f := 2046;
        ELSIF x = 14752 THEN
            sigmoid_f := 2046;
        ELSIF x = 14753 THEN
            sigmoid_f := 2046;
        ELSIF x = 14754 THEN
            sigmoid_f := 2046;
        ELSIF x = 14755 THEN
            sigmoid_f := 2046;
        ELSIF x = 14756 THEN
            sigmoid_f := 2046;
        ELSIF x = 14757 THEN
            sigmoid_f := 2046;
        ELSIF x = 14758 THEN
            sigmoid_f := 2046;
        ELSIF x = 14759 THEN
            sigmoid_f := 2046;
        ELSIF x = 14760 THEN
            sigmoid_f := 2046;
        ELSIF x = 14761 THEN
            sigmoid_f := 2046;
        ELSIF x = 14762 THEN
            sigmoid_f := 2046;
        ELSIF x = 14763 THEN
            sigmoid_f := 2046;
        ELSIF x = 14764 THEN
            sigmoid_f := 2046;
        ELSIF x = 14765 THEN
            sigmoid_f := 2046;
        ELSIF x = 14766 THEN
            sigmoid_f := 2046;
        ELSIF x = 14767 THEN
            sigmoid_f := 2046;
        ELSIF x = 14768 THEN
            sigmoid_f := 2046;
        ELSIF x = 14769 THEN
            sigmoid_f := 2046;
        ELSIF x = 14770 THEN
            sigmoid_f := 2046;
        ELSIF x = 14771 THEN
            sigmoid_f := 2046;
        ELSIF x = 14772 THEN
            sigmoid_f := 2046;
        ELSIF x = 14773 THEN
            sigmoid_f := 2046;
        ELSIF x = 14774 THEN
            sigmoid_f := 2046;
        ELSIF x = 14775 THEN
            sigmoid_f := 2046;
        ELSIF x = 14776 THEN
            sigmoid_f := 2046;
        ELSIF x = 14777 THEN
            sigmoid_f := 2046;
        ELSIF x = 14778 THEN
            sigmoid_f := 2046;
        ELSIF x = 14779 THEN
            sigmoid_f := 2046;
        ELSIF x = 14780 THEN
            sigmoid_f := 2046;
        ELSIF x = 14781 THEN
            sigmoid_f := 2046;
        ELSIF x = 14782 THEN
            sigmoid_f := 2046;
        ELSIF x = 14783 THEN
            sigmoid_f := 2046;
        ELSIF x = 14784 THEN
            sigmoid_f := 2046;
        ELSIF x = 14785 THEN
            sigmoid_f := 2046;
        ELSIF x = 14786 THEN
            sigmoid_f := 2046;
        ELSIF x = 14787 THEN
            sigmoid_f := 2046;
        ELSIF x = 14788 THEN
            sigmoid_f := 2046;
        ELSIF x = 14789 THEN
            sigmoid_f := 2046;
        ELSIF x = 14790 THEN
            sigmoid_f := 2046;
        ELSIF x = 14791 THEN
            sigmoid_f := 2046;
        ELSIF x = 14792 THEN
            sigmoid_f := 2046;
        ELSIF x = 14793 THEN
            sigmoid_f := 2046;
        ELSIF x = 14794 THEN
            sigmoid_f := 2046;
        ELSIF x = 14795 THEN
            sigmoid_f := 2046;
        ELSIF x = 14796 THEN
            sigmoid_f := 2046;
        ELSIF x = 14797 THEN
            sigmoid_f := 2046;
        ELSIF x = 14798 THEN
            sigmoid_f := 2046;
        ELSIF x = 14799 THEN
            sigmoid_f := 2046;
        ELSIF x = 14800 THEN
            sigmoid_f := 2046;
        ELSIF x = 14801 THEN
            sigmoid_f := 2046;
        ELSIF x = 14802 THEN
            sigmoid_f := 2046;
        ELSIF x = 14803 THEN
            sigmoid_f := 2046;
        ELSIF x = 14804 THEN
            sigmoid_f := 2046;
        ELSIF x = 14805 THEN
            sigmoid_f := 2046;
        ELSIF x = 14806 THEN
            sigmoid_f := 2046;
        ELSIF x = 14807 THEN
            sigmoid_f := 2046;
        ELSIF x = 14808 THEN
            sigmoid_f := 2046;
        ELSIF x = 14809 THEN
            sigmoid_f := 2046;
        ELSIF x = 14810 THEN
            sigmoid_f := 2046;
        ELSIF x = 14811 THEN
            sigmoid_f := 2046;
        ELSIF x = 14812 THEN
            sigmoid_f := 2046;
        ELSIF x = 14813 THEN
            sigmoid_f := 2046;
        ELSIF x = 14814 THEN
            sigmoid_f := 2046;
        ELSIF x = 14815 THEN
            sigmoid_f := 2046;
        ELSIF x = 14816 THEN
            sigmoid_f := 2046;
        ELSIF x = 14817 THEN
            sigmoid_f := 2046;
        ELSIF x = 14818 THEN
            sigmoid_f := 2046;
        ELSIF x = 14819 THEN
            sigmoid_f := 2046;
        ELSIF x = 14820 THEN
            sigmoid_f := 2046;
        ELSIF x = 14821 THEN
            sigmoid_f := 2046;
        ELSIF x = 14822 THEN
            sigmoid_f := 2046;
        ELSIF x = 14823 THEN
            sigmoid_f := 2046;
        ELSIF x = 14824 THEN
            sigmoid_f := 2046;
        ELSIF x = 14825 THEN
            sigmoid_f := 2046;
        ELSIF x = 14826 THEN
            sigmoid_f := 2046;
        ELSIF x = 14827 THEN
            sigmoid_f := 2046;
        ELSIF x = 14828 THEN
            sigmoid_f := 2046;
        ELSIF x = 14829 THEN
            sigmoid_f := 2046;
        ELSIF x = 14830 THEN
            sigmoid_f := 2046;
        ELSIF x = 14831 THEN
            sigmoid_f := 2046;
        ELSIF x = 14832 THEN
            sigmoid_f := 2046;
        ELSIF x = 14833 THEN
            sigmoid_f := 2046;
        ELSIF x = 14834 THEN
            sigmoid_f := 2046;
        ELSIF x = 14835 THEN
            sigmoid_f := 2046;
        ELSIF x = 14836 THEN
            sigmoid_f := 2046;
        ELSIF x = 14837 THEN
            sigmoid_f := 2046;
        ELSIF x = 14838 THEN
            sigmoid_f := 2046;
        ELSIF x = 14839 THEN
            sigmoid_f := 2046;
        ELSIF x = 14840 THEN
            sigmoid_f := 2046;
        ELSIF x = 14841 THEN
            sigmoid_f := 2046;
        ELSIF x = 14842 THEN
            sigmoid_f := 2046;
        ELSIF x = 14843 THEN
            sigmoid_f := 2046;
        ELSIF x = 14844 THEN
            sigmoid_f := 2046;
        ELSIF x = 14845 THEN
            sigmoid_f := 2046;
        ELSIF x = 14846 THEN
            sigmoid_f := 2046;
        ELSIF x = 14847 THEN
            sigmoid_f := 2046;
        ELSIF x = 14848 THEN
            sigmoid_f := 2047;
        ELSIF x = 14849 THEN
            sigmoid_f := 2047;
        ELSIF x = 14850 THEN
            sigmoid_f := 2047;
        ELSIF x = 14851 THEN
            sigmoid_f := 2047;
        ELSIF x = 14852 THEN
            sigmoid_f := 2047;
        ELSIF x = 14853 THEN
            sigmoid_f := 2047;
        ELSIF x = 14854 THEN
            sigmoid_f := 2047;
        ELSIF x = 14855 THEN
            sigmoid_f := 2047;
        ELSIF x = 14856 THEN
            sigmoid_f := 2047;
        ELSIF x = 14857 THEN
            sigmoid_f := 2047;
        ELSIF x = 14858 THEN
            sigmoid_f := 2047;
        ELSIF x = 14859 THEN
            sigmoid_f := 2047;
        ELSIF x = 14860 THEN
            sigmoid_f := 2047;
        ELSIF x = 14861 THEN
            sigmoid_f := 2047;
        ELSIF x = 14862 THEN
            sigmoid_f := 2047;
        ELSIF x = 14863 THEN
            sigmoid_f := 2047;
        ELSIF x = 14864 THEN
            sigmoid_f := 2047;
        ELSIF x = 14865 THEN
            sigmoid_f := 2047;
        ELSIF x = 14866 THEN
            sigmoid_f := 2047;
        ELSIF x = 14867 THEN
            sigmoid_f := 2047;
        ELSIF x = 14868 THEN
            sigmoid_f := 2047;
        ELSIF x = 14869 THEN
            sigmoid_f := 2047;
        ELSIF x = 14870 THEN
            sigmoid_f := 2047;
        ELSIF x = 14871 THEN
            sigmoid_f := 2047;
        ELSIF x = 14872 THEN
            sigmoid_f := 2047;
        ELSIF x = 14873 THEN
            sigmoid_f := 2047;
        ELSIF x = 14874 THEN
            sigmoid_f := 2047;
        ELSIF x = 14875 THEN
            sigmoid_f := 2047;
        ELSIF x = 14876 THEN
            sigmoid_f := 2047;
        ELSIF x = 14877 THEN
            sigmoid_f := 2047;
        ELSIF x = 14878 THEN
            sigmoid_f := 2047;
        ELSIF x = 14879 THEN
            sigmoid_f := 2047;
        ELSIF x = 14880 THEN
            sigmoid_f := 2047;
        ELSIF x = 14881 THEN
            sigmoid_f := 2047;
        ELSIF x = 14882 THEN
            sigmoid_f := 2047;
        ELSIF x = 14883 THEN
            sigmoid_f := 2047;
        ELSIF x = 14884 THEN
            sigmoid_f := 2047;
        ELSIF x = 14885 THEN
            sigmoid_f := 2047;
        ELSIF x = 14886 THEN
            sigmoid_f := 2047;
        ELSIF x = 14887 THEN
            sigmoid_f := 2047;
        ELSIF x = 14888 THEN
            sigmoid_f := 2047;
        ELSIF x = 14889 THEN
            sigmoid_f := 2047;
        ELSIF x = 14890 THEN
            sigmoid_f := 2047;
        ELSIF x = 14891 THEN
            sigmoid_f := 2047;
        ELSIF x = 14892 THEN
            sigmoid_f := 2047;
        ELSIF x = 14893 THEN
            sigmoid_f := 2047;
        ELSIF x = 14894 THEN
            sigmoid_f := 2047;
        ELSIF x = 14895 THEN
            sigmoid_f := 2047;
        ELSIF x = 14896 THEN
            sigmoid_f := 2047;
        ELSIF x = 14897 THEN
            sigmoid_f := 2047;
        ELSIF x = 14898 THEN
            sigmoid_f := 2047;
        ELSIF x = 14899 THEN
            sigmoid_f := 2047;
        ELSIF x = 14900 THEN
            sigmoid_f := 2047;
        ELSIF x = 14901 THEN
            sigmoid_f := 2047;
        ELSIF x = 14902 THEN
            sigmoid_f := 2047;
        ELSIF x = 14903 THEN
            sigmoid_f := 2047;
        ELSIF x = 14904 THEN
            sigmoid_f := 2047;
        ELSIF x = 14905 THEN
            sigmoid_f := 2047;
        ELSIF x = 14906 THEN
            sigmoid_f := 2047;
        ELSIF x = 14907 THEN
            sigmoid_f := 2047;
        ELSIF x = 14908 THEN
            sigmoid_f := 2047;
        ELSIF x = 14909 THEN
            sigmoid_f := 2047;
        ELSIF x = 14910 THEN
            sigmoid_f := 2047;
        ELSIF x = 14911 THEN
            sigmoid_f := 2047;
        ELSIF x = 14912 THEN
            sigmoid_f := 2047;
        ELSIF x = 14913 THEN
            sigmoid_f := 2047;
        ELSIF x = 14914 THEN
            sigmoid_f := 2047;
        ELSIF x = 14915 THEN
            sigmoid_f := 2047;
        ELSIF x = 14916 THEN
            sigmoid_f := 2047;
        ELSIF x = 14917 THEN
            sigmoid_f := 2047;
        ELSIF x = 14918 THEN
            sigmoid_f := 2047;
        ELSIF x = 14919 THEN
            sigmoid_f := 2047;
        ELSIF x = 14920 THEN
            sigmoid_f := 2047;
        ELSIF x = 14921 THEN
            sigmoid_f := 2047;
        ELSIF x = 14922 THEN
            sigmoid_f := 2047;
        ELSIF x = 14923 THEN
            sigmoid_f := 2047;
        ELSIF x = 14924 THEN
            sigmoid_f := 2047;
        ELSIF x = 14925 THEN
            sigmoid_f := 2047;
        ELSIF x = 14926 THEN
            sigmoid_f := 2047;
        ELSIF x = 14927 THEN
            sigmoid_f := 2047;
        ELSIF x = 14928 THEN
            sigmoid_f := 2047;
        ELSIF x = 14929 THEN
            sigmoid_f := 2047;
        ELSIF x = 14930 THEN
            sigmoid_f := 2047;
        ELSIF x = 14931 THEN
            sigmoid_f := 2047;
        ELSIF x = 14932 THEN
            sigmoid_f := 2047;
        ELSIF x = 14933 THEN
            sigmoid_f := 2047;
        ELSIF x = 14934 THEN
            sigmoid_f := 2047;
        ELSIF x = 14935 THEN
            sigmoid_f := 2047;
        ELSIF x = 14936 THEN
            sigmoid_f := 2047;
        ELSIF x = 14937 THEN
            sigmoid_f := 2047;
        ELSIF x = 14938 THEN
            sigmoid_f := 2047;
        ELSIF x = 14939 THEN
            sigmoid_f := 2047;
        ELSIF x = 14940 THEN
            sigmoid_f := 2047;
        ELSIF x = 14941 THEN
            sigmoid_f := 2047;
        ELSIF x = 14942 THEN
            sigmoid_f := 2047;
        ELSIF x = 14943 THEN
            sigmoid_f := 2047;
        ELSIF x = 14944 THEN
            sigmoid_f := 2047;
        ELSIF x = 14945 THEN
            sigmoid_f := 2047;
        ELSIF x = 14946 THEN
            sigmoid_f := 2047;
        ELSIF x = 14947 THEN
            sigmoid_f := 2047;
        ELSIF x = 14948 THEN
            sigmoid_f := 2047;
        ELSIF x = 14949 THEN
            sigmoid_f := 2047;
        ELSIF x = 14950 THEN
            sigmoid_f := 2047;
        ELSIF x = 14951 THEN
            sigmoid_f := 2047;
        ELSIF x = 14952 THEN
            sigmoid_f := 2047;
        ELSIF x = 14953 THEN
            sigmoid_f := 2047;
        ELSIF x = 14954 THEN
            sigmoid_f := 2047;
        ELSIF x = 14955 THEN
            sigmoid_f := 2047;
        ELSIF x = 14956 THEN
            sigmoid_f := 2047;
        ELSIF x = 14957 THEN
            sigmoid_f := 2047;
        ELSIF x = 14958 THEN
            sigmoid_f := 2047;
        ELSIF x = 14959 THEN
            sigmoid_f := 2047;
        ELSIF x = 14960 THEN
            sigmoid_f := 2047;
        ELSIF x = 14961 THEN
            sigmoid_f := 2047;
        ELSIF x = 14962 THEN
            sigmoid_f := 2047;
        ELSIF x = 14963 THEN
            sigmoid_f := 2047;
        ELSIF x = 14964 THEN
            sigmoid_f := 2047;
        ELSIF x = 14965 THEN
            sigmoid_f := 2047;
        ELSIF x = 14966 THEN
            sigmoid_f := 2047;
        ELSIF x = 14967 THEN
            sigmoid_f := 2047;
        ELSIF x = 14968 THEN
            sigmoid_f := 2047;
        ELSIF x = 14969 THEN
            sigmoid_f := 2047;
        ELSIF x = 14970 THEN
            sigmoid_f := 2047;
        ELSIF x = 14971 THEN
            sigmoid_f := 2047;
        ELSIF x = 14972 THEN
            sigmoid_f := 2047;
        ELSIF x = 14973 THEN
            sigmoid_f := 2047;
        ELSIF x = 14974 THEN
            sigmoid_f := 2047;
        ELSIF x = 14975 THEN
            sigmoid_f := 2047;
        ELSIF x = 14976 THEN
            sigmoid_f := 2047;
        ELSIF x = 14977 THEN
            sigmoid_f := 2047;
        ELSIF x = 14978 THEN
            sigmoid_f := 2047;
        ELSIF x = 14979 THEN
            sigmoid_f := 2047;
        ELSIF x = 14980 THEN
            sigmoid_f := 2047;
        ELSIF x = 14981 THEN
            sigmoid_f := 2047;
        ELSIF x = 14982 THEN
            sigmoid_f := 2047;
        ELSIF x = 14983 THEN
            sigmoid_f := 2047;
        ELSIF x = 14984 THEN
            sigmoid_f := 2047;
        ELSIF x = 14985 THEN
            sigmoid_f := 2047;
        ELSIF x = 14986 THEN
            sigmoid_f := 2047;
        ELSIF x = 14987 THEN
            sigmoid_f := 2047;
        ELSIF x = 14988 THEN
            sigmoid_f := 2047;
        ELSIF x = 14989 THEN
            sigmoid_f := 2047;
        ELSIF x = 14990 THEN
            sigmoid_f := 2047;
        ELSIF x = 14991 THEN
            sigmoid_f := 2047;
        ELSIF x = 14992 THEN
            sigmoid_f := 2047;
        ELSIF x = 14993 THEN
            sigmoid_f := 2047;
        ELSIF x = 14994 THEN
            sigmoid_f := 2047;
        ELSIF x = 14995 THEN
            sigmoid_f := 2047;
        ELSIF x = 14996 THEN
            sigmoid_f := 2047;
        ELSIF x = 14997 THEN
            sigmoid_f := 2047;
        ELSIF x = 14998 THEN
            sigmoid_f := 2047;
        ELSIF x = 14999 THEN
            sigmoid_f := 2047;
        ELSIF x = 15000 THEN
            sigmoid_f := 2047;
        ELSIF x = 15001 THEN
            sigmoid_f := 2047;
        ELSIF x = 15002 THEN
            sigmoid_f := 2047;
        ELSIF x = 15003 THEN
            sigmoid_f := 2047;
        ELSIF x = 15004 THEN
            sigmoid_f := 2047;
        ELSIF x = 15005 THEN
            sigmoid_f := 2047;
        ELSIF x = 15006 THEN
            sigmoid_f := 2047;
        ELSIF x = 15007 THEN
            sigmoid_f := 2047;
        ELSIF x = 15008 THEN
            sigmoid_f := 2047;
        ELSIF x = 15009 THEN
            sigmoid_f := 2047;
        ELSIF x = 15010 THEN
            sigmoid_f := 2047;
        ELSIF x = 15011 THEN
            sigmoid_f := 2047;
        ELSIF x = 15012 THEN
            sigmoid_f := 2047;
        ELSIF x = 15013 THEN
            sigmoid_f := 2047;
        ELSIF x = 15014 THEN
            sigmoid_f := 2047;
        ELSIF x = 15015 THEN
            sigmoid_f := 2047;
        ELSIF x = 15016 THEN
            sigmoid_f := 2047;
        ELSIF x = 15017 THEN
            sigmoid_f := 2047;
        ELSIF x = 15018 THEN
            sigmoid_f := 2047;
        ELSIF x = 15019 THEN
            sigmoid_f := 2047;
        ELSIF x = 15020 THEN
            sigmoid_f := 2047;
        ELSIF x = 15021 THEN
            sigmoid_f := 2047;
        ELSIF x = 15022 THEN
            sigmoid_f := 2047;
        ELSIF x = 15023 THEN
            sigmoid_f := 2047;
        ELSIF x = 15024 THEN
            sigmoid_f := 2047;
        ELSIF x = 15025 THEN
            sigmoid_f := 2047;
        ELSIF x = 15026 THEN
            sigmoid_f := 2047;
        ELSIF x = 15027 THEN
            sigmoid_f := 2047;
        ELSIF x = 15028 THEN
            sigmoid_f := 2047;
        ELSIF x = 15029 THEN
            sigmoid_f := 2047;
        ELSIF x = 15030 THEN
            sigmoid_f := 2047;
        ELSIF x = 15031 THEN
            sigmoid_f := 2047;
        ELSIF x = 15032 THEN
            sigmoid_f := 2047;
        ELSIF x = 15033 THEN
            sigmoid_f := 2047;
        ELSIF x = 15034 THEN
            sigmoid_f := 2047;
        ELSIF x = 15035 THEN
            sigmoid_f := 2047;
        ELSIF x = 15036 THEN
            sigmoid_f := 2047;
        ELSIF x = 15037 THEN
            sigmoid_f := 2047;
        ELSIF x = 15038 THEN
            sigmoid_f := 2047;
        ELSIF x = 15039 THEN
            sigmoid_f := 2047;
        ELSIF x = 15040 THEN
            sigmoid_f := 2047;
        ELSIF x = 15041 THEN
            sigmoid_f := 2047;
        ELSIF x = 15042 THEN
            sigmoid_f := 2047;
        ELSIF x = 15043 THEN
            sigmoid_f := 2047;
        ELSIF x = 15044 THEN
            sigmoid_f := 2047;
        ELSIF x = 15045 THEN
            sigmoid_f := 2047;
        ELSIF x = 15046 THEN
            sigmoid_f := 2047;
        ELSIF x = 15047 THEN
            sigmoid_f := 2047;
        ELSIF x = 15048 THEN
            sigmoid_f := 2047;
        ELSIF x = 15049 THEN
            sigmoid_f := 2047;
        ELSIF x = 15050 THEN
            sigmoid_f := 2047;
        ELSIF x = 15051 THEN
            sigmoid_f := 2047;
        ELSIF x = 15052 THEN
            sigmoid_f := 2047;
        ELSIF x = 15053 THEN
            sigmoid_f := 2047;
        ELSIF x = 15054 THEN
            sigmoid_f := 2047;
        ELSIF x = 15055 THEN
            sigmoid_f := 2047;
        ELSIF x = 15056 THEN
            sigmoid_f := 2047;
        ELSIF x = 15057 THEN
            sigmoid_f := 2047;
        ELSIF x = 15058 THEN
            sigmoid_f := 2047;
        ELSIF x = 15059 THEN
            sigmoid_f := 2047;
        ELSIF x = 15060 THEN
            sigmoid_f := 2047;
        ELSIF x = 15061 THEN
            sigmoid_f := 2047;
        ELSIF x = 15062 THEN
            sigmoid_f := 2047;
        ELSIF x = 15063 THEN
            sigmoid_f := 2047;
        ELSIF x = 15064 THEN
            sigmoid_f := 2047;
        ELSIF x = 15065 THEN
            sigmoid_f := 2047;
        ELSIF x = 15066 THEN
            sigmoid_f := 2047;
        ELSIF x = 15067 THEN
            sigmoid_f := 2047;
        ELSIF x = 15068 THEN
            sigmoid_f := 2047;
        ELSIF x = 15069 THEN
            sigmoid_f := 2047;
        ELSIF x = 15070 THEN
            sigmoid_f := 2047;
        ELSIF x = 15071 THEN
            sigmoid_f := 2047;
        ELSIF x = 15072 THEN
            sigmoid_f := 2047;
        ELSIF x = 15073 THEN
            sigmoid_f := 2047;
        ELSIF x = 15074 THEN
            sigmoid_f := 2047;
        ELSIF x = 15075 THEN
            sigmoid_f := 2047;
        ELSIF x = 15076 THEN
            sigmoid_f := 2047;
        ELSIF x = 15077 THEN
            sigmoid_f := 2047;
        ELSIF x = 15078 THEN
            sigmoid_f := 2047;
        ELSIF x = 15079 THEN
            sigmoid_f := 2047;
        ELSIF x = 15080 THEN
            sigmoid_f := 2047;
        ELSIF x = 15081 THEN
            sigmoid_f := 2047;
        ELSIF x = 15082 THEN
            sigmoid_f := 2047;
        ELSIF x = 15083 THEN
            sigmoid_f := 2047;
        ELSIF x = 15084 THEN
            sigmoid_f := 2047;
        ELSIF x = 15085 THEN
            sigmoid_f := 2047;
        ELSIF x = 15086 THEN
            sigmoid_f := 2047;
        ELSIF x = 15087 THEN
            sigmoid_f := 2047;
        ELSIF x = 15088 THEN
            sigmoid_f := 2047;
        ELSIF x = 15089 THEN
            sigmoid_f := 2047;
        ELSIF x = 15090 THEN
            sigmoid_f := 2047;
        ELSIF x = 15091 THEN
            sigmoid_f := 2047;
        ELSIF x = 15092 THEN
            sigmoid_f := 2047;
        ELSIF x = 15093 THEN
            sigmoid_f := 2047;
        ELSIF x = 15094 THEN
            sigmoid_f := 2047;
        ELSIF x = 15095 THEN
            sigmoid_f := 2047;
        ELSIF x = 15096 THEN
            sigmoid_f := 2047;
        ELSIF x = 15097 THEN
            sigmoid_f := 2047;
        ELSIF x = 15098 THEN
            sigmoid_f := 2047;
        ELSIF x = 15099 THEN
            sigmoid_f := 2047;
        ELSIF x = 15100 THEN
            sigmoid_f := 2047;
        ELSIF x = 15101 THEN
            sigmoid_f := 2047;
        ELSIF x = 15102 THEN
            sigmoid_f := 2047;
        ELSIF x = 15103 THEN
            sigmoid_f := 2047;
        ELSIF x = 15104 THEN
            sigmoid_f := 2047;
        ELSIF x = 15105 THEN
            sigmoid_f := 2047;
        ELSIF x = 15106 THEN
            sigmoid_f := 2047;
        ELSIF x = 15107 THEN
            sigmoid_f := 2047;
        ELSIF x = 15108 THEN
            sigmoid_f := 2047;
        ELSIF x = 15109 THEN
            sigmoid_f := 2047;
        ELSIF x = 15110 THEN
            sigmoid_f := 2047;
        ELSIF x = 15111 THEN
            sigmoid_f := 2047;
        ELSIF x = 15112 THEN
            sigmoid_f := 2047;
        ELSIF x = 15113 THEN
            sigmoid_f := 2047;
        ELSIF x = 15114 THEN
            sigmoid_f := 2047;
        ELSIF x = 15115 THEN
            sigmoid_f := 2047;
        ELSIF x = 15116 THEN
            sigmoid_f := 2047;
        ELSIF x = 15117 THEN
            sigmoid_f := 2047;
        ELSIF x = 15118 THEN
            sigmoid_f := 2047;
        ELSIF x = 15119 THEN
            sigmoid_f := 2047;
        ELSIF x = 15120 THEN
            sigmoid_f := 2047;
        ELSIF x = 15121 THEN
            sigmoid_f := 2047;
        ELSIF x = 15122 THEN
            sigmoid_f := 2047;
        ELSIF x = 15123 THEN
            sigmoid_f := 2047;
        ELSIF x = 15124 THEN
            sigmoid_f := 2047;
        ELSIF x = 15125 THEN
            sigmoid_f := 2047;
        ELSIF x = 15126 THEN
            sigmoid_f := 2047;
        ELSIF x = 15127 THEN
            sigmoid_f := 2047;
        ELSIF x = 15128 THEN
            sigmoid_f := 2047;
        ELSIF x = 15129 THEN
            sigmoid_f := 2047;
        ELSIF x = 15130 THEN
            sigmoid_f := 2047;
        ELSIF x = 15131 THEN
            sigmoid_f := 2047;
        ELSIF x = 15132 THEN
            sigmoid_f := 2047;
        ELSIF x = 15133 THEN
            sigmoid_f := 2047;
        ELSIF x = 15134 THEN
            sigmoid_f := 2047;
        ELSIF x = 15135 THEN
            sigmoid_f := 2047;
        ELSIF x = 15136 THEN
            sigmoid_f := 2047;
        ELSIF x = 15137 THEN
            sigmoid_f := 2047;
        ELSIF x = 15138 THEN
            sigmoid_f := 2047;
        ELSIF x = 15139 THEN
            sigmoid_f := 2047;
        ELSIF x = 15140 THEN
            sigmoid_f := 2047;
        ELSIF x = 15141 THEN
            sigmoid_f := 2047;
        ELSIF x = 15142 THEN
            sigmoid_f := 2047;
        ELSIF x = 15143 THEN
            sigmoid_f := 2047;
        ELSIF x = 15144 THEN
            sigmoid_f := 2047;
        ELSIF x = 15145 THEN
            sigmoid_f := 2047;
        ELSIF x = 15146 THEN
            sigmoid_f := 2047;
        ELSIF x = 15147 THEN
            sigmoid_f := 2047;
        ELSIF x = 15148 THEN
            sigmoid_f := 2047;
        ELSIF x = 15149 THEN
            sigmoid_f := 2047;
        ELSIF x = 15150 THEN
            sigmoid_f := 2047;
        ELSIF x = 15151 THEN
            sigmoid_f := 2047;
        ELSIF x = 15152 THEN
            sigmoid_f := 2047;
        ELSIF x = 15153 THEN
            sigmoid_f := 2047;
        ELSIF x = 15154 THEN
            sigmoid_f := 2047;
        ELSIF x = 15155 THEN
            sigmoid_f := 2047;
        ELSIF x = 15156 THEN
            sigmoid_f := 2047;
        ELSIF x = 15157 THEN
            sigmoid_f := 2047;
        ELSIF x = 15158 THEN
            sigmoid_f := 2047;
        ELSIF x = 15159 THEN
            sigmoid_f := 2047;
        ELSIF x = 15160 THEN
            sigmoid_f := 2047;
        ELSIF x = 15161 THEN
            sigmoid_f := 2047;
        ELSIF x = 15162 THEN
            sigmoid_f := 2047;
        ELSIF x = 15163 THEN
            sigmoid_f := 2047;
        ELSIF x = 15164 THEN
            sigmoid_f := 2047;
        ELSIF x = 15165 THEN
            sigmoid_f := 2047;
        ELSIF x = 15166 THEN
            sigmoid_f := 2047;
        ELSIF x = 15167 THEN
            sigmoid_f := 2047;
        ELSIF x = 15168 THEN
            sigmoid_f := 2047;
        ELSIF x = 15169 THEN
            sigmoid_f := 2047;
        ELSIF x = 15170 THEN
            sigmoid_f := 2047;
        ELSIF x = 15171 THEN
            sigmoid_f := 2047;
        ELSIF x = 15172 THEN
            sigmoid_f := 2047;
        ELSIF x = 15173 THEN
            sigmoid_f := 2047;
        ELSIF x = 15174 THEN
            sigmoid_f := 2047;
        ELSIF x = 15175 THEN
            sigmoid_f := 2047;
        ELSIF x = 15176 THEN
            sigmoid_f := 2047;
        ELSIF x = 15177 THEN
            sigmoid_f := 2047;
        ELSIF x = 15178 THEN
            sigmoid_f := 2047;
        ELSIF x = 15179 THEN
            sigmoid_f := 2047;
        ELSIF x = 15180 THEN
            sigmoid_f := 2047;
        ELSIF x = 15181 THEN
            sigmoid_f := 2047;
        ELSIF x = 15182 THEN
            sigmoid_f := 2047;
        ELSIF x = 15183 THEN
            sigmoid_f := 2047;
        ELSIF x = 15184 THEN
            sigmoid_f := 2047;
        ELSIF x = 15185 THEN
            sigmoid_f := 2047;
        ELSIF x = 15186 THEN
            sigmoid_f := 2047;
        ELSIF x = 15187 THEN
            sigmoid_f := 2047;
        ELSIF x = 15188 THEN
            sigmoid_f := 2047;
        ELSIF x = 15189 THEN
            sigmoid_f := 2047;
        ELSIF x = 15190 THEN
            sigmoid_f := 2047;
        ELSIF x = 15191 THEN
            sigmoid_f := 2047;
        ELSIF x = 15192 THEN
            sigmoid_f := 2047;
        ELSIF x = 15193 THEN
            sigmoid_f := 2047;
        ELSIF x = 15194 THEN
            sigmoid_f := 2047;
        ELSIF x = 15195 THEN
            sigmoid_f := 2047;
        ELSIF x = 15196 THEN
            sigmoid_f := 2047;
        ELSIF x = 15197 THEN
            sigmoid_f := 2047;
        ELSIF x = 15198 THEN
            sigmoid_f := 2047;
        ELSIF x = 15199 THEN
            sigmoid_f := 2047;
        ELSIF x = 15200 THEN
            sigmoid_f := 2047;
        ELSIF x = 15201 THEN
            sigmoid_f := 2047;
        ELSIF x = 15202 THEN
            sigmoid_f := 2047;
        ELSIF x = 15203 THEN
            sigmoid_f := 2047;
        ELSIF x = 15204 THEN
            sigmoid_f := 2047;
        ELSIF x = 15205 THEN
            sigmoid_f := 2047;
        ELSIF x = 15206 THEN
            sigmoid_f := 2047;
        ELSIF x = 15207 THEN
            sigmoid_f := 2047;
        ELSIF x = 15208 THEN
            sigmoid_f := 2047;
        ELSIF x = 15209 THEN
            sigmoid_f := 2047;
        ELSIF x = 15210 THEN
            sigmoid_f := 2047;
        ELSIF x = 15211 THEN
            sigmoid_f := 2047;
        ELSIF x = 15212 THEN
            sigmoid_f := 2047;
        ELSIF x = 15213 THEN
            sigmoid_f := 2047;
        ELSIF x = 15214 THEN
            sigmoid_f := 2047;
        ELSIF x = 15215 THEN
            sigmoid_f := 2047;
        ELSIF x = 15216 THEN
            sigmoid_f := 2047;
        ELSIF x = 15217 THEN
            sigmoid_f := 2047;
        ELSIF x = 15218 THEN
            sigmoid_f := 2047;
        ELSIF x = 15219 THEN
            sigmoid_f := 2047;
        ELSIF x = 15220 THEN
            sigmoid_f := 2047;
        ELSIF x = 15221 THEN
            sigmoid_f := 2047;
        ELSIF x = 15222 THEN
            sigmoid_f := 2047;
        ELSIF x = 15223 THEN
            sigmoid_f := 2047;
        ELSIF x = 15224 THEN
            sigmoid_f := 2047;
        ELSIF x = 15225 THEN
            sigmoid_f := 2047;
        ELSIF x = 15226 THEN
            sigmoid_f := 2047;
        ELSIF x = 15227 THEN
            sigmoid_f := 2047;
        ELSIF x = 15228 THEN
            sigmoid_f := 2047;
        ELSIF x = 15229 THEN
            sigmoid_f := 2047;
        ELSIF x = 15230 THEN
            sigmoid_f := 2047;
        ELSIF x = 15231 THEN
            sigmoid_f := 2047;
        ELSIF x = 15232 THEN
            sigmoid_f := 2047;
        ELSIF x = 15233 THEN
            sigmoid_f := 2047;
        ELSIF x = 15234 THEN
            sigmoid_f := 2047;
        ELSIF x = 15235 THEN
            sigmoid_f := 2047;
        ELSIF x = 15236 THEN
            sigmoid_f := 2047;
        ELSIF x = 15237 THEN
            sigmoid_f := 2047;
        ELSIF x = 15238 THEN
            sigmoid_f := 2047;
        ELSIF x = 15239 THEN
            sigmoid_f := 2047;
        ELSIF x = 15240 THEN
            sigmoid_f := 2047;
        ELSIF x = 15241 THEN
            sigmoid_f := 2047;
        ELSIF x = 15242 THEN
            sigmoid_f := 2047;
        ELSIF x = 15243 THEN
            sigmoid_f := 2047;
        ELSIF x = 15244 THEN
            sigmoid_f := 2047;
        ELSIF x = 15245 THEN
            sigmoid_f := 2047;
        ELSIF x = 15246 THEN
            sigmoid_f := 2047;
        ELSIF x = 15247 THEN
            sigmoid_f := 2047;
        ELSIF x = 15248 THEN
            sigmoid_f := 2047;
        ELSIF x = 15249 THEN
            sigmoid_f := 2047;
        ELSIF x = 15250 THEN
            sigmoid_f := 2047;
        ELSIF x = 15251 THEN
            sigmoid_f := 2047;
        ELSIF x = 15252 THEN
            sigmoid_f := 2047;
        ELSIF x = 15253 THEN
            sigmoid_f := 2047;
        ELSIF x = 15254 THEN
            sigmoid_f := 2047;
        ELSIF x = 15255 THEN
            sigmoid_f := 2047;
        ELSIF x = 15256 THEN
            sigmoid_f := 2047;
        ELSIF x = 15257 THEN
            sigmoid_f := 2047;
        ELSIF x = 15258 THEN
            sigmoid_f := 2047;
        ELSIF x = 15259 THEN
            sigmoid_f := 2047;
        ELSIF x = 15260 THEN
            sigmoid_f := 2047;
        ELSIF x = 15261 THEN
            sigmoid_f := 2047;
        ELSIF x = 15262 THEN
            sigmoid_f := 2047;
        ELSIF x = 15263 THEN
            sigmoid_f := 2047;
        ELSIF x = 15264 THEN
            sigmoid_f := 2047;
        ELSIF x = 15265 THEN
            sigmoid_f := 2047;
        ELSIF x = 15266 THEN
            sigmoid_f := 2047;
        ELSIF x = 15267 THEN
            sigmoid_f := 2047;
        ELSIF x = 15268 THEN
            sigmoid_f := 2047;
        ELSIF x = 15269 THEN
            sigmoid_f := 2047;
        ELSIF x = 15270 THEN
            sigmoid_f := 2047;
        ELSIF x = 15271 THEN
            sigmoid_f := 2047;
        ELSIF x = 15272 THEN
            sigmoid_f := 2047;
        ELSIF x = 15273 THEN
            sigmoid_f := 2047;
        ELSIF x = 15274 THEN
            sigmoid_f := 2047;
        ELSIF x = 15275 THEN
            sigmoid_f := 2047;
        ELSIF x = 15276 THEN
            sigmoid_f := 2047;
        ELSIF x = 15277 THEN
            sigmoid_f := 2047;
        ELSIF x = 15278 THEN
            sigmoid_f := 2047;
        ELSIF x = 15279 THEN
            sigmoid_f := 2047;
        ELSIF x = 15280 THEN
            sigmoid_f := 2047;
        ELSIF x = 15281 THEN
            sigmoid_f := 2047;
        ELSIF x = 15282 THEN
            sigmoid_f := 2047;
        ELSIF x = 15283 THEN
            sigmoid_f := 2047;
        ELSIF x = 15284 THEN
            sigmoid_f := 2047;
        ELSIF x = 15285 THEN
            sigmoid_f := 2047;
        ELSIF x = 15286 THEN
            sigmoid_f := 2047;
        ELSIF x = 15287 THEN
            sigmoid_f := 2047;
        ELSIF x = 15288 THEN
            sigmoid_f := 2047;
        ELSIF x = 15289 THEN
            sigmoid_f := 2047;
        ELSIF x = 15290 THEN
            sigmoid_f := 2047;
        ELSIF x = 15291 THEN
            sigmoid_f := 2047;
        ELSIF x = 15292 THEN
            sigmoid_f := 2047;
        ELSIF x = 15293 THEN
            sigmoid_f := 2047;
        ELSIF x = 15294 THEN
            sigmoid_f := 2047;
        ELSIF x = 15295 THEN
            sigmoid_f := 2047;
        ELSIF x = 15296 THEN
            sigmoid_f := 2047;
        ELSIF x = 15297 THEN
            sigmoid_f := 2047;
        ELSIF x = 15298 THEN
            sigmoid_f := 2047;
        ELSIF x = 15299 THEN
            sigmoid_f := 2047;
        ELSIF x = 15300 THEN
            sigmoid_f := 2047;
        ELSIF x = 15301 THEN
            sigmoid_f := 2047;
        ELSIF x = 15302 THEN
            sigmoid_f := 2047;
        ELSIF x = 15303 THEN
            sigmoid_f := 2047;
        ELSIF x = 15304 THEN
            sigmoid_f := 2047;
        ELSIF x = 15305 THEN
            sigmoid_f := 2047;
        ELSIF x = 15306 THEN
            sigmoid_f := 2047;
        ELSIF x = 15307 THEN
            sigmoid_f := 2047;
        ELSIF x = 15308 THEN
            sigmoid_f := 2047;
        ELSIF x = 15309 THEN
            sigmoid_f := 2047;
        ELSIF x = 15310 THEN
            sigmoid_f := 2047;
        ELSIF x = 15311 THEN
            sigmoid_f := 2047;
        ELSIF x = 15312 THEN
            sigmoid_f := 2047;
        ELSIF x = 15313 THEN
            sigmoid_f := 2047;
        ELSIF x = 15314 THEN
            sigmoid_f := 2047;
        ELSIF x = 15315 THEN
            sigmoid_f := 2047;
        ELSIF x = 15316 THEN
            sigmoid_f := 2047;
        ELSIF x = 15317 THEN
            sigmoid_f := 2047;
        ELSIF x = 15318 THEN
            sigmoid_f := 2047;
        ELSIF x = 15319 THEN
            sigmoid_f := 2047;
        ELSIF x = 15320 THEN
            sigmoid_f := 2047;
        ELSIF x = 15321 THEN
            sigmoid_f := 2047;
        ELSIF x = 15322 THEN
            sigmoid_f := 2047;
        ELSIF x = 15323 THEN
            sigmoid_f := 2047;
        ELSIF x = 15324 THEN
            sigmoid_f := 2047;
        ELSIF x = 15325 THEN
            sigmoid_f := 2047;
        ELSIF x = 15326 THEN
            sigmoid_f := 2047;
        ELSIF x = 15327 THEN
            sigmoid_f := 2047;
        ELSIF x = 15328 THEN
            sigmoid_f := 2047;
        ELSIF x = 15329 THEN
            sigmoid_f := 2047;
        ELSIF x = 15330 THEN
            sigmoid_f := 2047;
        ELSIF x = 15331 THEN
            sigmoid_f := 2047;
        ELSIF x = 15332 THEN
            sigmoid_f := 2047;
        ELSIF x = 15333 THEN
            sigmoid_f := 2047;
        ELSIF x = 15334 THEN
            sigmoid_f := 2047;
        ELSIF x = 15335 THEN
            sigmoid_f := 2047;
        ELSIF x = 15336 THEN
            sigmoid_f := 2047;
        ELSIF x = 15337 THEN
            sigmoid_f := 2047;
        ELSIF x = 15338 THEN
            sigmoid_f := 2047;
        ELSIF x = 15339 THEN
            sigmoid_f := 2047;
        ELSIF x = 15340 THEN
            sigmoid_f := 2047;
        ELSIF x = 15341 THEN
            sigmoid_f := 2047;
        ELSIF x = 15342 THEN
            sigmoid_f := 2047;
        ELSIF x = 15343 THEN
            sigmoid_f := 2047;
        ELSIF x = 15344 THEN
            sigmoid_f := 2047;
        ELSIF x = 15345 THEN
            sigmoid_f := 2047;
        ELSIF x = 15346 THEN
            sigmoid_f := 2047;
        ELSIF x = 15347 THEN
            sigmoid_f := 2047;
        ELSIF x = 15348 THEN
            sigmoid_f := 2047;
        ELSIF x = 15349 THEN
            sigmoid_f := 2047;
        ELSIF x = 15350 THEN
            sigmoid_f := 2047;
        ELSIF x = 15351 THEN
            sigmoid_f := 2047;
        ELSIF x = 15352 THEN
            sigmoid_f := 2047;
        ELSIF x = 15353 THEN
            sigmoid_f := 2047;
        ELSIF x = 15354 THEN
            sigmoid_f := 2047;
        ELSIF x = 15355 THEN
            sigmoid_f := 2047;
        ELSIF x = 15356 THEN
            sigmoid_f := 2047;
        ELSIF x = 15357 THEN
            sigmoid_f := 2047;
        ELSIF x = 15358 THEN
            sigmoid_f := 2047;
        ELSIF x = 15359 THEN
            sigmoid_f := 2047;
        ELSIF x = 15360 THEN
            sigmoid_f := 2047;
        ELSIF x = 15361 THEN
            sigmoid_f := 2047;
        ELSIF x = 15362 THEN
            sigmoid_f := 2047;
        ELSIF x = 15363 THEN
            sigmoid_f := 2047;
        ELSIF x = 15364 THEN
            sigmoid_f := 2047;
        ELSIF x = 15365 THEN
            sigmoid_f := 2047;
        ELSIF x = 15366 THEN
            sigmoid_f := 2047;
        ELSIF x = 15367 THEN
            sigmoid_f := 2047;
        ELSIF x = 15368 THEN
            sigmoid_f := 2047;
        ELSIF x = 15369 THEN
            sigmoid_f := 2047;
        ELSIF x = 15370 THEN
            sigmoid_f := 2047;
        ELSIF x = 15371 THEN
            sigmoid_f := 2047;
        ELSIF x = 15372 THEN
            sigmoid_f := 2047;
        ELSIF x = 15373 THEN
            sigmoid_f := 2047;
        ELSIF x = 15374 THEN
            sigmoid_f := 2047;
        ELSIF x = 15375 THEN
            sigmoid_f := 2047;
        ELSIF x = 15376 THEN
            sigmoid_f := 2047;
        ELSIF x = 15377 THEN
            sigmoid_f := 2047;
        ELSIF x = 15378 THEN
            sigmoid_f := 2047;
        ELSIF x = 15379 THEN
            sigmoid_f := 2047;
        ELSIF x = 15380 THEN
            sigmoid_f := 2047;
        ELSIF x = 15381 THEN
            sigmoid_f := 2047;
        ELSIF x = 15382 THEN
            sigmoid_f := 2047;
        ELSIF x = 15383 THEN
            sigmoid_f := 2047;
        ELSIF x = 15384 THEN
            sigmoid_f := 2047;
        ELSIF x = 15385 THEN
            sigmoid_f := 2047;
        ELSIF x = 15386 THEN
            sigmoid_f := 2047;
        ELSIF x = 15387 THEN
            sigmoid_f := 2047;
        ELSIF x = 15388 THEN
            sigmoid_f := 2047;
        ELSIF x = 15389 THEN
            sigmoid_f := 2047;
        ELSIF x = 15390 THEN
            sigmoid_f := 2047;
        ELSIF x = 15391 THEN
            sigmoid_f := 2047;
        ELSIF x = 15392 THEN
            sigmoid_f := 2047;
        ELSIF x = 15393 THEN
            sigmoid_f := 2047;
        ELSIF x = 15394 THEN
            sigmoid_f := 2047;
        ELSIF x = 15395 THEN
            sigmoid_f := 2047;
        ELSIF x = 15396 THEN
            sigmoid_f := 2047;
        ELSIF x = 15397 THEN
            sigmoid_f := 2047;
        ELSIF x = 15398 THEN
            sigmoid_f := 2047;
        ELSIF x = 15399 THEN
            sigmoid_f := 2047;
        ELSIF x = 15400 THEN
            sigmoid_f := 2047;
        ELSIF x = 15401 THEN
            sigmoid_f := 2047;
        ELSIF x = 15402 THEN
            sigmoid_f := 2047;
        ELSIF x = 15403 THEN
            sigmoid_f := 2047;
        ELSIF x = 15404 THEN
            sigmoid_f := 2047;
        ELSIF x = 15405 THEN
            sigmoid_f := 2047;
        ELSIF x = 15406 THEN
            sigmoid_f := 2047;
        ELSIF x = 15407 THEN
            sigmoid_f := 2047;
        ELSIF x = 15408 THEN
            sigmoid_f := 2047;
        ELSIF x = 15409 THEN
            sigmoid_f := 2047;
        ELSIF x = 15410 THEN
            sigmoid_f := 2047;
        ELSIF x = 15411 THEN
            sigmoid_f := 2047;
        ELSIF x = 15412 THEN
            sigmoid_f := 2047;
        ELSIF x = 15413 THEN
            sigmoid_f := 2047;
        ELSIF x = 15414 THEN
            sigmoid_f := 2047;
        ELSIF x = 15415 THEN
            sigmoid_f := 2047;
        ELSIF x = 15416 THEN
            sigmoid_f := 2047;
        ELSIF x = 15417 THEN
            sigmoid_f := 2047;
        ELSIF x = 15418 THEN
            sigmoid_f := 2047;
        ELSIF x = 15419 THEN
            sigmoid_f := 2047;
        ELSIF x = 15420 THEN
            sigmoid_f := 2047;
        ELSIF x = 15421 THEN
            sigmoid_f := 2047;
        ELSIF x = 15422 THEN
            sigmoid_f := 2047;
        ELSIF x = 15423 THEN
            sigmoid_f := 2047;
        ELSIF x = 15424 THEN
            sigmoid_f := 2047;
        ELSIF x = 15425 THEN
            sigmoid_f := 2047;
        ELSIF x = 15426 THEN
            sigmoid_f := 2047;
        ELSIF x = 15427 THEN
            sigmoid_f := 2047;
        ELSIF x = 15428 THEN
            sigmoid_f := 2047;
        ELSIF x = 15429 THEN
            sigmoid_f := 2047;
        ELSIF x = 15430 THEN
            sigmoid_f := 2047;
        ELSIF x = 15431 THEN
            sigmoid_f := 2047;
        ELSIF x = 15432 THEN
            sigmoid_f := 2047;
        ELSIF x = 15433 THEN
            sigmoid_f := 2047;
        ELSIF x = 15434 THEN
            sigmoid_f := 2047;
        ELSIF x = 15435 THEN
            sigmoid_f := 2047;
        ELSIF x = 15436 THEN
            sigmoid_f := 2047;
        ELSIF x = 15437 THEN
            sigmoid_f := 2047;
        ELSIF x = 15438 THEN
            sigmoid_f := 2047;
        ELSIF x = 15439 THEN
            sigmoid_f := 2047;
        ELSIF x = 15440 THEN
            sigmoid_f := 2047;
        ELSIF x = 15441 THEN
            sigmoid_f := 2047;
        ELSIF x = 15442 THEN
            sigmoid_f := 2047;
        ELSIF x = 15443 THEN
            sigmoid_f := 2047;
        ELSIF x = 15444 THEN
            sigmoid_f := 2047;
        ELSIF x = 15445 THEN
            sigmoid_f := 2047;
        ELSIF x = 15446 THEN
            sigmoid_f := 2047;
        ELSIF x = 15447 THEN
            sigmoid_f := 2047;
        ELSIF x = 15448 THEN
            sigmoid_f := 2047;
        ELSIF x = 15449 THEN
            sigmoid_f := 2047;
        ELSIF x = 15450 THEN
            sigmoid_f := 2047;
        ELSIF x = 15451 THEN
            sigmoid_f := 2047;
        ELSIF x = 15452 THEN
            sigmoid_f := 2047;
        ELSIF x = 15453 THEN
            sigmoid_f := 2047;
        ELSIF x = 15454 THEN
            sigmoid_f := 2047;
        ELSIF x = 15455 THEN
            sigmoid_f := 2047;
        ELSIF x = 15456 THEN
            sigmoid_f := 2047;
        ELSIF x = 15457 THEN
            sigmoid_f := 2047;
        ELSIF x = 15458 THEN
            sigmoid_f := 2047;
        ELSIF x = 15459 THEN
            sigmoid_f := 2047;
        ELSIF x = 15460 THEN
            sigmoid_f := 2047;
        ELSIF x = 15461 THEN
            sigmoid_f := 2047;
        ELSIF x = 15462 THEN
            sigmoid_f := 2047;
        ELSIF x = 15463 THEN
            sigmoid_f := 2047;
        ELSIF x = 15464 THEN
            sigmoid_f := 2047;
        ELSIF x = 15465 THEN
            sigmoid_f := 2047;
        ELSIF x = 15466 THEN
            sigmoid_f := 2047;
        ELSIF x = 15467 THEN
            sigmoid_f := 2047;
        ELSIF x = 15468 THEN
            sigmoid_f := 2047;
        ELSIF x = 15469 THEN
            sigmoid_f := 2047;
        ELSIF x = 15470 THEN
            sigmoid_f := 2047;
        ELSIF x = 15471 THEN
            sigmoid_f := 2047;
        ELSIF x = 15472 THEN
            sigmoid_f := 2047;
        ELSIF x = 15473 THEN
            sigmoid_f := 2047;
        ELSIF x = 15474 THEN
            sigmoid_f := 2047;
        ELSIF x = 15475 THEN
            sigmoid_f := 2047;
        ELSIF x = 15476 THEN
            sigmoid_f := 2047;
        ELSIF x = 15477 THEN
            sigmoid_f := 2047;
        ELSIF x = 15478 THEN
            sigmoid_f := 2047;
        ELSIF x = 15479 THEN
            sigmoid_f := 2047;
        ELSIF x = 15480 THEN
            sigmoid_f := 2047;
        ELSIF x = 15481 THEN
            sigmoid_f := 2047;
        ELSIF x = 15482 THEN
            sigmoid_f := 2047;
        ELSIF x = 15483 THEN
            sigmoid_f := 2047;
        ELSIF x = 15484 THEN
            sigmoid_f := 2047;
        ELSIF x = 15485 THEN
            sigmoid_f := 2047;
        ELSIF x = 15486 THEN
            sigmoid_f := 2047;
        ELSIF x = 15487 THEN
            sigmoid_f := 2047;
        ELSIF x = 15488 THEN
            sigmoid_f := 2047;
        ELSIF x = 15489 THEN
            sigmoid_f := 2047;
        ELSIF x = 15490 THEN
            sigmoid_f := 2047;
        ELSIF x = 15491 THEN
            sigmoid_f := 2047;
        ELSIF x = 15492 THEN
            sigmoid_f := 2047;
        ELSIF x = 15493 THEN
            sigmoid_f := 2047;
        ELSIF x = 15494 THEN
            sigmoid_f := 2047;
        ELSIF x = 15495 THEN
            sigmoid_f := 2047;
        ELSIF x = 15496 THEN
            sigmoid_f := 2047;
        ELSIF x = 15497 THEN
            sigmoid_f := 2047;
        ELSIF x = 15498 THEN
            sigmoid_f := 2047;
        ELSIF x = 15499 THEN
            sigmoid_f := 2047;
        ELSIF x = 15500 THEN
            sigmoid_f := 2047;
        ELSIF x = 15501 THEN
            sigmoid_f := 2047;
        ELSIF x = 15502 THEN
            sigmoid_f := 2047;
        ELSIF x = 15503 THEN
            sigmoid_f := 2047;
        ELSIF x = 15504 THEN
            sigmoid_f := 2047;
        ELSIF x = 15505 THEN
            sigmoid_f := 2047;
        ELSIF x = 15506 THEN
            sigmoid_f := 2047;
        ELSIF x = 15507 THEN
            sigmoid_f := 2047;
        ELSIF x = 15508 THEN
            sigmoid_f := 2047;
        ELSIF x = 15509 THEN
            sigmoid_f := 2047;
        ELSIF x = 15510 THEN
            sigmoid_f := 2047;
        ELSIF x = 15511 THEN
            sigmoid_f := 2047;
        ELSIF x = 15512 THEN
            sigmoid_f := 2047;
        ELSIF x = 15513 THEN
            sigmoid_f := 2047;
        ELSIF x = 15514 THEN
            sigmoid_f := 2047;
        ELSIF x = 15515 THEN
            sigmoid_f := 2047;
        ELSIF x = 15516 THEN
            sigmoid_f := 2047;
        ELSIF x = 15517 THEN
            sigmoid_f := 2047;
        ELSIF x = 15518 THEN
            sigmoid_f := 2047;
        ELSIF x = 15519 THEN
            sigmoid_f := 2047;
        ELSIF x = 15520 THEN
            sigmoid_f := 2047;
        ELSIF x = 15521 THEN
            sigmoid_f := 2047;
        ELSIF x = 15522 THEN
            sigmoid_f := 2047;
        ELSIF x = 15523 THEN
            sigmoid_f := 2047;
        ELSIF x = 15524 THEN
            sigmoid_f := 2047;
        ELSIF x = 15525 THEN
            sigmoid_f := 2047;
        ELSIF x = 15526 THEN
            sigmoid_f := 2047;
        ELSIF x = 15527 THEN
            sigmoid_f := 2047;
        ELSIF x = 15528 THEN
            sigmoid_f := 2047;
        ELSIF x = 15529 THEN
            sigmoid_f := 2047;
        ELSIF x = 15530 THEN
            sigmoid_f := 2047;
        ELSIF x = 15531 THEN
            sigmoid_f := 2047;
        ELSIF x = 15532 THEN
            sigmoid_f := 2047;
        ELSIF x = 15533 THEN
            sigmoid_f := 2047;
        ELSIF x = 15534 THEN
            sigmoid_f := 2047;
        ELSIF x = 15535 THEN
            sigmoid_f := 2047;
        ELSIF x = 15536 THEN
            sigmoid_f := 2047;
        ELSIF x = 15537 THEN
            sigmoid_f := 2047;
        ELSIF x = 15538 THEN
            sigmoid_f := 2047;
        ELSIF x = 15539 THEN
            sigmoid_f := 2047;
        ELSIF x = 15540 THEN
            sigmoid_f := 2047;
        ELSIF x = 15541 THEN
            sigmoid_f := 2047;
        ELSIF x = 15542 THEN
            sigmoid_f := 2047;
        ELSIF x = 15543 THEN
            sigmoid_f := 2047;
        ELSIF x = 15544 THEN
            sigmoid_f := 2047;
        ELSIF x = 15545 THEN
            sigmoid_f := 2047;
        ELSIF x = 15546 THEN
            sigmoid_f := 2047;
        ELSIF x = 15547 THEN
            sigmoid_f := 2047;
        ELSIF x = 15548 THEN
            sigmoid_f := 2047;
        ELSIF x = 15549 THEN
            sigmoid_f := 2047;
        ELSIF x = 15550 THEN
            sigmoid_f := 2047;
        ELSIF x = 15551 THEN
            sigmoid_f := 2047;
        ELSIF x = 15552 THEN
            sigmoid_f := 2047;
        ELSIF x = 15553 THEN
            sigmoid_f := 2047;
        ELSIF x = 15554 THEN
            sigmoid_f := 2047;
        ELSIF x = 15555 THEN
            sigmoid_f := 2047;
        ELSIF x = 15556 THEN
            sigmoid_f := 2047;
        ELSIF x = 15557 THEN
            sigmoid_f := 2047;
        ELSIF x = 15558 THEN
            sigmoid_f := 2047;
        ELSIF x = 15559 THEN
            sigmoid_f := 2047;
        ELSIF x = 15560 THEN
            sigmoid_f := 2047;
        ELSIF x = 15561 THEN
            sigmoid_f := 2047;
        ELSIF x = 15562 THEN
            sigmoid_f := 2047;
        ELSIF x = 15563 THEN
            sigmoid_f := 2047;
        ELSIF x = 15564 THEN
            sigmoid_f := 2047;
        ELSIF x = 15565 THEN
            sigmoid_f := 2047;
        ELSIF x = 15566 THEN
            sigmoid_f := 2047;
        ELSIF x = 15567 THEN
            sigmoid_f := 2047;
        ELSIF x = 15568 THEN
            sigmoid_f := 2047;
        ELSIF x = 15569 THEN
            sigmoid_f := 2047;
        ELSIF x = 15570 THEN
            sigmoid_f := 2047;
        ELSIF x = 15571 THEN
            sigmoid_f := 2047;
        ELSIF x = 15572 THEN
            sigmoid_f := 2047;
        ELSIF x = 15573 THEN
            sigmoid_f := 2047;
        ELSIF x = 15574 THEN
            sigmoid_f := 2047;
        ELSIF x = 15575 THEN
            sigmoid_f := 2047;
        ELSIF x = 15576 THEN
            sigmoid_f := 2047;
        ELSIF x = 15577 THEN
            sigmoid_f := 2047;
        ELSIF x = 15578 THEN
            sigmoid_f := 2047;
        ELSIF x = 15579 THEN
            sigmoid_f := 2047;
        ELSIF x = 15580 THEN
            sigmoid_f := 2047;
        ELSIF x = 15581 THEN
            sigmoid_f := 2047;
        ELSIF x = 15582 THEN
            sigmoid_f := 2047;
        ELSIF x = 15583 THEN
            sigmoid_f := 2047;
        ELSIF x = 15584 THEN
            sigmoid_f := 2047;
        ELSIF x = 15585 THEN
            sigmoid_f := 2047;
        ELSIF x = 15586 THEN
            sigmoid_f := 2047;
        ELSIF x = 15587 THEN
            sigmoid_f := 2047;
        ELSIF x = 15588 THEN
            sigmoid_f := 2047;
        ELSIF x = 15589 THEN
            sigmoid_f := 2047;
        ELSIF x = 15590 THEN
            sigmoid_f := 2047;
        ELSIF x = 15591 THEN
            sigmoid_f := 2047;
        ELSIF x = 15592 THEN
            sigmoid_f := 2047;
        ELSIF x = 15593 THEN
            sigmoid_f := 2047;
        ELSIF x = 15594 THEN
            sigmoid_f := 2047;
        ELSIF x = 15595 THEN
            sigmoid_f := 2047;
        ELSIF x = 15596 THEN
            sigmoid_f := 2047;
        ELSIF x = 15597 THEN
            sigmoid_f := 2047;
        ELSIF x = 15598 THEN
            sigmoid_f := 2047;
        ELSIF x = 15599 THEN
            sigmoid_f := 2047;
        ELSIF x = 15600 THEN
            sigmoid_f := 2047;
        ELSIF x = 15601 THEN
            sigmoid_f := 2047;
        ELSIF x = 15602 THEN
            sigmoid_f := 2047;
        ELSIF x = 15603 THEN
            sigmoid_f := 2047;
        ELSIF x = 15604 THEN
            sigmoid_f := 2047;
        ELSIF x = 15605 THEN
            sigmoid_f := 2047;
        ELSIF x = 15606 THEN
            sigmoid_f := 2047;
        ELSIF x = 15607 THEN
            sigmoid_f := 2047;
        ELSIF x = 15608 THEN
            sigmoid_f := 2047;
        ELSIF x = 15609 THEN
            sigmoid_f := 2047;
        ELSIF x = 15610 THEN
            sigmoid_f := 2047;
        ELSIF x = 15611 THEN
            sigmoid_f := 2047;
        ELSIF x = 15612 THEN
            sigmoid_f := 2047;
        ELSIF x = 15613 THEN
            sigmoid_f := 2047;
        ELSIF x = 15614 THEN
            sigmoid_f := 2047;
        ELSIF x = 15615 THEN
            sigmoid_f := 2047;
        ELSIF x = 15616 THEN
            sigmoid_f := 2047;
        ELSIF x = 15617 THEN
            sigmoid_f := 2047;
        ELSIF x = 15618 THEN
            sigmoid_f := 2047;
        ELSIF x = 15619 THEN
            sigmoid_f := 2047;
        ELSIF x = 15620 THEN
            sigmoid_f := 2047;
        ELSIF x = 15621 THEN
            sigmoid_f := 2047;
        ELSIF x = 15622 THEN
            sigmoid_f := 2047;
        ELSIF x = 15623 THEN
            sigmoid_f := 2047;
        ELSIF x = 15624 THEN
            sigmoid_f := 2047;
        ELSIF x = 15625 THEN
            sigmoid_f := 2047;
        ELSIF x = 15626 THEN
            sigmoid_f := 2047;
        ELSIF x = 15627 THEN
            sigmoid_f := 2047;
        ELSIF x = 15628 THEN
            sigmoid_f := 2047;
        ELSIF x = 15629 THEN
            sigmoid_f := 2047;
        ELSIF x = 15630 THEN
            sigmoid_f := 2047;
        ELSIF x = 15631 THEN
            sigmoid_f := 2047;
        ELSIF x = 15632 THEN
            sigmoid_f := 2047;
        ELSIF x = 15633 THEN
            sigmoid_f := 2047;
        ELSIF x = 15634 THEN
            sigmoid_f := 2047;
        ELSIF x = 15635 THEN
            sigmoid_f := 2047;
        ELSIF x = 15636 THEN
            sigmoid_f := 2047;
        ELSIF x = 15637 THEN
            sigmoid_f := 2047;
        ELSIF x = 15638 THEN
            sigmoid_f := 2047;
        ELSIF x = 15639 THEN
            sigmoid_f := 2047;
        ELSIF x = 15640 THEN
            sigmoid_f := 2047;
        ELSIF x = 15641 THEN
            sigmoid_f := 2047;
        ELSIF x = 15642 THEN
            sigmoid_f := 2047;
        ELSIF x = 15643 THEN
            sigmoid_f := 2047;
        ELSIF x = 15644 THEN
            sigmoid_f := 2047;
        ELSIF x = 15645 THEN
            sigmoid_f := 2047;
        ELSIF x = 15646 THEN
            sigmoid_f := 2047;
        ELSIF x = 15647 THEN
            sigmoid_f := 2047;
        ELSIF x = 15648 THEN
            sigmoid_f := 2047;
        ELSIF x = 15649 THEN
            sigmoid_f := 2047;
        ELSIF x = 15650 THEN
            sigmoid_f := 2047;
        ELSIF x = 15651 THEN
            sigmoid_f := 2047;
        ELSIF x = 15652 THEN
            sigmoid_f := 2047;
        ELSIF x = 15653 THEN
            sigmoid_f := 2047;
        ELSIF x = 15654 THEN
            sigmoid_f := 2047;
        ELSIF x = 15655 THEN
            sigmoid_f := 2047;
        ELSIF x = 15656 THEN
            sigmoid_f := 2047;
        ELSIF x = 15657 THEN
            sigmoid_f := 2047;
        ELSIF x = 15658 THEN
            sigmoid_f := 2047;
        ELSIF x = 15659 THEN
            sigmoid_f := 2047;
        ELSIF x = 15660 THEN
            sigmoid_f := 2047;
        ELSIF x = 15661 THEN
            sigmoid_f := 2047;
        ELSIF x = 15662 THEN
            sigmoid_f := 2047;
        ELSIF x = 15663 THEN
            sigmoid_f := 2047;
        ELSIF x = 15664 THEN
            sigmoid_f := 2047;
        ELSIF x = 15665 THEN
            sigmoid_f := 2047;
        ELSIF x = 15666 THEN
            sigmoid_f := 2047;
        ELSIF x = 15667 THEN
            sigmoid_f := 2047;
        ELSIF x = 15668 THEN
            sigmoid_f := 2047;
        ELSIF x = 15669 THEN
            sigmoid_f := 2047;
        ELSIF x = 15670 THEN
            sigmoid_f := 2047;
        ELSIF x = 15671 THEN
            sigmoid_f := 2047;
        ELSIF x = 15672 THEN
            sigmoid_f := 2047;
        ELSIF x = 15673 THEN
            sigmoid_f := 2047;
        ELSIF x = 15674 THEN
            sigmoid_f := 2047;
        ELSIF x = 15675 THEN
            sigmoid_f := 2047;
        ELSIF x = 15676 THEN
            sigmoid_f := 2047;
        ELSIF x = 15677 THEN
            sigmoid_f := 2047;
        ELSIF x = 15678 THEN
            sigmoid_f := 2047;
        ELSIF x = 15679 THEN
            sigmoid_f := 2047;
        ELSIF x = 15680 THEN
            sigmoid_f := 2047;
        ELSIF x = 15681 THEN
            sigmoid_f := 2047;
        ELSIF x = 15682 THEN
            sigmoid_f := 2047;
        ELSIF x = 15683 THEN
            sigmoid_f := 2047;
        ELSIF x = 15684 THEN
            sigmoid_f := 2047;
        ELSIF x = 15685 THEN
            sigmoid_f := 2047;
        ELSIF x = 15686 THEN
            sigmoid_f := 2047;
        ELSIF x = 15687 THEN
            sigmoid_f := 2047;
        ELSIF x = 15688 THEN
            sigmoid_f := 2047;
        ELSIF x = 15689 THEN
            sigmoid_f := 2047;
        ELSIF x = 15690 THEN
            sigmoid_f := 2047;
        ELSIF x = 15691 THEN
            sigmoid_f := 2047;
        ELSIF x = 15692 THEN
            sigmoid_f := 2047;
        ELSIF x = 15693 THEN
            sigmoid_f := 2047;
        ELSIF x = 15694 THEN
            sigmoid_f := 2047;
        ELSIF x = 15695 THEN
            sigmoid_f := 2047;
        ELSIF x = 15696 THEN
            sigmoid_f := 2047;
        ELSIF x = 15697 THEN
            sigmoid_f := 2047;
        ELSIF x = 15698 THEN
            sigmoid_f := 2047;
        ELSIF x = 15699 THEN
            sigmoid_f := 2047;
        ELSIF x = 15700 THEN
            sigmoid_f := 2047;
        ELSIF x = 15701 THEN
            sigmoid_f := 2047;
        ELSIF x = 15702 THEN
            sigmoid_f := 2047;
        ELSIF x = 15703 THEN
            sigmoid_f := 2047;
        ELSIF x = 15704 THEN
            sigmoid_f := 2047;
        ELSIF x = 15705 THEN
            sigmoid_f := 2047;
        ELSIF x = 15706 THEN
            sigmoid_f := 2047;
        ELSIF x = 15707 THEN
            sigmoid_f := 2047;
        ELSIF x = 15708 THEN
            sigmoid_f := 2047;
        ELSIF x = 15709 THEN
            sigmoid_f := 2047;
        ELSIF x = 15710 THEN
            sigmoid_f := 2047;
        ELSIF x = 15711 THEN
            sigmoid_f := 2047;
        ELSIF x = 15712 THEN
            sigmoid_f := 2047;
        ELSIF x = 15713 THEN
            sigmoid_f := 2047;
        ELSIF x = 15714 THEN
            sigmoid_f := 2047;
        ELSIF x = 15715 THEN
            sigmoid_f := 2047;
        ELSIF x = 15716 THEN
            sigmoid_f := 2047;
        ELSIF x = 15717 THEN
            sigmoid_f := 2047;
        ELSIF x = 15718 THEN
            sigmoid_f := 2047;
        ELSIF x = 15719 THEN
            sigmoid_f := 2047;
        ELSIF x = 15720 THEN
            sigmoid_f := 2047;
        ELSIF x = 15721 THEN
            sigmoid_f := 2047;
        ELSIF x = 15722 THEN
            sigmoid_f := 2047;
        ELSIF x = 15723 THEN
            sigmoid_f := 2047;
        ELSIF x = 15724 THEN
            sigmoid_f := 2047;
        ELSIF x = 15725 THEN
            sigmoid_f := 2047;
        ELSIF x = 15726 THEN
            sigmoid_f := 2047;
        ELSIF x = 15727 THEN
            sigmoid_f := 2047;
        ELSIF x = 15728 THEN
            sigmoid_f := 2047;
        ELSIF x = 15729 THEN
            sigmoid_f := 2047;
        ELSIF x = 15730 THEN
            sigmoid_f := 2047;
        ELSIF x = 15731 THEN
            sigmoid_f := 2047;
        ELSIF x = 15732 THEN
            sigmoid_f := 2047;
        ELSIF x = 15733 THEN
            sigmoid_f := 2047;
        ELSIF x = 15734 THEN
            sigmoid_f := 2047;
        ELSIF x = 15735 THEN
            sigmoid_f := 2047;
        ELSIF x = 15736 THEN
            sigmoid_f := 2047;
        ELSIF x = 15737 THEN
            sigmoid_f := 2047;
        ELSIF x = 15738 THEN
            sigmoid_f := 2047;
        ELSIF x = 15739 THEN
            sigmoid_f := 2047;
        ELSIF x = 15740 THEN
            sigmoid_f := 2047;
        ELSIF x = 15741 THEN
            sigmoid_f := 2047;
        ELSIF x = 15742 THEN
            sigmoid_f := 2047;
        ELSIF x = 15743 THEN
            sigmoid_f := 2047;
        ELSIF x = 15744 THEN
            sigmoid_f := 2047;
        ELSIF x = 15745 THEN
            sigmoid_f := 2047;
        ELSIF x = 15746 THEN
            sigmoid_f := 2047;
        ELSIF x = 15747 THEN
            sigmoid_f := 2047;
        ELSIF x = 15748 THEN
            sigmoid_f := 2047;
        ELSIF x = 15749 THEN
            sigmoid_f := 2047;
        ELSIF x = 15750 THEN
            sigmoid_f := 2047;
        ELSIF x = 15751 THEN
            sigmoid_f := 2047;
        ELSIF x = 15752 THEN
            sigmoid_f := 2047;
        ELSIF x = 15753 THEN
            sigmoid_f := 2047;
        ELSIF x = 15754 THEN
            sigmoid_f := 2047;
        ELSIF x = 15755 THEN
            sigmoid_f := 2047;
        ELSIF x = 15756 THEN
            sigmoid_f := 2047;
        ELSIF x = 15757 THEN
            sigmoid_f := 2047;
        ELSIF x = 15758 THEN
            sigmoid_f := 2047;
        ELSIF x = 15759 THEN
            sigmoid_f := 2047;
        ELSIF x = 15760 THEN
            sigmoid_f := 2047;
        ELSIF x = 15761 THEN
            sigmoid_f := 2047;
        ELSIF x = 15762 THEN
            sigmoid_f := 2047;
        ELSIF x = 15763 THEN
            sigmoid_f := 2047;
        ELSIF x = 15764 THEN
            sigmoid_f := 2047;
        ELSIF x = 15765 THEN
            sigmoid_f := 2047;
        ELSIF x = 15766 THEN
            sigmoid_f := 2047;
        ELSIF x = 15767 THEN
            sigmoid_f := 2047;
        ELSIF x = 15768 THEN
            sigmoid_f := 2047;
        ELSIF x = 15769 THEN
            sigmoid_f := 2047;
        ELSIF x = 15770 THEN
            sigmoid_f := 2047;
        ELSIF x = 15771 THEN
            sigmoid_f := 2047;
        ELSIF x = 15772 THEN
            sigmoid_f := 2047;
        ELSIF x = 15773 THEN
            sigmoid_f := 2047;
        ELSIF x = 15774 THEN
            sigmoid_f := 2047;
        ELSIF x = 15775 THEN
            sigmoid_f := 2047;
        ELSIF x = 15776 THEN
            sigmoid_f := 2047;
        ELSIF x = 15777 THEN
            sigmoid_f := 2047;
        ELSIF x = 15778 THEN
            sigmoid_f := 2047;
        ELSIF x = 15779 THEN
            sigmoid_f := 2047;
        ELSIF x = 15780 THEN
            sigmoid_f := 2047;
        ELSIF x = 15781 THEN
            sigmoid_f := 2047;
        ELSIF x = 15782 THEN
            sigmoid_f := 2047;
        ELSIF x = 15783 THEN
            sigmoid_f := 2047;
        ELSIF x = 15784 THEN
            sigmoid_f := 2047;
        ELSIF x = 15785 THEN
            sigmoid_f := 2047;
        ELSIF x = 15786 THEN
            sigmoid_f := 2047;
        ELSIF x = 15787 THEN
            sigmoid_f := 2047;
        ELSIF x = 15788 THEN
            sigmoid_f := 2047;
        ELSIF x = 15789 THEN
            sigmoid_f := 2047;
        ELSIF x = 15790 THEN
            sigmoid_f := 2047;
        ELSIF x = 15791 THEN
            sigmoid_f := 2047;
        ELSIF x = 15792 THEN
            sigmoid_f := 2047;
        ELSIF x = 15793 THEN
            sigmoid_f := 2047;
        ELSIF x = 15794 THEN
            sigmoid_f := 2047;
        ELSIF x = 15795 THEN
            sigmoid_f := 2047;
        ELSIF x = 15796 THEN
            sigmoid_f := 2047;
        ELSIF x = 15797 THEN
            sigmoid_f := 2047;
        ELSIF x = 15798 THEN
            sigmoid_f := 2047;
        ELSIF x = 15799 THEN
            sigmoid_f := 2047;
        ELSIF x = 15800 THEN
            sigmoid_f := 2047;
        ELSIF x = 15801 THEN
            sigmoid_f := 2047;
        ELSIF x = 15802 THEN
            sigmoid_f := 2047;
        ELSIF x = 15803 THEN
            sigmoid_f := 2047;
        ELSIF x = 15804 THEN
            sigmoid_f := 2047;
        ELSIF x = 15805 THEN
            sigmoid_f := 2047;
        ELSIF x = 15806 THEN
            sigmoid_f := 2047;
        ELSIF x = 15807 THEN
            sigmoid_f := 2047;
        ELSIF x = 15808 THEN
            sigmoid_f := 2047;
        ELSIF x = 15809 THEN
            sigmoid_f := 2047;
        ELSIF x = 15810 THEN
            sigmoid_f := 2047;
        ELSIF x = 15811 THEN
            sigmoid_f := 2047;
        ELSIF x = 15812 THEN
            sigmoid_f := 2047;
        ELSIF x = 15813 THEN
            sigmoid_f := 2047;
        ELSIF x = 15814 THEN
            sigmoid_f := 2047;
        ELSIF x = 15815 THEN
            sigmoid_f := 2047;
        ELSIF x = 15816 THEN
            sigmoid_f := 2047;
        ELSIF x = 15817 THEN
            sigmoid_f := 2047;
        ELSIF x = 15818 THEN
            sigmoid_f := 2047;
        ELSIF x = 15819 THEN
            sigmoid_f := 2047;
        ELSIF x = 15820 THEN
            sigmoid_f := 2047;
        ELSIF x = 15821 THEN
            sigmoid_f := 2047;
        ELSIF x = 15822 THEN
            sigmoid_f := 2047;
        ELSIF x = 15823 THEN
            sigmoid_f := 2047;
        ELSIF x = 15824 THEN
            sigmoid_f := 2047;
        ELSIF x = 15825 THEN
            sigmoid_f := 2047;
        ELSIF x = 15826 THEN
            sigmoid_f := 2047;
        ELSIF x = 15827 THEN
            sigmoid_f := 2047;
        ELSIF x = 15828 THEN
            sigmoid_f := 2047;
        ELSIF x = 15829 THEN
            sigmoid_f := 2047;
        ELSIF x = 15830 THEN
            sigmoid_f := 2047;
        ELSIF x = 15831 THEN
            sigmoid_f := 2047;
        ELSIF x = 15832 THEN
            sigmoid_f := 2047;
        ELSIF x = 15833 THEN
            sigmoid_f := 2047;
        ELSIF x = 15834 THEN
            sigmoid_f := 2047;
        ELSIF x = 15835 THEN
            sigmoid_f := 2047;
        ELSIF x = 15836 THEN
            sigmoid_f := 2047;
        ELSIF x = 15837 THEN
            sigmoid_f := 2047;
        ELSIF x = 15838 THEN
            sigmoid_f := 2047;
        ELSIF x = 15839 THEN
            sigmoid_f := 2047;
        ELSIF x = 15840 THEN
            sigmoid_f := 2047;
        ELSIF x = 15841 THEN
            sigmoid_f := 2047;
        ELSIF x = 15842 THEN
            sigmoid_f := 2047;
        ELSIF x = 15843 THEN
            sigmoid_f := 2047;
        ELSIF x = 15844 THEN
            sigmoid_f := 2047;
        ELSIF x = 15845 THEN
            sigmoid_f := 2047;
        ELSIF x = 15846 THEN
            sigmoid_f := 2047;
        ELSIF x = 15847 THEN
            sigmoid_f := 2047;
        ELSIF x = 15848 THEN
            sigmoid_f := 2047;
        ELSIF x = 15849 THEN
            sigmoid_f := 2047;
        ELSIF x = 15850 THEN
            sigmoid_f := 2047;
        ELSIF x = 15851 THEN
            sigmoid_f := 2047;
        ELSIF x = 15852 THEN
            sigmoid_f := 2047;
        ELSIF x = 15853 THEN
            sigmoid_f := 2047;
        ELSIF x = 15854 THEN
            sigmoid_f := 2047;
        ELSIF x = 15855 THEN
            sigmoid_f := 2047;
        ELSIF x = 15856 THEN
            sigmoid_f := 2047;
        ELSIF x = 15857 THEN
            sigmoid_f := 2047;
        ELSIF x = 15858 THEN
            sigmoid_f := 2047;
        ELSIF x = 15859 THEN
            sigmoid_f := 2047;
        ELSIF x = 15860 THEN
            sigmoid_f := 2047;
        ELSIF x = 15861 THEN
            sigmoid_f := 2047;
        ELSIF x = 15862 THEN
            sigmoid_f := 2047;
        ELSIF x = 15863 THEN
            sigmoid_f := 2047;
        ELSIF x = 15864 THEN
            sigmoid_f := 2047;
        ELSIF x = 15865 THEN
            sigmoid_f := 2047;
        ELSIF x = 15866 THEN
            sigmoid_f := 2047;
        ELSIF x = 15867 THEN
            sigmoid_f := 2047;
        ELSIF x = 15868 THEN
            sigmoid_f := 2047;
        ELSIF x = 15869 THEN
            sigmoid_f := 2047;
        ELSIF x = 15870 THEN
            sigmoid_f := 2047;
        ELSIF x = 15871 THEN
            sigmoid_f := 2047;
        ELSIF x = 15872 THEN
            sigmoid_f := 2047;
        ELSIF x = 15873 THEN
            sigmoid_f := 2047;
        ELSIF x = 15874 THEN
            sigmoid_f := 2047;
        ELSIF x = 15875 THEN
            sigmoid_f := 2047;
        ELSIF x = 15876 THEN
            sigmoid_f := 2047;
        ELSIF x = 15877 THEN
            sigmoid_f := 2047;
        ELSIF x = 15878 THEN
            sigmoid_f := 2047;
        ELSIF x = 15879 THEN
            sigmoid_f := 2047;
        ELSIF x = 15880 THEN
            sigmoid_f := 2047;
        ELSIF x = 15881 THEN
            sigmoid_f := 2047;
        ELSIF x = 15882 THEN
            sigmoid_f := 2047;
        ELSIF x = 15883 THEN
            sigmoid_f := 2047;
        ELSIF x = 15884 THEN
            sigmoid_f := 2047;
        ELSIF x = 15885 THEN
            sigmoid_f := 2047;
        ELSIF x = 15886 THEN
            sigmoid_f := 2047;
        ELSIF x = 15887 THEN
            sigmoid_f := 2047;
        ELSIF x = 15888 THEN
            sigmoid_f := 2047;
        ELSIF x = 15889 THEN
            sigmoid_f := 2047;
        ELSIF x = 15890 THEN
            sigmoid_f := 2047;
        ELSIF x = 15891 THEN
            sigmoid_f := 2047;
        ELSIF x = 15892 THEN
            sigmoid_f := 2047;
        ELSIF x = 15893 THEN
            sigmoid_f := 2047;
        ELSIF x = 15894 THEN
            sigmoid_f := 2047;
        ELSIF x = 15895 THEN
            sigmoid_f := 2047;
        ELSIF x = 15896 THEN
            sigmoid_f := 2047;
        ELSIF x = 15897 THEN
            sigmoid_f := 2047;
        ELSIF x = 15898 THEN
            sigmoid_f := 2047;
        ELSIF x = 15899 THEN
            sigmoid_f := 2047;
        ELSIF x = 15900 THEN
            sigmoid_f := 2047;
        ELSIF x = 15901 THEN
            sigmoid_f := 2047;
        ELSIF x = 15902 THEN
            sigmoid_f := 2047;
        ELSIF x = 15903 THEN
            sigmoid_f := 2047;
        ELSIF x = 15904 THEN
            sigmoid_f := 2047;
        ELSIF x = 15905 THEN
            sigmoid_f := 2047;
        ELSIF x = 15906 THEN
            sigmoid_f := 2047;
        ELSIF x = 15907 THEN
            sigmoid_f := 2047;
        ELSIF x = 15908 THEN
            sigmoid_f := 2047;
        ELSIF x = 15909 THEN
            sigmoid_f := 2047;
        ELSIF x = 15910 THEN
            sigmoid_f := 2047;
        ELSIF x = 15911 THEN
            sigmoid_f := 2047;
        ELSIF x = 15912 THEN
            sigmoid_f := 2047;
        ELSIF x = 15913 THEN
            sigmoid_f := 2047;
        ELSIF x = 15914 THEN
            sigmoid_f := 2047;
        ELSIF x = 15915 THEN
            sigmoid_f := 2047;
        ELSIF x = 15916 THEN
            sigmoid_f := 2047;
        ELSIF x = 15917 THEN
            sigmoid_f := 2047;
        ELSIF x = 15918 THEN
            sigmoid_f := 2047;
        ELSIF x = 15919 THEN
            sigmoid_f := 2047;
        ELSIF x = 15920 THEN
            sigmoid_f := 2047;
        ELSIF x = 15921 THEN
            sigmoid_f := 2047;
        ELSIF x = 15922 THEN
            sigmoid_f := 2047;
        ELSIF x = 15923 THEN
            sigmoid_f := 2047;
        ELSIF x = 15924 THEN
            sigmoid_f := 2047;
        ELSIF x = 15925 THEN
            sigmoid_f := 2047;
        ELSIF x = 15926 THEN
            sigmoid_f := 2047;
        ELSIF x = 15927 THEN
            sigmoid_f := 2047;
        ELSIF x = 15928 THEN
            sigmoid_f := 2047;
        ELSIF x = 15929 THEN
            sigmoid_f := 2047;
        ELSIF x = 15930 THEN
            sigmoid_f := 2047;
        ELSIF x = 15931 THEN
            sigmoid_f := 2047;
        ELSIF x = 15932 THEN
            sigmoid_f := 2047;
        ELSIF x = 15933 THEN
            sigmoid_f := 2047;
        ELSIF x = 15934 THEN
            sigmoid_f := 2047;
        ELSIF x = 15935 THEN
            sigmoid_f := 2047;
        ELSIF x = 15936 THEN
            sigmoid_f := 2047;
        ELSIF x = 15937 THEN
            sigmoid_f := 2047;
        ELSIF x = 15938 THEN
            sigmoid_f := 2047;
        ELSIF x = 15939 THEN
            sigmoid_f := 2047;
        ELSIF x = 15940 THEN
            sigmoid_f := 2047;
        ELSIF x = 15941 THEN
            sigmoid_f := 2047;
        ELSIF x = 15942 THEN
            sigmoid_f := 2047;
        ELSIF x = 15943 THEN
            sigmoid_f := 2047;
        ELSIF x = 15944 THEN
            sigmoid_f := 2047;
        ELSIF x = 15945 THEN
            sigmoid_f := 2047;
        ELSIF x = 15946 THEN
            sigmoid_f := 2047;
        ELSIF x = 15947 THEN
            sigmoid_f := 2047;
        ELSIF x = 15948 THEN
            sigmoid_f := 2047;
        ELSIF x = 15949 THEN
            sigmoid_f := 2047;
        ELSIF x = 15950 THEN
            sigmoid_f := 2047;
        ELSIF x = 15951 THEN
            sigmoid_f := 2047;
        ELSIF x = 15952 THEN
            sigmoid_f := 2047;
        ELSIF x = 15953 THEN
            sigmoid_f := 2047;
        ELSIF x = 15954 THEN
            sigmoid_f := 2047;
        ELSIF x = 15955 THEN
            sigmoid_f := 2047;
        ELSIF x = 15956 THEN
            sigmoid_f := 2047;
        ELSIF x = 15957 THEN
            sigmoid_f := 2047;
        ELSIF x = 15958 THEN
            sigmoid_f := 2047;
        ELSIF x = 15959 THEN
            sigmoid_f := 2047;
        ELSIF x = 15960 THEN
            sigmoid_f := 2047;
        ELSIF x = 15961 THEN
            sigmoid_f := 2047;
        ELSIF x = 15962 THEN
            sigmoid_f := 2047;
        ELSIF x = 15963 THEN
            sigmoid_f := 2047;
        ELSIF x = 15964 THEN
            sigmoid_f := 2047;
        ELSIF x = 15965 THEN
            sigmoid_f := 2047;
        ELSIF x = 15966 THEN
            sigmoid_f := 2047;
        ELSIF x = 15967 THEN
            sigmoid_f := 2047;
        ELSIF x = 15968 THEN
            sigmoid_f := 2047;
        ELSIF x = 15969 THEN
            sigmoid_f := 2047;
        ELSIF x = 15970 THEN
            sigmoid_f := 2047;
        ELSIF x = 15971 THEN
            sigmoid_f := 2047;
        ELSIF x = 15972 THEN
            sigmoid_f := 2047;
        ELSIF x = 15973 THEN
            sigmoid_f := 2047;
        ELSIF x = 15974 THEN
            sigmoid_f := 2047;
        ELSIF x = 15975 THEN
            sigmoid_f := 2047;
        ELSIF x = 15976 THEN
            sigmoid_f := 2047;
        ELSIF x = 15977 THEN
            sigmoid_f := 2047;
        ELSIF x = 15978 THEN
            sigmoid_f := 2047;
        ELSIF x = 15979 THEN
            sigmoid_f := 2047;
        ELSIF x = 15980 THEN
            sigmoid_f := 2047;
        ELSIF x = 15981 THEN
            sigmoid_f := 2047;
        ELSIF x = 15982 THEN
            sigmoid_f := 2047;
        ELSIF x = 15983 THEN
            sigmoid_f := 2047;
        ELSIF x = 15984 THEN
            sigmoid_f := 2047;
        ELSIF x = 15985 THEN
            sigmoid_f := 2047;
        ELSIF x = 15986 THEN
            sigmoid_f := 2047;
        ELSIF x = 15987 THEN
            sigmoid_f := 2047;
        ELSIF x = 15988 THEN
            sigmoid_f := 2047;
        ELSIF x = 15989 THEN
            sigmoid_f := 2047;
        ELSIF x = 15990 THEN
            sigmoid_f := 2047;
        ELSIF x = 15991 THEN
            sigmoid_f := 2047;
        ELSIF x = 15992 THEN
            sigmoid_f := 2047;
        ELSIF x = 15993 THEN
            sigmoid_f := 2047;
        ELSIF x = 15994 THEN
            sigmoid_f := 2047;
        ELSIF x = 15995 THEN
            sigmoid_f := 2047;
        ELSIF x = 15996 THEN
            sigmoid_f := 2047;
        ELSIF x = 15997 THEN
            sigmoid_f := 2047;
        ELSIF x = 15998 THEN
            sigmoid_f := 2047;
        ELSIF x = 15999 THEN
            sigmoid_f := 2047;
        ELSIF x = 16000 THEN
            sigmoid_f := 2047;
        ELSIF x = 16001 THEN
            sigmoid_f := 2047;
        ELSIF x = 16002 THEN
            sigmoid_f := 2047;
        ELSIF x = 16003 THEN
            sigmoid_f := 2047;
        ELSIF x = 16004 THEN
            sigmoid_f := 2047;
        ELSIF x = 16005 THEN
            sigmoid_f := 2047;
        ELSIF x = 16006 THEN
            sigmoid_f := 2047;
        ELSIF x = 16007 THEN
            sigmoid_f := 2047;
        ELSIF x = 16008 THEN
            sigmoid_f := 2047;
        ELSIF x = 16009 THEN
            sigmoid_f := 2047;
        ELSIF x = 16010 THEN
            sigmoid_f := 2047;
        ELSIF x = 16011 THEN
            sigmoid_f := 2047;
        ELSIF x = 16012 THEN
            sigmoid_f := 2047;
        ELSIF x = 16013 THEN
            sigmoid_f := 2047;
        ELSIF x = 16014 THEN
            sigmoid_f := 2047;
        ELSIF x = 16015 THEN
            sigmoid_f := 2047;
        ELSIF x = 16016 THEN
            sigmoid_f := 2047;
        ELSIF x = 16017 THEN
            sigmoid_f := 2047;
        ELSIF x = 16018 THEN
            sigmoid_f := 2047;
        ELSIF x = 16019 THEN
            sigmoid_f := 2047;
        ELSIF x = 16020 THEN
            sigmoid_f := 2047;
        ELSIF x = 16021 THEN
            sigmoid_f := 2047;
        ELSIF x = 16022 THEN
            sigmoid_f := 2047;
        ELSIF x = 16023 THEN
            sigmoid_f := 2047;
        ELSIF x = 16024 THEN
            sigmoid_f := 2047;
        ELSIF x = 16025 THEN
            sigmoid_f := 2047;
        ELSIF x = 16026 THEN
            sigmoid_f := 2047;
        ELSIF x = 16027 THEN
            sigmoid_f := 2047;
        ELSIF x = 16028 THEN
            sigmoid_f := 2047;
        ELSIF x = 16029 THEN
            sigmoid_f := 2047;
        ELSIF x = 16030 THEN
            sigmoid_f := 2047;
        ELSIF x = 16031 THEN
            sigmoid_f := 2047;
        ELSIF x = 16032 THEN
            sigmoid_f := 2047;
        ELSIF x = 16033 THEN
            sigmoid_f := 2047;
        ELSIF x = 16034 THEN
            sigmoid_f := 2047;
        ELSIF x = 16035 THEN
            sigmoid_f := 2047;
        ELSIF x = 16036 THEN
            sigmoid_f := 2047;
        ELSIF x = 16037 THEN
            sigmoid_f := 2047;
        ELSIF x = 16038 THEN
            sigmoid_f := 2047;
        ELSIF x = 16039 THEN
            sigmoid_f := 2047;
        ELSIF x = 16040 THEN
            sigmoid_f := 2047;
        ELSIF x = 16041 THEN
            sigmoid_f := 2047;
        ELSIF x = 16042 THEN
            sigmoid_f := 2047;
        ELSIF x = 16043 THEN
            sigmoid_f := 2047;
        ELSIF x = 16044 THEN
            sigmoid_f := 2047;
        ELSIF x = 16045 THEN
            sigmoid_f := 2047;
        ELSIF x = 16046 THEN
            sigmoid_f := 2047;
        ELSIF x = 16047 THEN
            sigmoid_f := 2047;
        ELSIF x = 16048 THEN
            sigmoid_f := 2047;
        ELSIF x = 16049 THEN
            sigmoid_f := 2047;
        ELSIF x = 16050 THEN
            sigmoid_f := 2047;
        ELSIF x = 16051 THEN
            sigmoid_f := 2047;
        ELSIF x = 16052 THEN
            sigmoid_f := 2047;
        ELSIF x = 16053 THEN
            sigmoid_f := 2047;
        ELSIF x = 16054 THEN
            sigmoid_f := 2047;
        ELSIF x = 16055 THEN
            sigmoid_f := 2047;
        ELSIF x = 16056 THEN
            sigmoid_f := 2047;
        ELSIF x = 16057 THEN
            sigmoid_f := 2047;
        ELSIF x = 16058 THEN
            sigmoid_f := 2047;
        ELSIF x = 16059 THEN
            sigmoid_f := 2047;
        ELSIF x = 16060 THEN
            sigmoid_f := 2047;
        ELSIF x = 16061 THEN
            sigmoid_f := 2047;
        ELSIF x = 16062 THEN
            sigmoid_f := 2047;
        ELSIF x = 16063 THEN
            sigmoid_f := 2047;
        ELSIF x = 16064 THEN
            sigmoid_f := 2047;
        ELSIF x = 16065 THEN
            sigmoid_f := 2047;
        ELSIF x = 16066 THEN
            sigmoid_f := 2047;
        ELSIF x = 16067 THEN
            sigmoid_f := 2047;
        ELSIF x = 16068 THEN
            sigmoid_f := 2047;
        ELSIF x = 16069 THEN
            sigmoid_f := 2047;
        ELSIF x = 16070 THEN
            sigmoid_f := 2047;
        ELSIF x = 16071 THEN
            sigmoid_f := 2047;
        ELSIF x = 16072 THEN
            sigmoid_f := 2047;
        ELSIF x = 16073 THEN
            sigmoid_f := 2047;
        ELSIF x = 16074 THEN
            sigmoid_f := 2047;
        ELSIF x = 16075 THEN
            sigmoid_f := 2047;
        ELSIF x = 16076 THEN
            sigmoid_f := 2047;
        ELSIF x = 16077 THEN
            sigmoid_f := 2047;
        ELSIF x = 16078 THEN
            sigmoid_f := 2047;
        ELSIF x = 16079 THEN
            sigmoid_f := 2047;
        ELSIF x = 16080 THEN
            sigmoid_f := 2047;
        ELSIF x = 16081 THEN
            sigmoid_f := 2047;
        ELSIF x = 16082 THEN
            sigmoid_f := 2047;
        ELSIF x = 16083 THEN
            sigmoid_f := 2047;
        ELSIF x = 16084 THEN
            sigmoid_f := 2047;
        ELSIF x = 16085 THEN
            sigmoid_f := 2047;
        ELSIF x = 16086 THEN
            sigmoid_f := 2047;
        ELSIF x = 16087 THEN
            sigmoid_f := 2047;
        ELSIF x = 16088 THEN
            sigmoid_f := 2047;
        ELSIF x = 16089 THEN
            sigmoid_f := 2047;
        ELSIF x = 16090 THEN
            sigmoid_f := 2047;
        ELSIF x = 16091 THEN
            sigmoid_f := 2047;
        ELSIF x = 16092 THEN
            sigmoid_f := 2047;
        ELSIF x = 16093 THEN
            sigmoid_f := 2047;
        ELSIF x = 16094 THEN
            sigmoid_f := 2047;
        ELSIF x = 16095 THEN
            sigmoid_f := 2047;
        ELSIF x = 16096 THEN
            sigmoid_f := 2047;
        ELSIF x = 16097 THEN
            sigmoid_f := 2047;
        ELSIF x = 16098 THEN
            sigmoid_f := 2047;
        ELSIF x = 16099 THEN
            sigmoid_f := 2047;
        ELSIF x = 16100 THEN
            sigmoid_f := 2047;
        ELSIF x = 16101 THEN
            sigmoid_f := 2047;
        ELSIF x = 16102 THEN
            sigmoid_f := 2047;
        ELSIF x = 16103 THEN
            sigmoid_f := 2047;
        ELSIF x = 16104 THEN
            sigmoid_f := 2047;
        ELSIF x = 16105 THEN
            sigmoid_f := 2047;
        ELSIF x = 16106 THEN
            sigmoid_f := 2047;
        ELSIF x = 16107 THEN
            sigmoid_f := 2047;
        ELSIF x = 16108 THEN
            sigmoid_f := 2047;
        ELSIF x = 16109 THEN
            sigmoid_f := 2047;
        ELSIF x = 16110 THEN
            sigmoid_f := 2047;
        ELSIF x = 16111 THEN
            sigmoid_f := 2047;
        ELSIF x = 16112 THEN
            sigmoid_f := 2047;
        ELSIF x = 16113 THEN
            sigmoid_f := 2047;
        ELSIF x = 16114 THEN
            sigmoid_f := 2047;
        ELSIF x = 16115 THEN
            sigmoid_f := 2047;
        ELSIF x = 16116 THEN
            sigmoid_f := 2047;
        ELSIF x = 16117 THEN
            sigmoid_f := 2047;
        ELSIF x = 16118 THEN
            sigmoid_f := 2047;
        ELSIF x = 16119 THEN
            sigmoid_f := 2047;
        ELSIF x = 16120 THEN
            sigmoid_f := 2047;
        ELSIF x = 16121 THEN
            sigmoid_f := 2047;
        ELSIF x = 16122 THEN
            sigmoid_f := 2047;
        ELSIF x = 16123 THEN
            sigmoid_f := 2047;
        ELSIF x = 16124 THEN
            sigmoid_f := 2047;
        ELSIF x = 16125 THEN
            sigmoid_f := 2047;
        ELSIF x = 16126 THEN
            sigmoid_f := 2047;
        ELSIF x = 16127 THEN
            sigmoid_f := 2047;
        ELSIF x = 16128 THEN
            sigmoid_f := 2047;
        ELSIF x = 16129 THEN
            sigmoid_f := 2047;
        ELSIF x = 16130 THEN
            sigmoid_f := 2047;
        ELSIF x = 16131 THEN
            sigmoid_f := 2047;
        ELSIF x = 16132 THEN
            sigmoid_f := 2047;
        ELSIF x = 16133 THEN
            sigmoid_f := 2047;
        ELSIF x = 16134 THEN
            sigmoid_f := 2047;
        ELSIF x = 16135 THEN
            sigmoid_f := 2047;
        ELSIF x = 16136 THEN
            sigmoid_f := 2047;
        ELSIF x = 16137 THEN
            sigmoid_f := 2047;
        ELSIF x = 16138 THEN
            sigmoid_f := 2047;
        ELSIF x = 16139 THEN
            sigmoid_f := 2047;
        ELSIF x = 16140 THEN
            sigmoid_f := 2047;
        ELSIF x = 16141 THEN
            sigmoid_f := 2047;
        ELSIF x = 16142 THEN
            sigmoid_f := 2047;
        ELSIF x = 16143 THEN
            sigmoid_f := 2047;
        ELSIF x = 16144 THEN
            sigmoid_f := 2047;
        ELSIF x = 16145 THEN
            sigmoid_f := 2047;
        ELSIF x = 16146 THEN
            sigmoid_f := 2047;
        ELSIF x = 16147 THEN
            sigmoid_f := 2047;
        ELSIF x = 16148 THEN
            sigmoid_f := 2047;
        ELSIF x = 16149 THEN
            sigmoid_f := 2047;
        ELSIF x = 16150 THEN
            sigmoid_f := 2047;
        ELSIF x = 16151 THEN
            sigmoid_f := 2047;
        ELSIF x = 16152 THEN
            sigmoid_f := 2047;
        ELSIF x = 16153 THEN
            sigmoid_f := 2047;
        ELSIF x = 16154 THEN
            sigmoid_f := 2047;
        ELSIF x = 16155 THEN
            sigmoid_f := 2047;
        ELSIF x = 16156 THEN
            sigmoid_f := 2047;
        ELSIF x = 16157 THEN
            sigmoid_f := 2047;
        ELSIF x = 16158 THEN
            sigmoid_f := 2047;
        ELSIF x = 16159 THEN
            sigmoid_f := 2047;
        ELSIF x = 16160 THEN
            sigmoid_f := 2047;
        ELSIF x = 16161 THEN
            sigmoid_f := 2047;
        ELSIF x = 16162 THEN
            sigmoid_f := 2047;
        ELSIF x = 16163 THEN
            sigmoid_f := 2047;
        ELSIF x = 16164 THEN
            sigmoid_f := 2047;
        ELSIF x = 16165 THEN
            sigmoid_f := 2047;
        ELSIF x = 16166 THEN
            sigmoid_f := 2047;
        ELSIF x = 16167 THEN
            sigmoid_f := 2047;
        ELSIF x = 16168 THEN
            sigmoid_f := 2047;
        ELSIF x = 16169 THEN
            sigmoid_f := 2047;
        ELSIF x = 16170 THEN
            sigmoid_f := 2047;
        ELSIF x = 16171 THEN
            sigmoid_f := 2047;
        ELSIF x = 16172 THEN
            sigmoid_f := 2047;
        ELSIF x = 16173 THEN
            sigmoid_f := 2047;
        ELSIF x = 16174 THEN
            sigmoid_f := 2047;
        ELSIF x = 16175 THEN
            sigmoid_f := 2047;
        ELSIF x = 16176 THEN
            sigmoid_f := 2047;
        ELSIF x = 16177 THEN
            sigmoid_f := 2047;
        ELSIF x = 16178 THEN
            sigmoid_f := 2047;
        ELSIF x = 16179 THEN
            sigmoid_f := 2047;
        ELSIF x = 16180 THEN
            sigmoid_f := 2047;
        ELSIF x = 16181 THEN
            sigmoid_f := 2047;
        ELSIF x = 16182 THEN
            sigmoid_f := 2047;
        ELSIF x = 16183 THEN
            sigmoid_f := 2047;
        ELSIF x = 16184 THEN
            sigmoid_f := 2047;
        ELSIF x = 16185 THEN
            sigmoid_f := 2047;
        ELSIF x = 16186 THEN
            sigmoid_f := 2047;
        ELSIF x = 16187 THEN
            sigmoid_f := 2047;
        ELSIF x = 16188 THEN
            sigmoid_f := 2047;
        ELSIF x = 16189 THEN
            sigmoid_f := 2047;
        ELSIF x = 16190 THEN
            sigmoid_f := 2047;
        ELSIF x = 16191 THEN
            sigmoid_f := 2047;
        ELSIF x = 16192 THEN
            sigmoid_f := 2047;
        ELSIF x = 16193 THEN
            sigmoid_f := 2047;
        ELSIF x = 16194 THEN
            sigmoid_f := 2047;
        ELSIF x = 16195 THEN
            sigmoid_f := 2047;
        ELSIF x = 16196 THEN
            sigmoid_f := 2047;
        ELSIF x = 16197 THEN
            sigmoid_f := 2047;
        ELSIF x = 16198 THEN
            sigmoid_f := 2047;
        ELSIF x = 16199 THEN
            sigmoid_f := 2047;
        ELSIF x = 16200 THEN
            sigmoid_f := 2047;
        ELSIF x = 16201 THEN
            sigmoid_f := 2047;
        ELSIF x = 16202 THEN
            sigmoid_f := 2047;
        ELSIF x = 16203 THEN
            sigmoid_f := 2047;
        ELSIF x = 16204 THEN
            sigmoid_f := 2047;
        ELSIF x = 16205 THEN
            sigmoid_f := 2047;
        ELSIF x = 16206 THEN
            sigmoid_f := 2047;
        ELSIF x = 16207 THEN
            sigmoid_f := 2047;
        ELSIF x = 16208 THEN
            sigmoid_f := 2047;
        ELSIF x = 16209 THEN
            sigmoid_f := 2047;
        ELSIF x = 16210 THEN
            sigmoid_f := 2047;
        ELSIF x = 16211 THEN
            sigmoid_f := 2047;
        ELSIF x = 16212 THEN
            sigmoid_f := 2047;
        ELSIF x = 16213 THEN
            sigmoid_f := 2047;
        ELSIF x = 16214 THEN
            sigmoid_f := 2047;
        ELSIF x = 16215 THEN
            sigmoid_f := 2047;
        ELSIF x = 16216 THEN
            sigmoid_f := 2047;
        ELSIF x = 16217 THEN
            sigmoid_f := 2047;
        ELSIF x = 16218 THEN
            sigmoid_f := 2047;
        ELSIF x = 16219 THEN
            sigmoid_f := 2047;
        ELSIF x = 16220 THEN
            sigmoid_f := 2047;
        ELSIF x = 16221 THEN
            sigmoid_f := 2047;
        ELSIF x = 16222 THEN
            sigmoid_f := 2047;
        ELSIF x = 16223 THEN
            sigmoid_f := 2047;
        ELSIF x = 16224 THEN
            sigmoid_f := 2047;
        ELSIF x = 16225 THEN
            sigmoid_f := 2047;
        ELSIF x = 16226 THEN
            sigmoid_f := 2047;
        ELSIF x = 16227 THEN
            sigmoid_f := 2047;
        ELSIF x = 16228 THEN
            sigmoid_f := 2047;
        ELSIF x = 16229 THEN
            sigmoid_f := 2047;
        ELSIF x = 16230 THEN
            sigmoid_f := 2047;
        ELSIF x = 16231 THEN
            sigmoid_f := 2047;
        ELSIF x = 16232 THEN
            sigmoid_f := 2047;
        ELSIF x = 16233 THEN
            sigmoid_f := 2047;
        ELSIF x = 16234 THEN
            sigmoid_f := 2047;
        ELSIF x = 16235 THEN
            sigmoid_f := 2047;
        ELSIF x = 16236 THEN
            sigmoid_f := 2047;
        ELSIF x = 16237 THEN
            sigmoid_f := 2047;
        ELSIF x = 16238 THEN
            sigmoid_f := 2047;
        ELSIF x = 16239 THEN
            sigmoid_f := 2047;
        ELSIF x = 16240 THEN
            sigmoid_f := 2047;
        ELSIF x = 16241 THEN
            sigmoid_f := 2047;
        ELSIF x = 16242 THEN
            sigmoid_f := 2047;
        ELSIF x = 16243 THEN
            sigmoid_f := 2047;
        ELSIF x = 16244 THEN
            sigmoid_f := 2047;
        ELSIF x = 16245 THEN
            sigmoid_f := 2047;
        ELSIF x = 16246 THEN
            sigmoid_f := 2047;
        ELSIF x = 16247 THEN
            sigmoid_f := 2047;
        ELSIF x = 16248 THEN
            sigmoid_f := 2047;
        ELSIF x = 16249 THEN
            sigmoid_f := 2047;
        ELSIF x = 16250 THEN
            sigmoid_f := 2047;
        ELSIF x = 16251 THEN
            sigmoid_f := 2047;
        ELSIF x = 16252 THEN
            sigmoid_f := 2047;
        ELSIF x = 16253 THEN
            sigmoid_f := 2047;
        ELSIF x = 16254 THEN
            sigmoid_f := 2047;
        ELSIF x = 16255 THEN
            sigmoid_f := 2047;
        ELSIF x = 16256 THEN
            sigmoid_f := 2047;
        ELSIF x = 16257 THEN
            sigmoid_f := 2047;
        ELSIF x = 16258 THEN
            sigmoid_f := 2047;
        ELSIF x = 16259 THEN
            sigmoid_f := 2047;
        ELSIF x = 16260 THEN
            sigmoid_f := 2047;
        ELSIF x = 16261 THEN
            sigmoid_f := 2047;
        ELSIF x = 16262 THEN
            sigmoid_f := 2047;
        ELSIF x = 16263 THEN
            sigmoid_f := 2047;
        ELSIF x = 16264 THEN
            sigmoid_f := 2047;
        ELSIF x = 16265 THEN
            sigmoid_f := 2047;
        ELSIF x = 16266 THEN
            sigmoid_f := 2047;
        ELSIF x = 16267 THEN
            sigmoid_f := 2047;
        ELSIF x = 16268 THEN
            sigmoid_f := 2047;
        ELSIF x = 16269 THEN
            sigmoid_f := 2047;
        ELSIF x = 16270 THEN
            sigmoid_f := 2047;
        ELSIF x = 16271 THEN
            sigmoid_f := 2047;
        ELSIF x = 16272 THEN
            sigmoid_f := 2047;
        ELSIF x = 16273 THEN
            sigmoid_f := 2047;
        ELSIF x = 16274 THEN
            sigmoid_f := 2047;
        ELSIF x = 16275 THEN
            sigmoid_f := 2047;
        ELSIF x = 16276 THEN
            sigmoid_f := 2047;
        ELSIF x = 16277 THEN
            sigmoid_f := 2047;
        ELSIF x = 16278 THEN
            sigmoid_f := 2047;
        ELSIF x = 16279 THEN
            sigmoid_f := 2047;
        ELSIF x = 16280 THEN
            sigmoid_f := 2047;
        ELSIF x = 16281 THEN
            sigmoid_f := 2047;
        ELSIF x = 16282 THEN
            sigmoid_f := 2047;
        ELSIF x = 16283 THEN
            sigmoid_f := 2047;
        ELSIF x = 16284 THEN
            sigmoid_f := 2047;
        ELSIF x = 16285 THEN
            sigmoid_f := 2047;
        ELSIF x = 16286 THEN
            sigmoid_f := 2047;
        ELSIF x = 16287 THEN
            sigmoid_f := 2047;
        ELSIF x = 16288 THEN
            sigmoid_f := 2047;
        ELSIF x = 16289 THEN
            sigmoid_f := 2047;
        ELSIF x = 16290 THEN
            sigmoid_f := 2047;
        ELSIF x = 16291 THEN
            sigmoid_f := 2047;
        ELSIF x = 16292 THEN
            sigmoid_f := 2047;
        ELSIF x = 16293 THEN
            sigmoid_f := 2047;
        ELSIF x = 16294 THEN
            sigmoid_f := 2047;
        ELSIF x = 16295 THEN
            sigmoid_f := 2047;
        ELSIF x = 16296 THEN
            sigmoid_f := 2047;
        ELSIF x = 16297 THEN
            sigmoid_f := 2047;
        ELSIF x = 16298 THEN
            sigmoid_f := 2047;
        ELSIF x = 16299 THEN
            sigmoid_f := 2047;
        ELSIF x = 16300 THEN
            sigmoid_f := 2047;
        ELSIF x = 16301 THEN
            sigmoid_f := 2047;
        ELSIF x = 16302 THEN
            sigmoid_f := 2047;
        ELSIF x = 16303 THEN
            sigmoid_f := 2047;
        ELSIF x = 16304 THEN
            sigmoid_f := 2047;
        ELSIF x = 16305 THEN
            sigmoid_f := 2047;
        ELSIF x = 16306 THEN
            sigmoid_f := 2047;
        ELSIF x = 16307 THEN
            sigmoid_f := 2047;
        ELSIF x = 16308 THEN
            sigmoid_f := 2047;
        ELSIF x = 16309 THEN
            sigmoid_f := 2047;
        ELSIF x = 16310 THEN
            sigmoid_f := 2047;
        ELSIF x = 16311 THEN
            sigmoid_f := 2047;
        ELSIF x = 16312 THEN
            sigmoid_f := 2047;
        ELSIF x = 16313 THEN
            sigmoid_f := 2047;
        ELSIF x = 16314 THEN
            sigmoid_f := 2047;
        ELSIF x = 16315 THEN
            sigmoid_f := 2047;
        ELSIF x = 16316 THEN
            sigmoid_f := 2047;
        ELSIF x = 16317 THEN
            sigmoid_f := 2047;
        ELSIF x = 16318 THEN
            sigmoid_f := 2047;
        ELSIF x = 16319 THEN
            sigmoid_f := 2047;
        ELSIF x = 16320 THEN
            sigmoid_f := 2047;
        ELSIF x = 16321 THEN
            sigmoid_f := 2047;
        ELSIF x = 16322 THEN
            sigmoid_f := 2047;
        ELSIF x = 16323 THEN
            sigmoid_f := 2047;
        ELSIF x = 16324 THEN
            sigmoid_f := 2047;
        ELSIF x = 16325 THEN
            sigmoid_f := 2047;
        ELSIF x = 16326 THEN
            sigmoid_f := 2047;
        ELSIF x = 16327 THEN
            sigmoid_f := 2047;
        ELSIF x = 16328 THEN
            sigmoid_f := 2047;
        ELSIF x = 16329 THEN
            sigmoid_f := 2047;
        ELSIF x = 16330 THEN
            sigmoid_f := 2047;
        ELSIF x = 16331 THEN
            sigmoid_f := 2047;
        ELSIF x = 16332 THEN
            sigmoid_f := 2047;
        ELSIF x = 16333 THEN
            sigmoid_f := 2047;
        ELSIF x = 16334 THEN
            sigmoid_f := 2047;
        ELSIF x = 16335 THEN
            sigmoid_f := 2047;
        ELSIF x = 16336 THEN
            sigmoid_f := 2047;
        ELSIF x = 16337 THEN
            sigmoid_f := 2047;
        ELSIF x = 16338 THEN
            sigmoid_f := 2047;
        ELSIF x = 16339 THEN
            sigmoid_f := 2047;
        ELSIF x = 16340 THEN
            sigmoid_f := 2047;
        ELSIF x = 16341 THEN
            sigmoid_f := 2047;
        ELSIF x = 16342 THEN
            sigmoid_f := 2047;
        ELSIF x = 16343 THEN
            sigmoid_f := 2047;
        ELSIF x = 16344 THEN
            sigmoid_f := 2047;
        ELSIF x = 16345 THEN
            sigmoid_f := 2047;
        ELSIF x = 16346 THEN
            sigmoid_f := 2047;
        ELSIF x = 16347 THEN
            sigmoid_f := 2047;
        ELSIF x = 16348 THEN
            sigmoid_f := 2047;
        ELSIF x = 16349 THEN
            sigmoid_f := 2047;
        ELSIF x = 16350 THEN
            sigmoid_f := 2047;
        ELSIF x = 16351 THEN
            sigmoid_f := 2047;
        ELSIF x = 16352 THEN
            sigmoid_f := 2047;
        ELSIF x = 16353 THEN
            sigmoid_f := 2047;
        ELSIF x = 16354 THEN
            sigmoid_f := 2047;
        ELSIF x = 16355 THEN
            sigmoid_f := 2047;
        ELSIF x = 16356 THEN
            sigmoid_f := 2047;
        ELSIF x = 16357 THEN
            sigmoid_f := 2047;
        ELSIF x = 16358 THEN
            sigmoid_f := 2047;
        ELSIF x = 16359 THEN
            sigmoid_f := 2047;
        ELSIF x = 16360 THEN
            sigmoid_f := 2047;
        ELSIF x = 16361 THEN
            sigmoid_f := 2047;
        ELSIF x = 16362 THEN
            sigmoid_f := 2047;
        ELSIF x = 16363 THEN
            sigmoid_f := 2047;
        ELSIF x = 16364 THEN
            sigmoid_f := 2047;
        ELSIF x = 16365 THEN
            sigmoid_f := 2047;
        ELSIF x = 16366 THEN
            sigmoid_f := 2047;
        ELSIF x = 16367 THEN
            sigmoid_f := 2047;
        ELSIF x = 16368 THEN
            sigmoid_f := 2047;
        ELSIF x = 16369 THEN
            sigmoid_f := 2047;
        ELSIF x = 16370 THEN
            sigmoid_f := 2047;
        ELSIF x = 16371 THEN
            sigmoid_f := 2047;
        ELSIF x = 16372 THEN
            sigmoid_f := 2047;
        ELSIF x = 16373 THEN
            sigmoid_f := 2047;
        ELSIF x = 16374 THEN
            sigmoid_f := 2047;
        ELSIF x = 16375 THEN
            sigmoid_f := 2047;
        ELSIF x = 16376 THEN
            sigmoid_f := 2047;
        ELSIF x = 16377 THEN
            sigmoid_f := 2047;
        ELSIF x = 16378 THEN
            sigmoid_f := 2047;
        ELSIF x = 16379 THEN
            sigmoid_f := 2047;
        ELSIF x = 16380 THEN
            sigmoid_f := 2047;
        ELSIF x = 16381 THEN
            sigmoid_f := 2047;
        ELSIF x = 16382 THEN
            sigmoid_f := 2047;
        ELSIF x = 16383 THEN
            sigmoid_f := 2047;
        ELSIF x = 16384 THEN
            sigmoid_f := 2047;
        ELSIF x = 16385 THEN
            sigmoid_f := 2047;
        ELSIF x = 16386 THEN
            sigmoid_f := 2047;
        ELSIF x = 16387 THEN
            sigmoid_f := 2047;
        ELSIF x = 16388 THEN
            sigmoid_f := 2047;
        ELSIF x = 16389 THEN
            sigmoid_f := 2047;
        ELSIF x = 16390 THEN
            sigmoid_f := 2047;
        ELSIF x = 16391 THEN
            sigmoid_f := 2047;
        ELSIF x = 16392 THEN
            sigmoid_f := 2047;
        ELSIF x = 16393 THEN
            sigmoid_f := 2047;
        ELSIF x = 16394 THEN
            sigmoid_f := 2047;
        ELSIF x = 16395 THEN
            sigmoid_f := 2047;
        ELSIF x = 16396 THEN
            sigmoid_f := 2047;
        ELSIF x = 16397 THEN
            sigmoid_f := 2047;
        ELSIF x = 16398 THEN
            sigmoid_f := 2047;
        ELSIF x = 16399 THEN
            sigmoid_f := 2047;
        ELSIF x = 16400 THEN
            sigmoid_f := 2047;
        ELSIF x = 16401 THEN
            sigmoid_f := 2047;
        ELSIF x = 16402 THEN
            sigmoid_f := 2047;
        ELSIF x = 16403 THEN
            sigmoid_f := 2047;
        ELSIF x = 16404 THEN
            sigmoid_f := 2047;
        ELSIF x = 16405 THEN
            sigmoid_f := 2047;
        ELSIF x = 16406 THEN
            sigmoid_f := 2047;
        ELSIF x = 16407 THEN
            sigmoid_f := 2047;
        ELSIF x = 16408 THEN
            sigmoid_f := 2047;
        ELSIF x = 16409 THEN
            sigmoid_f := 2047;
        ELSIF x = 16410 THEN
            sigmoid_f := 2047;
        ELSIF x = 16411 THEN
            sigmoid_f := 2047;
        ELSIF x = 16412 THEN
            sigmoid_f := 2047;
        ELSIF x = 16413 THEN
            sigmoid_f := 2047;
        ELSIF x = 16414 THEN
            sigmoid_f := 2047;
        ELSIF x = 16415 THEN
            sigmoid_f := 2047;
        ELSIF x = 16416 THEN
            sigmoid_f := 2047;
        ELSIF x = 16417 THEN
            sigmoid_f := 2047;
        ELSIF x = 16418 THEN
            sigmoid_f := 2047;
        ELSIF x = 16419 THEN
            sigmoid_f := 2047;
        ELSIF x = 16420 THEN
            sigmoid_f := 2047;
        ELSIF x = 16421 THEN
            sigmoid_f := 2047;
        ELSIF x = 16422 THEN
            sigmoid_f := 2047;
        ELSIF x = 16423 THEN
            sigmoid_f := 2047;
        ELSIF x = 16424 THEN
            sigmoid_f := 2047;
        ELSIF x = 16425 THEN
            sigmoid_f := 2047;
        ELSIF x = 16426 THEN
            sigmoid_f := 2047;
        ELSIF x = 16427 THEN
            sigmoid_f := 2047;
        ELSIF x = 16428 THEN
            sigmoid_f := 2047;
        ELSIF x = 16429 THEN
            sigmoid_f := 2047;
        ELSIF x = 16430 THEN
            sigmoid_f := 2047;
        ELSIF x = 16431 THEN
            sigmoid_f := 2047;
        ELSIF x = 16432 THEN
            sigmoid_f := 2047;
        ELSIF x = 16433 THEN
            sigmoid_f := 2047;
        ELSIF x = 16434 THEN
            sigmoid_f := 2047;
        ELSIF x = 16435 THEN
            sigmoid_f := 2047;
        ELSIF x = 16436 THEN
            sigmoid_f := 2047;
        ELSIF x = 16437 THEN
            sigmoid_f := 2047;
        ELSIF x = 16438 THEN
            sigmoid_f := 2047;
        ELSIF x = 16439 THEN
            sigmoid_f := 2047;
        ELSIF x = 16440 THEN
            sigmoid_f := 2047;
        ELSIF x = 16441 THEN
            sigmoid_f := 2047;
        ELSIF x = 16442 THEN
            sigmoid_f := 2047;
        ELSIF x = 16443 THEN
            sigmoid_f := 2047;
        ELSIF x = 16444 THEN
            sigmoid_f := 2047;
        ELSIF x = 16445 THEN
            sigmoid_f := 2047;
        ELSIF x = 16446 THEN
            sigmoid_f := 2047;
        ELSIF x = 16447 THEN
            sigmoid_f := 2047;
        ELSIF x = 16448 THEN
            sigmoid_f := 2047;
        ELSIF x = 16449 THEN
            sigmoid_f := 2047;
        ELSIF x = 16450 THEN
            sigmoid_f := 2047;
        ELSIF x = 16451 THEN
            sigmoid_f := 2047;
        ELSIF x = 16452 THEN
            sigmoid_f := 2047;
        ELSIF x = 16453 THEN
            sigmoid_f := 2047;
        ELSIF x = 16454 THEN
            sigmoid_f := 2047;
        ELSIF x = 16455 THEN
            sigmoid_f := 2047;
        ELSIF x = 16456 THEN
            sigmoid_f := 2047;
        ELSIF x = 16457 THEN
            sigmoid_f := 2047;
        ELSIF x = 16458 THEN
            sigmoid_f := 2047;
        ELSIF x = 16459 THEN
            sigmoid_f := 2047;
        ELSIF x = 16460 THEN
            sigmoid_f := 2047;
        ELSIF x = 16461 THEN
            sigmoid_f := 2047;
        ELSIF x = 16462 THEN
            sigmoid_f := 2047;
        ELSIF x = 16463 THEN
            sigmoid_f := 2047;
        ELSIF x = 16464 THEN
            sigmoid_f := 2047;
        ELSIF x = 16465 THEN
            sigmoid_f := 2047;
        ELSIF x = 16466 THEN
            sigmoid_f := 2047;
        ELSIF x = 16467 THEN
            sigmoid_f := 2047;
        ELSIF x = 16468 THEN
            sigmoid_f := 2047;
        ELSIF x = 16469 THEN
            sigmoid_f := 2047;
        ELSIF x = 16470 THEN
            sigmoid_f := 2047;
        ELSIF x = 16471 THEN
            sigmoid_f := 2047;
        ELSIF x = 16472 THEN
            sigmoid_f := 2047;
        ELSIF x = 16473 THEN
            sigmoid_f := 2047;
        ELSIF x = 16474 THEN
            sigmoid_f := 2047;
        ELSIF x = 16475 THEN
            sigmoid_f := 2047;
        ELSIF x = 16476 THEN
            sigmoid_f := 2047;
        ELSIF x = 16477 THEN
            sigmoid_f := 2047;
        ELSIF x = 16478 THEN
            sigmoid_f := 2047;
        ELSIF x = 16479 THEN
            sigmoid_f := 2047;
        ELSIF x = 16480 THEN
            sigmoid_f := 2047;
        ELSIF x = 16481 THEN
            sigmoid_f := 2047;
        ELSIF x = 16482 THEN
            sigmoid_f := 2047;
        ELSIF x = 16483 THEN
            sigmoid_f := 2047;
        ELSIF x = 16484 THEN
            sigmoid_f := 2047;
        ELSIF x = 16485 THEN
            sigmoid_f := 2047;
        ELSIF x = 16486 THEN
            sigmoid_f := 2047;
        ELSIF x = 16487 THEN
            sigmoid_f := 2047;
        ELSIF x = 16488 THEN
            sigmoid_f := 2047;
        ELSIF x = 16489 THEN
            sigmoid_f := 2047;
        ELSIF x = 16490 THEN
            sigmoid_f := 2047;
        ELSIF x = 16491 THEN
            sigmoid_f := 2047;
        ELSIF x = 16492 THEN
            sigmoid_f := 2047;
        ELSIF x = 16493 THEN
            sigmoid_f := 2047;
        ELSIF x = 16494 THEN
            sigmoid_f := 2047;
        ELSIF x = 16495 THEN
            sigmoid_f := 2047;
        ELSIF x = 16496 THEN
            sigmoid_f := 2047;
        ELSIF x = 16497 THEN
            sigmoid_f := 2047;
        ELSIF x = 16498 THEN
            sigmoid_f := 2047;
        ELSIF x = 16499 THEN
            sigmoid_f := 2047;
        ELSIF x = 16500 THEN
            sigmoid_f := 2047;
        ELSIF x = 16501 THEN
            sigmoid_f := 2047;
        ELSIF x = 16502 THEN
            sigmoid_f := 2047;
        ELSIF x = 16503 THEN
            sigmoid_f := 2047;
        ELSIF x = 16504 THEN
            sigmoid_f := 2047;
        ELSIF x = 16505 THEN
            sigmoid_f := 2047;
        ELSIF x = 16506 THEN
            sigmoid_f := 2047;
        ELSIF x = 16507 THEN
            sigmoid_f := 2047;
        ELSIF x = 16508 THEN
            sigmoid_f := 2047;
        ELSIF x = 16509 THEN
            sigmoid_f := 2047;
        ELSIF x = 16510 THEN
            sigmoid_f := 2047;
        ELSIF x = 16511 THEN
            sigmoid_f := 2047;
        ELSIF x = 16512 THEN
            sigmoid_f := 2047;
        ELSIF x = 16513 THEN
            sigmoid_f := 2047;
        ELSIF x = 16514 THEN
            sigmoid_f := 2047;
        ELSIF x = 16515 THEN
            sigmoid_f := 2047;
        ELSIF x = 16516 THEN
            sigmoid_f := 2047;
        ELSIF x = 16517 THEN
            sigmoid_f := 2047;
        ELSIF x = 16518 THEN
            sigmoid_f := 2047;
        ELSIF x = 16519 THEN
            sigmoid_f := 2047;
        ELSIF x = 16520 THEN
            sigmoid_f := 2047;
        ELSIF x = 16521 THEN
            sigmoid_f := 2047;
        ELSIF x = 16522 THEN
            sigmoid_f := 2047;
        ELSIF x = 16523 THEN
            sigmoid_f := 2047;
        ELSIF x = 16524 THEN
            sigmoid_f := 2047;
        ELSIF x = 16525 THEN
            sigmoid_f := 2047;
        ELSIF x = 16526 THEN
            sigmoid_f := 2047;
        ELSIF x = 16527 THEN
            sigmoid_f := 2047;
        ELSIF x = 16528 THEN
            sigmoid_f := 2047;
        ELSIF x = 16529 THEN
            sigmoid_f := 2047;
        ELSIF x = 16530 THEN
            sigmoid_f := 2047;
        ELSIF x = 16531 THEN
            sigmoid_f := 2047;
        ELSIF x = 16532 THEN
            sigmoid_f := 2047;
        ELSIF x = 16533 THEN
            sigmoid_f := 2047;
        ELSIF x = 16534 THEN
            sigmoid_f := 2047;
        ELSIF x = 16535 THEN
            sigmoid_f := 2047;
        ELSIF x = 16536 THEN
            sigmoid_f := 2047;
        ELSIF x = 16537 THEN
            sigmoid_f := 2047;
        ELSIF x = 16538 THEN
            sigmoid_f := 2047;
        ELSIF x = 16539 THEN
            sigmoid_f := 2047;
        ELSIF x = 16540 THEN
            sigmoid_f := 2047;
        ELSIF x = 16541 THEN
            sigmoid_f := 2047;
        ELSIF x = 16542 THEN
            sigmoid_f := 2047;
        ELSIF x = 16543 THEN
            sigmoid_f := 2047;
        ELSIF x = 16544 THEN
            sigmoid_f := 2047;
        ELSIF x = 16545 THEN
            sigmoid_f := 2047;
        ELSIF x = 16546 THEN
            sigmoid_f := 2047;
        ELSIF x = 16547 THEN
            sigmoid_f := 2047;
        ELSIF x = 16548 THEN
            sigmoid_f := 2047;
        ELSIF x = 16549 THEN
            sigmoid_f := 2047;
        ELSIF x = 16550 THEN
            sigmoid_f := 2047;
        ELSIF x = 16551 THEN
            sigmoid_f := 2047;
        ELSIF x = 16552 THEN
            sigmoid_f := 2047;
        ELSIF x = 16553 THEN
            sigmoid_f := 2047;
        ELSIF x = 16554 THEN
            sigmoid_f := 2047;
        ELSIF x = 16555 THEN
            sigmoid_f := 2047;
        ELSIF x = 16556 THEN
            sigmoid_f := 2047;
        ELSIF x = 16557 THEN
            sigmoid_f := 2047;
        ELSIF x = 16558 THEN
            sigmoid_f := 2047;
        ELSIF x = 16559 THEN
            sigmoid_f := 2047;
        ELSIF x = 16560 THEN
            sigmoid_f := 2047;
        ELSIF x = 16561 THEN
            sigmoid_f := 2047;
        ELSIF x = 16562 THEN
            sigmoid_f := 2047;
        ELSIF x = 16563 THEN
            sigmoid_f := 2047;
        ELSIF x = 16564 THEN
            sigmoid_f := 2047;
        ELSIF x = 16565 THEN
            sigmoid_f := 2047;
        ELSIF x = 16566 THEN
            sigmoid_f := 2047;
        ELSIF x = 16567 THEN
            sigmoid_f := 2047;
        ELSIF x = 16568 THEN
            sigmoid_f := 2047;
        ELSIF x = 16569 THEN
            sigmoid_f := 2047;
        ELSIF x = 16570 THEN
            sigmoid_f := 2047;
        ELSIF x = 16571 THEN
            sigmoid_f := 2047;
        ELSIF x = 16572 THEN
            sigmoid_f := 2047;
        ELSIF x = 16573 THEN
            sigmoid_f := 2047;
        ELSIF x = 16574 THEN
            sigmoid_f := 2047;
        ELSIF x = 16575 THEN
            sigmoid_f := 2047;
        ELSIF x = 16576 THEN
            sigmoid_f := 2047;
        ELSIF x = 16577 THEN
            sigmoid_f := 2047;
        ELSIF x = 16578 THEN
            sigmoid_f := 2047;
        ELSIF x = 16579 THEN
            sigmoid_f := 2047;
        ELSIF x = 16580 THEN
            sigmoid_f := 2047;
        ELSIF x = 16581 THEN
            sigmoid_f := 2047;
        ELSIF x = 16582 THEN
            sigmoid_f := 2047;
        ELSIF x = 16583 THEN
            sigmoid_f := 2047;
        ELSIF x = 16584 THEN
            sigmoid_f := 2047;
        ELSIF x = 16585 THEN
            sigmoid_f := 2047;
        ELSIF x = 16586 THEN
            sigmoid_f := 2047;
        ELSIF x = 16587 THEN
            sigmoid_f := 2047;
        ELSIF x = 16588 THEN
            sigmoid_f := 2047;
        ELSIF x = 16589 THEN
            sigmoid_f := 2047;
        ELSIF x = 16590 THEN
            sigmoid_f := 2047;
        ELSIF x = 16591 THEN
            sigmoid_f := 2047;
        ELSIF x = 16592 THEN
            sigmoid_f := 2047;
        ELSIF x = 16593 THEN
            sigmoid_f := 2047;
        ELSIF x = 16594 THEN
            sigmoid_f := 2047;
        ELSIF x = 16595 THEN
            sigmoid_f := 2047;
        ELSIF x = 16596 THEN
            sigmoid_f := 2047;
        ELSIF x = 16597 THEN
            sigmoid_f := 2047;
        ELSIF x = 16598 THEN
            sigmoid_f := 2047;
        ELSIF x = 16599 THEN
            sigmoid_f := 2047;
        ELSIF x = 16600 THEN
            sigmoid_f := 2047;
        ELSIF x = 16601 THEN
            sigmoid_f := 2047;
        ELSIF x = 16602 THEN
            sigmoid_f := 2047;
        ELSIF x = 16603 THEN
            sigmoid_f := 2047;
        ELSIF x = 16604 THEN
            sigmoid_f := 2047;
        ELSIF x = 16605 THEN
            sigmoid_f := 2047;
        ELSIF x = 16606 THEN
            sigmoid_f := 2047;
        ELSIF x = 16607 THEN
            sigmoid_f := 2047;
        ELSIF x = 16608 THEN
            sigmoid_f := 2047;
        ELSIF x = 16609 THEN
            sigmoid_f := 2047;
        ELSIF x = 16610 THEN
            sigmoid_f := 2047;
        ELSIF x = 16611 THEN
            sigmoid_f := 2047;
        ELSIF x = 16612 THEN
            sigmoid_f := 2047;
        ELSIF x = 16613 THEN
            sigmoid_f := 2047;
        ELSIF x = 16614 THEN
            sigmoid_f := 2047;
        ELSIF x = 16615 THEN
            sigmoid_f := 2047;
        ELSIF x = 16616 THEN
            sigmoid_f := 2047;
        ELSIF x = 16617 THEN
            sigmoid_f := 2047;
        ELSIF x = 16618 THEN
            sigmoid_f := 2047;
        ELSIF x = 16619 THEN
            sigmoid_f := 2047;
        ELSIF x = 16620 THEN
            sigmoid_f := 2047;
        ELSIF x = 16621 THEN
            sigmoid_f := 2047;
        ELSIF x = 16622 THEN
            sigmoid_f := 2047;
        ELSIF x = 16623 THEN
            sigmoid_f := 2047;
        ELSIF x = 16624 THEN
            sigmoid_f := 2047;
        ELSIF x = 16625 THEN
            sigmoid_f := 2047;
        ELSIF x = 16626 THEN
            sigmoid_f := 2047;
        ELSIF x = 16627 THEN
            sigmoid_f := 2047;
        ELSIF x = 16628 THEN
            sigmoid_f := 2047;
        ELSIF x = 16629 THEN
            sigmoid_f := 2047;
        ELSIF x = 16630 THEN
            sigmoid_f := 2047;
        ELSIF x = 16631 THEN
            sigmoid_f := 2047;
        ELSIF x = 16632 THEN
            sigmoid_f := 2047;
        ELSIF x = 16633 THEN
            sigmoid_f := 2047;
        ELSIF x = 16634 THEN
            sigmoid_f := 2047;
        ELSIF x = 16635 THEN
            sigmoid_f := 2047;
        ELSIF x = 16636 THEN
            sigmoid_f := 2047;
        ELSIF x = 16637 THEN
            sigmoid_f := 2047;
        ELSIF x = 16638 THEN
            sigmoid_f := 2047;
        ELSIF x = 16639 THEN
            sigmoid_f := 2047;
        ELSIF x = 16640 THEN
            sigmoid_f := 2047;
        ELSIF x = 16641 THEN
            sigmoid_f := 2047;
        ELSIF x = 16642 THEN
            sigmoid_f := 2047;
        ELSIF x = 16643 THEN
            sigmoid_f := 2047;
        ELSIF x = 16644 THEN
            sigmoid_f := 2047;
        ELSIF x = 16645 THEN
            sigmoid_f := 2047;
        ELSIF x = 16646 THEN
            sigmoid_f := 2047;
        ELSIF x = 16647 THEN
            sigmoid_f := 2047;
        ELSIF x = 16648 THEN
            sigmoid_f := 2047;
        ELSIF x = 16649 THEN
            sigmoid_f := 2047;
        ELSIF x = 16650 THEN
            sigmoid_f := 2047;
        ELSIF x = 16651 THEN
            sigmoid_f := 2047;
        ELSIF x = 16652 THEN
            sigmoid_f := 2047;
        ELSIF x = 16653 THEN
            sigmoid_f := 2047;
        ELSIF x = 16654 THEN
            sigmoid_f := 2047;
        ELSIF x = 16655 THEN
            sigmoid_f := 2047;
        ELSIF x = 16656 THEN
            sigmoid_f := 2047;
        ELSIF x = 16657 THEN
            sigmoid_f := 2047;
        ELSIF x = 16658 THEN
            sigmoid_f := 2047;
        ELSIF x = 16659 THEN
            sigmoid_f := 2047;
        ELSIF x = 16660 THEN
            sigmoid_f := 2047;
        ELSIF x = 16661 THEN
            sigmoid_f := 2047;
        ELSIF x = 16662 THEN
            sigmoid_f := 2047;
        ELSIF x = 16663 THEN
            sigmoid_f := 2047;
        ELSIF x = 16664 THEN
            sigmoid_f := 2047;
        ELSIF x = 16665 THEN
            sigmoid_f := 2047;
        ELSIF x = 16666 THEN
            sigmoid_f := 2047;
        ELSIF x = 16667 THEN
            sigmoid_f := 2047;
        ELSIF x = 16668 THEN
            sigmoid_f := 2047;
        ELSIF x = 16669 THEN
            sigmoid_f := 2047;
        ELSIF x = 16670 THEN
            sigmoid_f := 2047;
        ELSIF x = 16671 THEN
            sigmoid_f := 2047;
        ELSIF x = 16672 THEN
            sigmoid_f := 2047;
        ELSIF x = 16673 THEN
            sigmoid_f := 2047;
        ELSIF x = 16674 THEN
            sigmoid_f := 2047;
        ELSIF x = 16675 THEN
            sigmoid_f := 2047;
        ELSIF x = 16676 THEN
            sigmoid_f := 2047;
        ELSIF x = 16677 THEN
            sigmoid_f := 2047;
        ELSIF x = 16678 THEN
            sigmoid_f := 2047;
        ELSIF x = 16679 THEN
            sigmoid_f := 2047;
        ELSIF x = 16680 THEN
            sigmoid_f := 2047;
        ELSIF x = 16681 THEN
            sigmoid_f := 2047;
        ELSIF x = 16682 THEN
            sigmoid_f := 2047;
        ELSIF x = 16683 THEN
            sigmoid_f := 2047;
        ELSIF x = 16684 THEN
            sigmoid_f := 2047;
        ELSIF x = 16685 THEN
            sigmoid_f := 2047;
        ELSIF x = 16686 THEN
            sigmoid_f := 2047;
        ELSIF x = 16687 THEN
            sigmoid_f := 2047;
        ELSIF x = 16688 THEN
            sigmoid_f := 2047;
        ELSIF x = 16689 THEN
            sigmoid_f := 2047;
        ELSIF x = 16690 THEN
            sigmoid_f := 2047;
        ELSIF x = 16691 THEN
            sigmoid_f := 2047;
        ELSIF x = 16692 THEN
            sigmoid_f := 2047;
        ELSIF x = 16693 THEN
            sigmoid_f := 2047;
        ELSIF x = 16694 THEN
            sigmoid_f := 2047;
        ELSIF x = 16695 THEN
            sigmoid_f := 2047;
        ELSIF x = 16696 THEN
            sigmoid_f := 2047;
        ELSIF x = 16697 THEN
            sigmoid_f := 2047;
        ELSIF x = 16698 THEN
            sigmoid_f := 2047;
        ELSIF x = 16699 THEN
            sigmoid_f := 2047;
        ELSIF x = 16700 THEN
            sigmoid_f := 2047;
        ELSIF x = 16701 THEN
            sigmoid_f := 2047;
        ELSIF x = 16702 THEN
            sigmoid_f := 2047;
        ELSIF x = 16703 THEN
            sigmoid_f := 2047;
        ELSIF x = 16704 THEN
            sigmoid_f := 2047;
        ELSIF x = 16705 THEN
            sigmoid_f := 2047;
        ELSIF x = 16706 THEN
            sigmoid_f := 2047;
        ELSIF x = 16707 THEN
            sigmoid_f := 2047;
        ELSIF x = 16708 THEN
            sigmoid_f := 2047;
        ELSIF x = 16709 THEN
            sigmoid_f := 2047;
        ELSIF x = 16710 THEN
            sigmoid_f := 2047;
        ELSIF x = 16711 THEN
            sigmoid_f := 2047;
        ELSIF x = 16712 THEN
            sigmoid_f := 2047;
        ELSIF x = 16713 THEN
            sigmoid_f := 2047;
        ELSIF x = 16714 THEN
            sigmoid_f := 2047;
        ELSIF x = 16715 THEN
            sigmoid_f := 2047;
        ELSIF x = 16716 THEN
            sigmoid_f := 2047;
        ELSIF x = 16717 THEN
            sigmoid_f := 2047;
        ELSIF x = 16718 THEN
            sigmoid_f := 2047;
        ELSIF x = 16719 THEN
            sigmoid_f := 2047;
        ELSIF x = 16720 THEN
            sigmoid_f := 2047;
        ELSIF x = 16721 THEN
            sigmoid_f := 2047;
        ELSIF x = 16722 THEN
            sigmoid_f := 2047;
        ELSIF x = 16723 THEN
            sigmoid_f := 2047;
        ELSIF x = 16724 THEN
            sigmoid_f := 2047;
        ELSIF x = 16725 THEN
            sigmoid_f := 2047;
        ELSIF x = 16726 THEN
            sigmoid_f := 2047;
        ELSIF x = 16727 THEN
            sigmoid_f := 2047;
        ELSIF x = 16728 THEN
            sigmoid_f := 2047;
        ELSIF x = 16729 THEN
            sigmoid_f := 2047;
        ELSIF x = 16730 THEN
            sigmoid_f := 2047;
        ELSIF x = 16731 THEN
            sigmoid_f := 2047;
        ELSIF x = 16732 THEN
            sigmoid_f := 2047;
        ELSIF x = 16733 THEN
            sigmoid_f := 2047;
        ELSIF x = 16734 THEN
            sigmoid_f := 2047;
        ELSIF x = 16735 THEN
            sigmoid_f := 2047;
        ELSIF x = 16736 THEN
            sigmoid_f := 2047;
        ELSIF x = 16737 THEN
            sigmoid_f := 2047;
        ELSIF x = 16738 THEN
            sigmoid_f := 2047;
        ELSIF x = 16739 THEN
            sigmoid_f := 2047;
        ELSIF x = 16740 THEN
            sigmoid_f := 2047;
        ELSIF x = 16741 THEN
            sigmoid_f := 2047;
        ELSIF x = 16742 THEN
            sigmoid_f := 2047;
        ELSIF x = 16743 THEN
            sigmoid_f := 2047;
        ELSIF x = 16744 THEN
            sigmoid_f := 2047;
        ELSIF x = 16745 THEN
            sigmoid_f := 2047;
        ELSIF x = 16746 THEN
            sigmoid_f := 2047;
        ELSIF x = 16747 THEN
            sigmoid_f := 2047;
        ELSIF x = 16748 THEN
            sigmoid_f := 2047;
        ELSIF x = 16749 THEN
            sigmoid_f := 2047;
        ELSIF x = 16750 THEN
            sigmoid_f := 2047;
        ELSIF x = 16751 THEN
            sigmoid_f := 2047;
        ELSIF x = 16752 THEN
            sigmoid_f := 2047;
        ELSIF x = 16753 THEN
            sigmoid_f := 2047;
        ELSIF x = 16754 THEN
            sigmoid_f := 2047;
        ELSIF x = 16755 THEN
            sigmoid_f := 2047;
        ELSIF x = 16756 THEN
            sigmoid_f := 2047;
        ELSIF x = 16757 THEN
            sigmoid_f := 2047;
        ELSIF x = 16758 THEN
            sigmoid_f := 2047;
        ELSIF x = 16759 THEN
            sigmoid_f := 2047;
        ELSIF x = 16760 THEN
            sigmoid_f := 2047;
        ELSIF x = 16761 THEN
            sigmoid_f := 2047;
        ELSIF x = 16762 THEN
            sigmoid_f := 2047;
        ELSIF x = 16763 THEN
            sigmoid_f := 2047;
        ELSIF x = 16764 THEN
            sigmoid_f := 2047;
        ELSIF x = 16765 THEN
            sigmoid_f := 2047;
        ELSIF x = 16766 THEN
            sigmoid_f := 2047;
        ELSIF x = 16767 THEN
            sigmoid_f := 2047;
        ELSIF x = 16768 THEN
            sigmoid_f := 2047;
        ELSIF x = 16769 THEN
            sigmoid_f := 2047;
        ELSIF x = 16770 THEN
            sigmoid_f := 2047;
        ELSIF x = 16771 THEN
            sigmoid_f := 2047;
        ELSIF x = 16772 THEN
            sigmoid_f := 2047;
        ELSIF x = 16773 THEN
            sigmoid_f := 2047;
        ELSIF x = 16774 THEN
            sigmoid_f := 2047;
        ELSIF x = 16775 THEN
            sigmoid_f := 2047;
        ELSIF x = 16776 THEN
            sigmoid_f := 2047;
        ELSIF x = 16777 THEN
            sigmoid_f := 2047;
        ELSIF x = 16778 THEN
            sigmoid_f := 2047;
        ELSIF x = 16779 THEN
            sigmoid_f := 2047;
        ELSIF x = 16780 THEN
            sigmoid_f := 2047;
        ELSIF x = 16781 THEN
            sigmoid_f := 2047;
        ELSIF x = 16782 THEN
            sigmoid_f := 2047;
        ELSIF x = 16783 THEN
            sigmoid_f := 2047;
        ELSIF x = 16784 THEN
            sigmoid_f := 2047;
        ELSIF x = 16785 THEN
            sigmoid_f := 2047;
        ELSIF x = 16786 THEN
            sigmoid_f := 2047;
        ELSIF x = 16787 THEN
            sigmoid_f := 2047;
        ELSIF x = 16788 THEN
            sigmoid_f := 2047;
        ELSIF x = 16789 THEN
            sigmoid_f := 2047;
        ELSIF x = 16790 THEN
            sigmoid_f := 2047;
        ELSIF x = 16791 THEN
            sigmoid_f := 2047;
        ELSIF x = 16792 THEN
            sigmoid_f := 2047;
        ELSIF x = 16793 THEN
            sigmoid_f := 2047;
        ELSIF x = 16794 THEN
            sigmoid_f := 2047;
        ELSIF x = 16795 THEN
            sigmoid_f := 2047;
        ELSIF x = 16796 THEN
            sigmoid_f := 2047;
        ELSIF x = 16797 THEN
            sigmoid_f := 2047;
        ELSIF x = 16798 THEN
            sigmoid_f := 2047;
        ELSIF x = 16799 THEN
            sigmoid_f := 2047;
        ELSIF x = 16800 THEN
            sigmoid_f := 2047;
        ELSIF x = 16801 THEN
            sigmoid_f := 2047;
        ELSIF x = 16802 THEN
            sigmoid_f := 2047;
        ELSIF x = 16803 THEN
            sigmoid_f := 2047;
        ELSIF x = 16804 THEN
            sigmoid_f := 2047;
        ELSIF x = 16805 THEN
            sigmoid_f := 2047;
        ELSIF x = 16806 THEN
            sigmoid_f := 2047;
        ELSIF x = 16807 THEN
            sigmoid_f := 2047;
        ELSIF x = 16808 THEN
            sigmoid_f := 2047;
        ELSIF x = 16809 THEN
            sigmoid_f := 2047;
        ELSIF x = 16810 THEN
            sigmoid_f := 2047;
        ELSIF x = 16811 THEN
            sigmoid_f := 2047;
        ELSIF x = 16812 THEN
            sigmoid_f := 2047;
        ELSIF x = 16813 THEN
            sigmoid_f := 2047;
        ELSIF x = 16814 THEN
            sigmoid_f := 2047;
        ELSIF x = 16815 THEN
            sigmoid_f := 2047;
        ELSIF x = 16816 THEN
            sigmoid_f := 2047;
        ELSIF x = 16817 THEN
            sigmoid_f := 2047;
        ELSIF x = 16818 THEN
            sigmoid_f := 2047;
        ELSIF x = 16819 THEN
            sigmoid_f := 2047;
        ELSIF x = 16820 THEN
            sigmoid_f := 2047;
        ELSIF x = 16821 THEN
            sigmoid_f := 2047;
        ELSIF x = 16822 THEN
            sigmoid_f := 2047;
        ELSIF x = 16823 THEN
            sigmoid_f := 2047;
        ELSIF x = 16824 THEN
            sigmoid_f := 2047;
        ELSIF x = 16825 THEN
            sigmoid_f := 2047;
        ELSIF x = 16826 THEN
            sigmoid_f := 2047;
        ELSIF x = 16827 THEN
            sigmoid_f := 2047;
        ELSIF x = 16828 THEN
            sigmoid_f := 2047;
        ELSIF x = 16829 THEN
            sigmoid_f := 2047;
        ELSIF x = 16830 THEN
            sigmoid_f := 2047;
        ELSIF x = 16831 THEN
            sigmoid_f := 2047;
        ELSIF x = 16832 THEN
            sigmoid_f := 2047;
        ELSIF x = 16833 THEN
            sigmoid_f := 2047;
        ELSIF x = 16834 THEN
            sigmoid_f := 2047;
        ELSIF x = 16835 THEN
            sigmoid_f := 2047;
        ELSIF x = 16836 THEN
            sigmoid_f := 2047;
        ELSIF x = 16837 THEN
            sigmoid_f := 2047;
        ELSIF x = 16838 THEN
            sigmoid_f := 2047;
        ELSIF x = 16839 THEN
            sigmoid_f := 2047;
        ELSIF x = 16840 THEN
            sigmoid_f := 2047;
        ELSIF x = 16841 THEN
            sigmoid_f := 2047;
        ELSIF x = 16842 THEN
            sigmoid_f := 2047;
        ELSIF x = 16843 THEN
            sigmoid_f := 2047;
        ELSIF x = 16844 THEN
            sigmoid_f := 2047;
        ELSIF x = 16845 THEN
            sigmoid_f := 2047;
        ELSIF x = 16846 THEN
            sigmoid_f := 2047;
        ELSIF x = 16847 THEN
            sigmoid_f := 2047;
        ELSIF x = 16848 THEN
            sigmoid_f := 2047;
        ELSIF x = 16849 THEN
            sigmoid_f := 2047;
        ELSIF x = 16850 THEN
            sigmoid_f := 2047;
        ELSIF x = 16851 THEN
            sigmoid_f := 2047;
        ELSIF x = 16852 THEN
            sigmoid_f := 2047;
        ELSIF x = 16853 THEN
            sigmoid_f := 2047;
        ELSIF x = 16854 THEN
            sigmoid_f := 2047;
        ELSIF x = 16855 THEN
            sigmoid_f := 2047;
        ELSIF x = 16856 THEN
            sigmoid_f := 2047;
        ELSIF x = 16857 THEN
            sigmoid_f := 2047;
        ELSIF x = 16858 THEN
            sigmoid_f := 2047;
        ELSIF x = 16859 THEN
            sigmoid_f := 2047;
        ELSIF x = 16860 THEN
            sigmoid_f := 2047;
        ELSIF x = 16861 THEN
            sigmoid_f := 2047;
        ELSIF x = 16862 THEN
            sigmoid_f := 2047;
        ELSIF x = 16863 THEN
            sigmoid_f := 2047;
        ELSIF x = 16864 THEN
            sigmoid_f := 2047;
        ELSIF x = 16865 THEN
            sigmoid_f := 2047;
        ELSIF x = 16866 THEN
            sigmoid_f := 2047;
        ELSIF x = 16867 THEN
            sigmoid_f := 2047;
        ELSIF x = 16868 THEN
            sigmoid_f := 2047;
        ELSIF x = 16869 THEN
            sigmoid_f := 2047;
        ELSIF x = 16870 THEN
            sigmoid_f := 2047;
        ELSIF x = 16871 THEN
            sigmoid_f := 2047;
        ELSIF x = 16872 THEN
            sigmoid_f := 2047;
        ELSIF x = 16873 THEN
            sigmoid_f := 2047;
        ELSIF x = 16874 THEN
            sigmoid_f := 2047;
        ELSIF x = 16875 THEN
            sigmoid_f := 2047;
        ELSIF x = 16876 THEN
            sigmoid_f := 2047;
        ELSIF x = 16877 THEN
            sigmoid_f := 2047;
        ELSIF x = 16878 THEN
            sigmoid_f := 2047;
        ELSIF x = 16879 THEN
            sigmoid_f := 2047;
        ELSIF x = 16880 THEN
            sigmoid_f := 2047;
        ELSIF x = 16881 THEN
            sigmoid_f := 2047;
        ELSIF x = 16882 THEN
            sigmoid_f := 2047;
        ELSIF x = 16883 THEN
            sigmoid_f := 2047;
        ELSIF x = 16884 THEN
            sigmoid_f := 2047;
        ELSIF x = 16885 THEN
            sigmoid_f := 2047;
        ELSIF x = 16886 THEN
            sigmoid_f := 2047;
        ELSIF x = 16887 THEN
            sigmoid_f := 2047;
        ELSIF x = 16888 THEN
            sigmoid_f := 2047;
        ELSIF x = 16889 THEN
            sigmoid_f := 2047;
        ELSIF x = 16890 THEN
            sigmoid_f := 2047;
        ELSIF x = 16891 THEN
            sigmoid_f := 2047;
        ELSIF x = 16892 THEN
            sigmoid_f := 2047;
        ELSIF x = 16893 THEN
            sigmoid_f := 2047;
        ELSIF x = 16894 THEN
            sigmoid_f := 2047;
        ELSIF x = 16895 THEN
            sigmoid_f := 2047;
        ELSIF x >= 16896 THEN
            sigmoid_f := 2048;
        END IF;
        RETURN sigmoid_f;
    END;
END PACKAGE BODY sigmoid_pkg;