-------------------------------------------------------
--! @file tanh_pkg.vhd
--! @brief Package Containing the lut for tanh (matlab generated)
--! @details 
--! @author Guido Baccelli
--! @version 1.0
--! @date 23/08/2019
--! @bug NONE
--! @todo NONE
--! @copyright  GNU Public License [GPL-3.0].
-------------------------------------------------------
---------------- Copyright (c) notice -----------------------------------------
--
-- The VHDL code, the logic and concepts described in this file constitute
-- the intellectual property of the authors listed below, who are affiliated
-- to KTH(Kungliga Tekniska Högskolan), School of ICT, Kista.
-- Any unauthorised use, copy or distribution is strictly prohibited.
-- Any authorised use, copy or distribution should carry this copyright notice
-- unaltered.
-------------------------------------------------------------------------------
-- Title      : Package Containing the lut for tanh (matlab generated)
-- Project    : SiLago
-------------------------------------------------------------------------------
-- File       : tanh_pkg.vhd
-- Author     : Guido Baccelli
-- Company    : KTH
-- Created    : 23/08/2019
-- Last update: 23/08/2019
-- Platform   : SiLago
-- Standard   : VHDL'08
-- Supervisor : Dimitrios Stathis
-------------------------------------------------------------------------------
-- Copyright (c) 2019
-------------------------------------------------------------------------------
-- Contact    : Dimitrios Stathis <stathis@kth.se>
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author                  Description
-- 23/08/2019  1.0      Guido Baccelli          Created
-------------------------------------------------------------------------------

--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#
--                                                                         #
--This file is part of SiLago.                                             #
--                                                                         #
--    SiLago platform source code is distributed freely: you can           #
--    redistribute it and/or modify it under the terms of the GNU          #
--    General Public License as published by the Free Software Foundation, #
--    either version 3 of the License, or (at your option) any             #
--    later version.                                                       #
--                                                                         #
--    SiLago is distributed in the hope that it will be useful,            #
--    but WITHOUT ANY WARRANTY; without even the implied warranty of       #
--    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the        #
--    GNU General Public License for more details.                         #
--                                                                         #
--    You should have received a copy of the GNU General Public License    #
--    along with SiLago.  If not, see <https://www.gnu.org/licenses/>.     #
--                                                                         #
--~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~#

--! Standard ieee library
LIBRARY ieee;
--! Standard logic package
USE ieee.std_logic_1164.ALL;
--! Standard numeric package for signed and unsigned
USE ieee.numeric_std.ALL;

--! Package file with Hyperbolic tangent behavior model for testbench

--! The only content is the 'tanh_fp11' function that emulates behavior of Hyperbolic Tangent operation inside 'ann_unit'
PACKAGE tanh_pkg IS

    FUNCTION tanh_fp11(
        x : INTEGER
    ) RETURN INTEGER;

END PACKAGE tanh_pkg;

--! @brief Contains body of function 'tanh_fp11'
--! @details The function 'tanh_fp11' (and the testbench) interpret input and output data words
--! as integer values instead of fixed-point values. This makes the model easier to describe.
--! The function describes the Hyperbolic tangent by assigning the corresponding output to each possible
--! input value representable on Q4.11.
PACKAGE BODY tanh_pkg IS
    FUNCTION tanh_fp11(
        x : INTEGER)
        RETURN INTEGER IS
        VARIABLE tanh_f : INTEGER;
    BEGIN
        IF x <= - 8448 THEN
            tanh_f := - 2048;
        ELSIF x =- 8447 THEN
            tanh_f := - 2046;
        ELSIF x =- 8446 THEN
            tanh_f := - 2046;
        ELSIF x =- 8445 THEN
            tanh_f := - 2046;
        ELSIF x =- 8444 THEN
            tanh_f := - 2046;
        ELSIF x =- 8443 THEN
            tanh_f := - 2046;
        ELSIF x =- 8442 THEN
            tanh_f := - 2046;
        ELSIF x =- 8441 THEN
            tanh_f := - 2046;
        ELSIF x =- 8440 THEN
            tanh_f := - 2046;
        ELSIF x =- 8439 THEN
            tanh_f := - 2046;
        ELSIF x =- 8438 THEN
            tanh_f := - 2046;
        ELSIF x =- 8437 THEN
            tanh_f := - 2046;
        ELSIF x =- 8436 THEN
            tanh_f := - 2046;
        ELSIF x =- 8435 THEN
            tanh_f := - 2046;
        ELSIF x =- 8434 THEN
            tanh_f := - 2046;
        ELSIF x =- 8433 THEN
            tanh_f := - 2046;
        ELSIF x =- 8432 THEN
            tanh_f := - 2046;
        ELSIF x =- 8431 THEN
            tanh_f := - 2046;
        ELSIF x =- 8430 THEN
            tanh_f := - 2046;
        ELSIF x =- 8429 THEN
            tanh_f := - 2046;
        ELSIF x =- 8428 THEN
            tanh_f := - 2046;
        ELSIF x =- 8427 THEN
            tanh_f := - 2046;
        ELSIF x =- 8426 THEN
            tanh_f := - 2046;
        ELSIF x =- 8425 THEN
            tanh_f := - 2046;
        ELSIF x =- 8424 THEN
            tanh_f := - 2046;
        ELSIF x =- 8423 THEN
            tanh_f := - 2046;
        ELSIF x =- 8422 THEN
            tanh_f := - 2046;
        ELSIF x =- 8421 THEN
            tanh_f := - 2046;
        ELSIF x =- 8420 THEN
            tanh_f := - 2046;
        ELSIF x =- 8419 THEN
            tanh_f := - 2046;
        ELSIF x =- 8418 THEN
            tanh_f := - 2046;
        ELSIF x =- 8417 THEN
            tanh_f := - 2046;
        ELSIF x =- 8416 THEN
            tanh_f := - 2046;
        ELSIF x =- 8415 THEN
            tanh_f := - 2046;
        ELSIF x =- 8414 THEN
            tanh_f := - 2046;
        ELSIF x =- 8413 THEN
            tanh_f := - 2046;
        ELSIF x =- 8412 THEN
            tanh_f := - 2046;
        ELSIF x =- 8411 THEN
            tanh_f := - 2046;
        ELSIF x =- 8410 THEN
            tanh_f := - 2046;
        ELSIF x =- 8409 THEN
            tanh_f := - 2046;
        ELSIF x =- 8408 THEN
            tanh_f := - 2046;
        ELSIF x =- 8407 THEN
            tanh_f := - 2046;
        ELSIF x =- 8406 THEN
            tanh_f := - 2046;
        ELSIF x =- 8405 THEN
            tanh_f := - 2046;
        ELSIF x =- 8404 THEN
            tanh_f := - 2046;
        ELSIF x =- 8403 THEN
            tanh_f := - 2046;
        ELSIF x =- 8402 THEN
            tanh_f := - 2046;
        ELSIF x =- 8401 THEN
            tanh_f := - 2046;
        ELSIF x =- 8400 THEN
            tanh_f := - 2046;
        ELSIF x =- 8399 THEN
            tanh_f := - 2046;
        ELSIF x =- 8398 THEN
            tanh_f := - 2046;
        ELSIF x =- 8397 THEN
            tanh_f := - 2046;
        ELSIF x =- 8396 THEN
            tanh_f := - 2046;
        ELSIF x =- 8395 THEN
            tanh_f := - 2046;
        ELSIF x =- 8394 THEN
            tanh_f := - 2046;
        ELSIF x =- 8393 THEN
            tanh_f := - 2046;
        ELSIF x =- 8392 THEN
            tanh_f := - 2046;
        ELSIF x =- 8391 THEN
            tanh_f := - 2046;
        ELSIF x =- 8390 THEN
            tanh_f := - 2046;
        ELSIF x =- 8389 THEN
            tanh_f := - 2046;
        ELSIF x =- 8388 THEN
            tanh_f := - 2046;
        ELSIF x =- 8387 THEN
            tanh_f := - 2046;
        ELSIF x =- 8386 THEN
            tanh_f := - 2046;
        ELSIF x =- 8385 THEN
            tanh_f := - 2046;
        ELSIF x =- 8384 THEN
            tanh_f := - 2046;
        ELSIF x =- 8383 THEN
            tanh_f := - 2046;
        ELSIF x =- 8382 THEN
            tanh_f := - 2046;
        ELSIF x =- 8381 THEN
            tanh_f := - 2046;
        ELSIF x =- 8380 THEN
            tanh_f := - 2046;
        ELSIF x =- 8379 THEN
            tanh_f := - 2046;
        ELSIF x =- 8378 THEN
            tanh_f := - 2046;
        ELSIF x =- 8377 THEN
            tanh_f := - 2046;
        ELSIF x =- 8376 THEN
            tanh_f := - 2046;
        ELSIF x =- 8375 THEN
            tanh_f := - 2046;
        ELSIF x =- 8374 THEN
            tanh_f := - 2046;
        ELSIF x =- 8373 THEN
            tanh_f := - 2046;
        ELSIF x =- 8372 THEN
            tanh_f := - 2046;
        ELSIF x =- 8371 THEN
            tanh_f := - 2046;
        ELSIF x =- 8370 THEN
            tanh_f := - 2046;
        ELSIF x =- 8369 THEN
            tanh_f := - 2046;
        ELSIF x =- 8368 THEN
            tanh_f := - 2046;
        ELSIF x =- 8367 THEN
            tanh_f := - 2046;
        ELSIF x =- 8366 THEN
            tanh_f := - 2046;
        ELSIF x =- 8365 THEN
            tanh_f := - 2046;
        ELSIF x =- 8364 THEN
            tanh_f := - 2046;
        ELSIF x =- 8363 THEN
            tanh_f := - 2046;
        ELSIF x =- 8362 THEN
            tanh_f := - 2046;
        ELSIF x =- 8361 THEN
            tanh_f := - 2046;
        ELSIF x =- 8360 THEN
            tanh_f := - 2046;
        ELSIF x =- 8359 THEN
            tanh_f := - 2046;
        ELSIF x =- 8358 THEN
            tanh_f := - 2046;
        ELSIF x =- 8357 THEN
            tanh_f := - 2046;
        ELSIF x =- 8356 THEN
            tanh_f := - 2046;
        ELSIF x =- 8355 THEN
            tanh_f := - 2046;
        ELSIF x =- 8354 THEN
            tanh_f := - 2046;
        ELSIF x =- 8353 THEN
            tanh_f := - 2046;
        ELSIF x =- 8352 THEN
            tanh_f := - 2046;
        ELSIF x =- 8351 THEN
            tanh_f := - 2046;
        ELSIF x =- 8350 THEN
            tanh_f := - 2046;
        ELSIF x =- 8349 THEN
            tanh_f := - 2046;
        ELSIF x =- 8348 THEN
            tanh_f := - 2046;
        ELSIF x =- 8347 THEN
            tanh_f := - 2046;
        ELSIF x =- 8346 THEN
            tanh_f := - 2046;
        ELSIF x =- 8345 THEN
            tanh_f := - 2046;
        ELSIF x =- 8344 THEN
            tanh_f := - 2046;
        ELSIF x =- 8343 THEN
            tanh_f := - 2046;
        ELSIF x =- 8342 THEN
            tanh_f := - 2046;
        ELSIF x =- 8341 THEN
            tanh_f := - 2046;
        ELSIF x =- 8340 THEN
            tanh_f := - 2046;
        ELSIF x =- 8339 THEN
            tanh_f := - 2046;
        ELSIF x =- 8338 THEN
            tanh_f := - 2046;
        ELSIF x =- 8337 THEN
            tanh_f := - 2046;
        ELSIF x =- 8336 THEN
            tanh_f := - 2046;
        ELSIF x =- 8335 THEN
            tanh_f := - 2046;
        ELSIF x =- 8334 THEN
            tanh_f := - 2046;
        ELSIF x =- 8333 THEN
            tanh_f := - 2046;
        ELSIF x =- 8332 THEN
            tanh_f := - 2046;
        ELSIF x =- 8331 THEN
            tanh_f := - 2046;
        ELSIF x =- 8330 THEN
            tanh_f := - 2046;
        ELSIF x =- 8329 THEN
            tanh_f := - 2046;
        ELSIF x =- 8328 THEN
            tanh_f := - 2046;
        ELSIF x =- 8327 THEN
            tanh_f := - 2046;
        ELSIF x =- 8326 THEN
            tanh_f := - 2046;
        ELSIF x =- 8325 THEN
            tanh_f := - 2046;
        ELSIF x =- 8324 THEN
            tanh_f := - 2046;
        ELSIF x =- 8323 THEN
            tanh_f := - 2046;
        ELSIF x =- 8322 THEN
            tanh_f := - 2046;
        ELSIF x =- 8321 THEN
            tanh_f := - 2046;
        ELSIF x =- 8320 THEN
            tanh_f := - 2046;
        ELSIF x =- 8319 THEN
            tanh_f := - 2046;
        ELSIF x =- 8318 THEN
            tanh_f := - 2046;
        ELSIF x =- 8317 THEN
            tanh_f := - 2046;
        ELSIF x =- 8316 THEN
            tanh_f := - 2046;
        ELSIF x =- 8315 THEN
            tanh_f := - 2046;
        ELSIF x =- 8314 THEN
            tanh_f := - 2046;
        ELSIF x =- 8313 THEN
            tanh_f := - 2046;
        ELSIF x =- 8312 THEN
            tanh_f := - 2046;
        ELSIF x =- 8311 THEN
            tanh_f := - 2046;
        ELSIF x =- 8310 THEN
            tanh_f := - 2046;
        ELSIF x =- 8309 THEN
            tanh_f := - 2046;
        ELSIF x =- 8308 THEN
            tanh_f := - 2046;
        ELSIF x =- 8307 THEN
            tanh_f := - 2046;
        ELSIF x =- 8306 THEN
            tanh_f := - 2046;
        ELSIF x =- 8305 THEN
            tanh_f := - 2046;
        ELSIF x =- 8304 THEN
            tanh_f := - 2046;
        ELSIF x =- 8303 THEN
            tanh_f := - 2046;
        ELSIF x =- 8302 THEN
            tanh_f := - 2046;
        ELSIF x =- 8301 THEN
            tanh_f := - 2046;
        ELSIF x =- 8300 THEN
            tanh_f := - 2046;
        ELSIF x =- 8299 THEN
            tanh_f := - 2046;
        ELSIF x =- 8298 THEN
            tanh_f := - 2046;
        ELSIF x =- 8297 THEN
            tanh_f := - 2046;
        ELSIF x =- 8296 THEN
            tanh_f := - 2046;
        ELSIF x =- 8295 THEN
            tanh_f := - 2046;
        ELSIF x =- 8294 THEN
            tanh_f := - 2046;
        ELSIF x =- 8293 THEN
            tanh_f := - 2046;
        ELSIF x =- 8292 THEN
            tanh_f := - 2046;
        ELSIF x =- 8291 THEN
            tanh_f := - 2046;
        ELSIF x =- 8290 THEN
            tanh_f := - 2046;
        ELSIF x =- 8289 THEN
            tanh_f := - 2046;
        ELSIF x =- 8288 THEN
            tanh_f := - 2046;
        ELSIF x =- 8287 THEN
            tanh_f := - 2046;
        ELSIF x =- 8286 THEN
            tanh_f := - 2046;
        ELSIF x =- 8285 THEN
            tanh_f := - 2046;
        ELSIF x =- 8284 THEN
            tanh_f := - 2046;
        ELSIF x =- 8283 THEN
            tanh_f := - 2046;
        ELSIF x =- 8282 THEN
            tanh_f := - 2046;
        ELSIF x =- 8281 THEN
            tanh_f := - 2046;
        ELSIF x =- 8280 THEN
            tanh_f := - 2046;
        ELSIF x =- 8279 THEN
            tanh_f := - 2046;
        ELSIF x =- 8278 THEN
            tanh_f := - 2046;
        ELSIF x =- 8277 THEN
            tanh_f := - 2046;
        ELSIF x =- 8276 THEN
            tanh_f := - 2046;
        ELSIF x =- 8275 THEN
            tanh_f := - 2046;
        ELSIF x =- 8274 THEN
            tanh_f := - 2046;
        ELSIF x =- 8273 THEN
            tanh_f := - 2046;
        ELSIF x =- 8272 THEN
            tanh_f := - 2046;
        ELSIF x =- 8271 THEN
            tanh_f := - 2046;
        ELSIF x =- 8270 THEN
            tanh_f := - 2046;
        ELSIF x =- 8269 THEN
            tanh_f := - 2046;
        ELSIF x =- 8268 THEN
            tanh_f := - 2046;
        ELSIF x =- 8267 THEN
            tanh_f := - 2046;
        ELSIF x =- 8266 THEN
            tanh_f := - 2046;
        ELSIF x =- 8265 THEN
            tanh_f := - 2046;
        ELSIF x =- 8264 THEN
            tanh_f := - 2046;
        ELSIF x =- 8263 THEN
            tanh_f := - 2046;
        ELSIF x =- 8262 THEN
            tanh_f := - 2046;
        ELSIF x =- 8261 THEN
            tanh_f := - 2046;
        ELSIF x =- 8260 THEN
            tanh_f := - 2046;
        ELSIF x =- 8259 THEN
            tanh_f := - 2046;
        ELSIF x =- 8258 THEN
            tanh_f := - 2046;
        ELSIF x =- 8257 THEN
            tanh_f := - 2046;
        ELSIF x =- 8256 THEN
            tanh_f := - 2046;
        ELSIF x =- 8255 THEN
            tanh_f := - 2046;
        ELSIF x =- 8254 THEN
            tanh_f := - 2046;
        ELSIF x =- 8253 THEN
            tanh_f := - 2046;
        ELSIF x =- 8252 THEN
            tanh_f := - 2046;
        ELSIF x =- 8251 THEN
            tanh_f := - 2046;
        ELSIF x =- 8250 THEN
            tanh_f := - 2046;
        ELSIF x =- 8249 THEN
            tanh_f := - 2046;
        ELSIF x =- 8248 THEN
            tanh_f := - 2046;
        ELSIF x =- 8247 THEN
            tanh_f := - 2046;
        ELSIF x =- 8246 THEN
            tanh_f := - 2046;
        ELSIF x =- 8245 THEN
            tanh_f := - 2046;
        ELSIF x =- 8244 THEN
            tanh_f := - 2046;
        ELSIF x =- 8243 THEN
            tanh_f := - 2046;
        ELSIF x =- 8242 THEN
            tanh_f := - 2046;
        ELSIF x =- 8241 THEN
            tanh_f := - 2046;
        ELSIF x =- 8240 THEN
            tanh_f := - 2046;
        ELSIF x =- 8239 THEN
            tanh_f := - 2046;
        ELSIF x =- 8238 THEN
            tanh_f := - 2046;
        ELSIF x =- 8237 THEN
            tanh_f := - 2046;
        ELSIF x =- 8236 THEN
            tanh_f := - 2046;
        ELSIF x =- 8235 THEN
            tanh_f := - 2046;
        ELSIF x =- 8234 THEN
            tanh_f := - 2046;
        ELSIF x =- 8233 THEN
            tanh_f := - 2046;
        ELSIF x =- 8232 THEN
            tanh_f := - 2046;
        ELSIF x =- 8231 THEN
            tanh_f := - 2046;
        ELSIF x =- 8230 THEN
            tanh_f := - 2046;
        ELSIF x =- 8229 THEN
            tanh_f := - 2046;
        ELSIF x =- 8228 THEN
            tanh_f := - 2046;
        ELSIF x =- 8227 THEN
            tanh_f := - 2046;
        ELSIF x =- 8226 THEN
            tanh_f := - 2046;
        ELSIF x =- 8225 THEN
            tanh_f := - 2046;
        ELSIF x =- 8224 THEN
            tanh_f := - 2046;
        ELSIF x =- 8223 THEN
            tanh_f := - 2046;
        ELSIF x =- 8222 THEN
            tanh_f := - 2046;
        ELSIF x =- 8221 THEN
            tanh_f := - 2046;
        ELSIF x =- 8220 THEN
            tanh_f := - 2046;
        ELSIF x =- 8219 THEN
            tanh_f := - 2046;
        ELSIF x =- 8218 THEN
            tanh_f := - 2046;
        ELSIF x =- 8217 THEN
            tanh_f := - 2046;
        ELSIF x =- 8216 THEN
            tanh_f := - 2046;
        ELSIF x =- 8215 THEN
            tanh_f := - 2046;
        ELSIF x =- 8214 THEN
            tanh_f := - 2046;
        ELSIF x =- 8213 THEN
            tanh_f := - 2046;
        ELSIF x =- 8212 THEN
            tanh_f := - 2046;
        ELSIF x =- 8211 THEN
            tanh_f := - 2046;
        ELSIF x =- 8210 THEN
            tanh_f := - 2046;
        ELSIF x =- 8209 THEN
            tanh_f := - 2046;
        ELSIF x =- 8208 THEN
            tanh_f := - 2046;
        ELSIF x =- 8207 THEN
            tanh_f := - 2046;
        ELSIF x =- 8206 THEN
            tanh_f := - 2046;
        ELSIF x =- 8205 THEN
            tanh_f := - 2046;
        ELSIF x =- 8204 THEN
            tanh_f := - 2046;
        ELSIF x =- 8203 THEN
            tanh_f := - 2046;
        ELSIF x =- 8202 THEN
            tanh_f := - 2046;
        ELSIF x =- 8201 THEN
            tanh_f := - 2046;
        ELSIF x =- 8200 THEN
            tanh_f := - 2046;
        ELSIF x =- 8199 THEN
            tanh_f := - 2046;
        ELSIF x =- 8198 THEN
            tanh_f := - 2046;
        ELSIF x =- 8197 THEN
            tanh_f := - 2046;
        ELSIF x =- 8196 THEN
            tanh_f := - 2046;
        ELSIF x =- 8195 THEN
            tanh_f := - 2046;
        ELSIF x =- 8194 THEN
            tanh_f := - 2046;
        ELSIF x =- 8193 THEN
            tanh_f := - 2046;
        ELSIF x =- 8192 THEN
            tanh_f := - 2046;
        ELSIF x =- 8191 THEN
            tanh_f := - 2046;
        ELSIF x =- 8190 THEN
            tanh_f := - 2046;
        ELSIF x =- 8189 THEN
            tanh_f := - 2046;
        ELSIF x =- 8188 THEN
            tanh_f := - 2046;
        ELSIF x =- 8187 THEN
            tanh_f := - 2046;
        ELSIF x =- 8186 THEN
            tanh_f := - 2046;
        ELSIF x =- 8185 THEN
            tanh_f := - 2046;
        ELSIF x =- 8184 THEN
            tanh_f := - 2046;
        ELSIF x =- 8183 THEN
            tanh_f := - 2046;
        ELSIF x =- 8182 THEN
            tanh_f := - 2046;
        ELSIF x =- 8181 THEN
            tanh_f := - 2046;
        ELSIF x =- 8180 THEN
            tanh_f := - 2046;
        ELSIF x =- 8179 THEN
            tanh_f := - 2046;
        ELSIF x =- 8178 THEN
            tanh_f := - 2046;
        ELSIF x =- 8177 THEN
            tanh_f := - 2046;
        ELSIF x =- 8176 THEN
            tanh_f := - 2046;
        ELSIF x =- 8175 THEN
            tanh_f := - 2046;
        ELSIF x =- 8174 THEN
            tanh_f := - 2046;
        ELSIF x =- 8173 THEN
            tanh_f := - 2046;
        ELSIF x =- 8172 THEN
            tanh_f := - 2046;
        ELSIF x =- 8171 THEN
            tanh_f := - 2046;
        ELSIF x =- 8170 THEN
            tanh_f := - 2046;
        ELSIF x =- 8169 THEN
            tanh_f := - 2046;
        ELSIF x =- 8168 THEN
            tanh_f := - 2046;
        ELSIF x =- 8167 THEN
            tanh_f := - 2046;
        ELSIF x =- 8166 THEN
            tanh_f := - 2046;
        ELSIF x =- 8165 THEN
            tanh_f := - 2046;
        ELSIF x =- 8164 THEN
            tanh_f := - 2046;
        ELSIF x =- 8163 THEN
            tanh_f := - 2046;
        ELSIF x =- 8162 THEN
            tanh_f := - 2046;
        ELSIF x =- 8161 THEN
            tanh_f := - 2046;
        ELSIF x =- 8160 THEN
            tanh_f := - 2046;
        ELSIF x =- 8159 THEN
            tanh_f := - 2046;
        ELSIF x =- 8158 THEN
            tanh_f := - 2046;
        ELSIF x =- 8157 THEN
            tanh_f := - 2046;
        ELSIF x =- 8156 THEN
            tanh_f := - 2046;
        ELSIF x =- 8155 THEN
            tanh_f := - 2046;
        ELSIF x =- 8154 THEN
            tanh_f := - 2046;
        ELSIF x =- 8153 THEN
            tanh_f := - 2046;
        ELSIF x =- 8152 THEN
            tanh_f := - 2046;
        ELSIF x =- 8151 THEN
            tanh_f := - 2046;
        ELSIF x =- 8150 THEN
            tanh_f := - 2046;
        ELSIF x =- 8149 THEN
            tanh_f := - 2046;
        ELSIF x =- 8148 THEN
            tanh_f := - 2046;
        ELSIF x =- 8147 THEN
            tanh_f := - 2046;
        ELSIF x =- 8146 THEN
            tanh_f := - 2046;
        ELSIF x =- 8145 THEN
            tanh_f := - 2046;
        ELSIF x =- 8144 THEN
            tanh_f := - 2046;
        ELSIF x =- 8143 THEN
            tanh_f := - 2046;
        ELSIF x =- 8142 THEN
            tanh_f := - 2046;
        ELSIF x =- 8141 THEN
            tanh_f := - 2046;
        ELSIF x =- 8140 THEN
            tanh_f := - 2046;
        ELSIF x =- 8139 THEN
            tanh_f := - 2046;
        ELSIF x =- 8138 THEN
            tanh_f := - 2046;
        ELSIF x =- 8137 THEN
            tanh_f := - 2046;
        ELSIF x =- 8136 THEN
            tanh_f := - 2046;
        ELSIF x =- 8135 THEN
            tanh_f := - 2046;
        ELSIF x =- 8134 THEN
            tanh_f := - 2046;
        ELSIF x =- 8133 THEN
            tanh_f := - 2046;
        ELSIF x =- 8132 THEN
            tanh_f := - 2046;
        ELSIF x =- 8131 THEN
            tanh_f := - 2046;
        ELSIF x =- 8130 THEN
            tanh_f := - 2046;
        ELSIF x =- 8129 THEN
            tanh_f := - 2046;
        ELSIF x =- 8128 THEN
            tanh_f := - 2046;
        ELSIF x =- 8127 THEN
            tanh_f := - 2046;
        ELSIF x =- 8126 THEN
            tanh_f := - 2046;
        ELSIF x =- 8125 THEN
            tanh_f := - 2046;
        ELSIF x =- 8124 THEN
            tanh_f := - 2046;
        ELSIF x =- 8123 THEN
            tanh_f := - 2046;
        ELSIF x =- 8122 THEN
            tanh_f := - 2046;
        ELSIF x =- 8121 THEN
            tanh_f := - 2046;
        ELSIF x =- 8120 THEN
            tanh_f := - 2046;
        ELSIF x =- 8119 THEN
            tanh_f := - 2046;
        ELSIF x =- 8118 THEN
            tanh_f := - 2046;
        ELSIF x =- 8117 THEN
            tanh_f := - 2046;
        ELSIF x =- 8116 THEN
            tanh_f := - 2046;
        ELSIF x =- 8115 THEN
            tanh_f := - 2046;
        ELSIF x =- 8114 THEN
            tanh_f := - 2046;
        ELSIF x =- 8113 THEN
            tanh_f := - 2046;
        ELSIF x =- 8112 THEN
            tanh_f := - 2046;
        ELSIF x =- 8111 THEN
            tanh_f := - 2046;
        ELSIF x =- 8110 THEN
            tanh_f := - 2046;
        ELSIF x =- 8109 THEN
            tanh_f := - 2046;
        ELSIF x =- 8108 THEN
            tanh_f := - 2046;
        ELSIF x =- 8107 THEN
            tanh_f := - 2046;
        ELSIF x =- 8106 THEN
            tanh_f := - 2046;
        ELSIF x =- 8105 THEN
            tanh_f := - 2046;
        ELSIF x =- 8104 THEN
            tanh_f := - 2046;
        ELSIF x =- 8103 THEN
            tanh_f := - 2046;
        ELSIF x =- 8102 THEN
            tanh_f := - 2046;
        ELSIF x =- 8101 THEN
            tanh_f := - 2046;
        ELSIF x =- 8100 THEN
            tanh_f := - 2046;
        ELSIF x =- 8099 THEN
            tanh_f := - 2046;
        ELSIF x =- 8098 THEN
            tanh_f := - 2046;
        ELSIF x =- 8097 THEN
            tanh_f := - 2046;
        ELSIF x =- 8096 THEN
            tanh_f := - 2046;
        ELSIF x =- 8095 THEN
            tanh_f := - 2046;
        ELSIF x =- 8094 THEN
            tanh_f := - 2046;
        ELSIF x =- 8093 THEN
            tanh_f := - 2046;
        ELSIF x =- 8092 THEN
            tanh_f := - 2046;
        ELSIF x =- 8091 THEN
            tanh_f := - 2046;
        ELSIF x =- 8090 THEN
            tanh_f := - 2046;
        ELSIF x =- 8089 THEN
            tanh_f := - 2046;
        ELSIF x =- 8088 THEN
            tanh_f := - 2046;
        ELSIF x =- 8087 THEN
            tanh_f := - 2046;
        ELSIF x =- 8086 THEN
            tanh_f := - 2046;
        ELSIF x =- 8085 THEN
            tanh_f := - 2046;
        ELSIF x =- 8084 THEN
            tanh_f := - 2046;
        ELSIF x =- 8083 THEN
            tanh_f := - 2046;
        ELSIF x =- 8082 THEN
            tanh_f := - 2046;
        ELSIF x =- 8081 THEN
            tanh_f := - 2046;
        ELSIF x =- 8080 THEN
            tanh_f := - 2046;
        ELSIF x =- 8079 THEN
            tanh_f := - 2046;
        ELSIF x =- 8078 THEN
            tanh_f := - 2046;
        ELSIF x =- 8077 THEN
            tanh_f := - 2046;
        ELSIF x =- 8076 THEN
            tanh_f := - 2046;
        ELSIF x =- 8075 THEN
            tanh_f := - 2046;
        ELSIF x =- 8074 THEN
            tanh_f := - 2046;
        ELSIF x =- 8073 THEN
            tanh_f := - 2046;
        ELSIF x =- 8072 THEN
            tanh_f := - 2046;
        ELSIF x =- 8071 THEN
            tanh_f := - 2046;
        ELSIF x =- 8070 THEN
            tanh_f := - 2046;
        ELSIF x =- 8069 THEN
            tanh_f := - 2046;
        ELSIF x =- 8068 THEN
            tanh_f := - 2046;
        ELSIF x =- 8067 THEN
            tanh_f := - 2046;
        ELSIF x =- 8066 THEN
            tanh_f := - 2046;
        ELSIF x =- 8065 THEN
            tanh_f := - 2046;
        ELSIF x =- 8064 THEN
            tanh_f := - 2046;
        ELSIF x =- 8063 THEN
            tanh_f := - 2046;
        ELSIF x =- 8062 THEN
            tanh_f := - 2046;
        ELSIF x =- 8061 THEN
            tanh_f := - 2046;
        ELSIF x =- 8060 THEN
            tanh_f := - 2046;
        ELSIF x =- 8059 THEN
            tanh_f := - 2046;
        ELSIF x =- 8058 THEN
            tanh_f := - 2046;
        ELSIF x =- 8057 THEN
            tanh_f := - 2046;
        ELSIF x =- 8056 THEN
            tanh_f := - 2046;
        ELSIF x =- 8055 THEN
            tanh_f := - 2046;
        ELSIF x =- 8054 THEN
            tanh_f := - 2046;
        ELSIF x =- 8053 THEN
            tanh_f := - 2046;
        ELSIF x =- 8052 THEN
            tanh_f := - 2046;
        ELSIF x =- 8051 THEN
            tanh_f := - 2046;
        ELSIF x =- 8050 THEN
            tanh_f := - 2046;
        ELSIF x =- 8049 THEN
            tanh_f := - 2046;
        ELSIF x =- 8048 THEN
            tanh_f := - 2046;
        ELSIF x =- 8047 THEN
            tanh_f := - 2046;
        ELSIF x =- 8046 THEN
            tanh_f := - 2046;
        ELSIF x =- 8045 THEN
            tanh_f := - 2046;
        ELSIF x =- 8044 THEN
            tanh_f := - 2046;
        ELSIF x =- 8043 THEN
            tanh_f := - 2046;
        ELSIF x =- 8042 THEN
            tanh_f := - 2046;
        ELSIF x =- 8041 THEN
            tanh_f := - 2046;
        ELSIF x =- 8040 THEN
            tanh_f := - 2046;
        ELSIF x =- 8039 THEN
            tanh_f := - 2046;
        ELSIF x =- 8038 THEN
            tanh_f := - 2046;
        ELSIF x =- 8037 THEN
            tanh_f := - 2046;
        ELSIF x =- 8036 THEN
            tanh_f := - 2046;
        ELSIF x =- 8035 THEN
            tanh_f := - 2046;
        ELSIF x =- 8034 THEN
            tanh_f := - 2046;
        ELSIF x =- 8033 THEN
            tanh_f := - 2046;
        ELSIF x =- 8032 THEN
            tanh_f := - 2046;
        ELSIF x =- 8031 THEN
            tanh_f := - 2046;
        ELSIF x =- 8030 THEN
            tanh_f := - 2046;
        ELSIF x =- 8029 THEN
            tanh_f := - 2046;
        ELSIF x =- 8028 THEN
            tanh_f := - 2046;
        ELSIF x =- 8027 THEN
            tanh_f := - 2046;
        ELSIF x =- 8026 THEN
            tanh_f := - 2046;
        ELSIF x =- 8025 THEN
            tanh_f := - 2046;
        ELSIF x =- 8024 THEN
            tanh_f := - 2046;
        ELSIF x =- 8023 THEN
            tanh_f := - 2046;
        ELSIF x =- 8022 THEN
            tanh_f := - 2046;
        ELSIF x =- 8021 THEN
            tanh_f := - 2046;
        ELSIF x =- 8020 THEN
            tanh_f := - 2046;
        ELSIF x =- 8019 THEN
            tanh_f := - 2046;
        ELSIF x =- 8018 THEN
            tanh_f := - 2046;
        ELSIF x =- 8017 THEN
            tanh_f := - 2046;
        ELSIF x =- 8016 THEN
            tanh_f := - 2046;
        ELSIF x =- 8015 THEN
            tanh_f := - 2046;
        ELSIF x =- 8014 THEN
            tanh_f := - 2046;
        ELSIF x =- 8013 THEN
            tanh_f := - 2046;
        ELSIF x =- 8012 THEN
            tanh_f := - 2046;
        ELSIF x =- 8011 THEN
            tanh_f := - 2046;
        ELSIF x =- 8010 THEN
            tanh_f := - 2046;
        ELSIF x =- 8009 THEN
            tanh_f := - 2046;
        ELSIF x =- 8008 THEN
            tanh_f := - 2046;
        ELSIF x =- 8007 THEN
            tanh_f := - 2046;
        ELSIF x =- 8006 THEN
            tanh_f := - 2046;
        ELSIF x =- 8005 THEN
            tanh_f := - 2046;
        ELSIF x =- 8004 THEN
            tanh_f := - 2046;
        ELSIF x =- 8003 THEN
            tanh_f := - 2046;
        ELSIF x =- 8002 THEN
            tanh_f := - 2046;
        ELSIF x =- 8001 THEN
            tanh_f := - 2046;
        ELSIF x =- 8000 THEN
            tanh_f := - 2046;
        ELSIF x =- 7999 THEN
            tanh_f := - 2046;
        ELSIF x =- 7998 THEN
            tanh_f := - 2046;
        ELSIF x =- 7997 THEN
            tanh_f := - 2046;
        ELSIF x =- 7996 THEN
            tanh_f := - 2046;
        ELSIF x =- 7995 THEN
            tanh_f := - 2046;
        ELSIF x =- 7994 THEN
            tanh_f := - 2046;
        ELSIF x =- 7993 THEN
            tanh_f := - 2046;
        ELSIF x =- 7992 THEN
            tanh_f := - 2046;
        ELSIF x =- 7991 THEN
            tanh_f := - 2046;
        ELSIF x =- 7990 THEN
            tanh_f := - 2046;
        ELSIF x =- 7989 THEN
            tanh_f := - 2046;
        ELSIF x =- 7988 THEN
            tanh_f := - 2046;
        ELSIF x =- 7987 THEN
            tanh_f := - 2046;
        ELSIF x =- 7986 THEN
            tanh_f := - 2046;
        ELSIF x =- 7985 THEN
            tanh_f := - 2046;
        ELSIF x =- 7984 THEN
            tanh_f := - 2046;
        ELSIF x =- 7983 THEN
            tanh_f := - 2046;
        ELSIF x =- 7982 THEN
            tanh_f := - 2046;
        ELSIF x =- 7981 THEN
            tanh_f := - 2046;
        ELSIF x =- 7980 THEN
            tanh_f := - 2046;
        ELSIF x =- 7979 THEN
            tanh_f := - 2046;
        ELSIF x =- 7978 THEN
            tanh_f := - 2046;
        ELSIF x =- 7977 THEN
            tanh_f := - 2046;
        ELSIF x =- 7976 THEN
            tanh_f := - 2046;
        ELSIF x =- 7975 THEN
            tanh_f := - 2046;
        ELSIF x =- 7974 THEN
            tanh_f := - 2046;
        ELSIF x =- 7973 THEN
            tanh_f := - 2046;
        ELSIF x =- 7972 THEN
            tanh_f := - 2046;
        ELSIF x =- 7971 THEN
            tanh_f := - 2046;
        ELSIF x =- 7970 THEN
            tanh_f := - 2046;
        ELSIF x =- 7969 THEN
            tanh_f := - 2046;
        ELSIF x =- 7968 THEN
            tanh_f := - 2046;
        ELSIF x =- 7967 THEN
            tanh_f := - 2046;
        ELSIF x =- 7966 THEN
            tanh_f := - 2046;
        ELSIF x =- 7965 THEN
            tanh_f := - 2046;
        ELSIF x =- 7964 THEN
            tanh_f := - 2046;
        ELSIF x =- 7963 THEN
            tanh_f := - 2046;
        ELSIF x =- 7962 THEN
            tanh_f := - 2046;
        ELSIF x =- 7961 THEN
            tanh_f := - 2046;
        ELSIF x =- 7960 THEN
            tanh_f := - 2046;
        ELSIF x =- 7959 THEN
            tanh_f := - 2046;
        ELSIF x =- 7958 THEN
            tanh_f := - 2046;
        ELSIF x =- 7957 THEN
            tanh_f := - 2046;
        ELSIF x =- 7956 THEN
            tanh_f := - 2046;
        ELSIF x =- 7955 THEN
            tanh_f := - 2046;
        ELSIF x =- 7954 THEN
            tanh_f := - 2046;
        ELSIF x =- 7953 THEN
            tanh_f := - 2046;
        ELSIF x =- 7952 THEN
            tanh_f := - 2046;
        ELSIF x =- 7951 THEN
            tanh_f := - 2046;
        ELSIF x =- 7950 THEN
            tanh_f := - 2046;
        ELSIF x =- 7949 THEN
            tanh_f := - 2046;
        ELSIF x =- 7948 THEN
            tanh_f := - 2046;
        ELSIF x =- 7947 THEN
            tanh_f := - 2046;
        ELSIF x =- 7946 THEN
            tanh_f := - 2046;
        ELSIF x =- 7945 THEN
            tanh_f := - 2046;
        ELSIF x =- 7944 THEN
            tanh_f := - 2046;
        ELSIF x =- 7943 THEN
            tanh_f := - 2046;
        ELSIF x =- 7942 THEN
            tanh_f := - 2046;
        ELSIF x =- 7941 THEN
            tanh_f := - 2046;
        ELSIF x =- 7940 THEN
            tanh_f := - 2046;
        ELSIF x =- 7939 THEN
            tanh_f := - 2046;
        ELSIF x =- 7938 THEN
            tanh_f := - 2046;
        ELSIF x =- 7937 THEN
            tanh_f := - 2046;
        ELSIF x =- 7936 THEN
            tanh_f := - 2046;
        ELSIF x =- 7935 THEN
            tanh_f := - 2046;
        ELSIF x =- 7934 THEN
            tanh_f := - 2046;
        ELSIF x =- 7933 THEN
            tanh_f := - 2046;
        ELSIF x =- 7932 THEN
            tanh_f := - 2046;
        ELSIF x =- 7931 THEN
            tanh_f := - 2046;
        ELSIF x =- 7930 THEN
            tanh_f := - 2046;
        ELSIF x =- 7929 THEN
            tanh_f := - 2046;
        ELSIF x =- 7928 THEN
            tanh_f := - 2046;
        ELSIF x =- 7927 THEN
            tanh_f := - 2046;
        ELSIF x =- 7926 THEN
            tanh_f := - 2046;
        ELSIF x =- 7925 THEN
            tanh_f := - 2046;
        ELSIF x =- 7924 THEN
            tanh_f := - 2046;
        ELSIF x =- 7923 THEN
            tanh_f := - 2046;
        ELSIF x =- 7922 THEN
            tanh_f := - 2046;
        ELSIF x =- 7921 THEN
            tanh_f := - 2046;
        ELSIF x =- 7920 THEN
            tanh_f := - 2046;
        ELSIF x =- 7919 THEN
            tanh_f := - 2046;
        ELSIF x =- 7918 THEN
            tanh_f := - 2046;
        ELSIF x =- 7917 THEN
            tanh_f := - 2046;
        ELSIF x =- 7916 THEN
            tanh_f := - 2046;
        ELSIF x =- 7915 THEN
            tanh_f := - 2046;
        ELSIF x =- 7914 THEN
            tanh_f := - 2046;
        ELSIF x =- 7913 THEN
            tanh_f := - 2046;
        ELSIF x =- 7912 THEN
            tanh_f := - 2046;
        ELSIF x =- 7911 THEN
            tanh_f := - 2046;
        ELSIF x =- 7910 THEN
            tanh_f := - 2046;
        ELSIF x =- 7909 THEN
            tanh_f := - 2046;
        ELSIF x =- 7908 THEN
            tanh_f := - 2046;
        ELSIF x =- 7907 THEN
            tanh_f := - 2046;
        ELSIF x =- 7906 THEN
            tanh_f := - 2046;
        ELSIF x =- 7905 THEN
            tanh_f := - 2046;
        ELSIF x =- 7904 THEN
            tanh_f := - 2046;
        ELSIF x =- 7903 THEN
            tanh_f := - 2046;
        ELSIF x =- 7902 THEN
            tanh_f := - 2046;
        ELSIF x =- 7901 THEN
            tanh_f := - 2046;
        ELSIF x =- 7900 THEN
            tanh_f := - 2046;
        ELSIF x =- 7899 THEN
            tanh_f := - 2046;
        ELSIF x =- 7898 THEN
            tanh_f := - 2046;
        ELSIF x =- 7897 THEN
            tanh_f := - 2046;
        ELSIF x =- 7896 THEN
            tanh_f := - 2046;
        ELSIF x =- 7895 THEN
            tanh_f := - 2046;
        ELSIF x =- 7894 THEN
            tanh_f := - 2046;
        ELSIF x =- 7893 THEN
            tanh_f := - 2046;
        ELSIF x =- 7892 THEN
            tanh_f := - 2046;
        ELSIF x =- 7891 THEN
            tanh_f := - 2046;
        ELSIF x =- 7890 THEN
            tanh_f := - 2046;
        ELSIF x =- 7889 THEN
            tanh_f := - 2046;
        ELSIF x =- 7888 THEN
            tanh_f := - 2046;
        ELSIF x =- 7887 THEN
            tanh_f := - 2046;
        ELSIF x =- 7886 THEN
            tanh_f := - 2046;
        ELSIF x =- 7885 THEN
            tanh_f := - 2046;
        ELSIF x =- 7884 THEN
            tanh_f := - 2046;
        ELSIF x =- 7883 THEN
            tanh_f := - 2046;
        ELSIF x =- 7882 THEN
            tanh_f := - 2046;
        ELSIF x =- 7881 THEN
            tanh_f := - 2046;
        ELSIF x =- 7880 THEN
            tanh_f := - 2046;
        ELSIF x =- 7879 THEN
            tanh_f := - 2046;
        ELSIF x =- 7878 THEN
            tanh_f := - 2046;
        ELSIF x =- 7877 THEN
            tanh_f := - 2046;
        ELSIF x =- 7876 THEN
            tanh_f := - 2046;
        ELSIF x =- 7875 THEN
            tanh_f := - 2046;
        ELSIF x =- 7874 THEN
            tanh_f := - 2046;
        ELSIF x =- 7873 THEN
            tanh_f := - 2046;
        ELSIF x =- 7872 THEN
            tanh_f := - 2046;
        ELSIF x =- 7871 THEN
            tanh_f := - 2046;
        ELSIF x =- 7870 THEN
            tanh_f := - 2046;
        ELSIF x =- 7869 THEN
            tanh_f := - 2046;
        ELSIF x =- 7868 THEN
            tanh_f := - 2046;
        ELSIF x =- 7867 THEN
            tanh_f := - 2046;
        ELSIF x =- 7866 THEN
            tanh_f := - 2046;
        ELSIF x =- 7865 THEN
            tanh_f := - 2046;
        ELSIF x =- 7864 THEN
            tanh_f := - 2046;
        ELSIF x =- 7863 THEN
            tanh_f := - 2046;
        ELSIF x =- 7862 THEN
            tanh_f := - 2046;
        ELSIF x =- 7861 THEN
            tanh_f := - 2046;
        ELSIF x =- 7860 THEN
            tanh_f := - 2046;
        ELSIF x =- 7859 THEN
            tanh_f := - 2046;
        ELSIF x =- 7858 THEN
            tanh_f := - 2046;
        ELSIF x =- 7857 THEN
            tanh_f := - 2046;
        ELSIF x =- 7856 THEN
            tanh_f := - 2046;
        ELSIF x =- 7855 THEN
            tanh_f := - 2046;
        ELSIF x =- 7854 THEN
            tanh_f := - 2046;
        ELSIF x =- 7853 THEN
            tanh_f := - 2046;
        ELSIF x =- 7852 THEN
            tanh_f := - 2046;
        ELSIF x =- 7851 THEN
            tanh_f := - 2046;
        ELSIF x =- 7850 THEN
            tanh_f := - 2046;
        ELSIF x =- 7849 THEN
            tanh_f := - 2046;
        ELSIF x =- 7848 THEN
            tanh_f := - 2046;
        ELSIF x =- 7847 THEN
            tanh_f := - 2046;
        ELSIF x =- 7846 THEN
            tanh_f := - 2046;
        ELSIF x =- 7845 THEN
            tanh_f := - 2046;
        ELSIF x =- 7844 THEN
            tanh_f := - 2046;
        ELSIF x =- 7843 THEN
            tanh_f := - 2046;
        ELSIF x =- 7842 THEN
            tanh_f := - 2046;
        ELSIF x =- 7841 THEN
            tanh_f := - 2046;
        ELSIF x =- 7840 THEN
            tanh_f := - 2046;
        ELSIF x =- 7839 THEN
            tanh_f := - 2046;
        ELSIF x =- 7838 THEN
            tanh_f := - 2046;
        ELSIF x =- 7837 THEN
            tanh_f := - 2046;
        ELSIF x =- 7836 THEN
            tanh_f := - 2046;
        ELSIF x =- 7835 THEN
            tanh_f := - 2046;
        ELSIF x =- 7834 THEN
            tanh_f := - 2046;
        ELSIF x =- 7833 THEN
            tanh_f := - 2046;
        ELSIF x =- 7832 THEN
            tanh_f := - 2046;
        ELSIF x =- 7831 THEN
            tanh_f := - 2046;
        ELSIF x =- 7830 THEN
            tanh_f := - 2046;
        ELSIF x =- 7829 THEN
            tanh_f := - 2046;
        ELSIF x =- 7828 THEN
            tanh_f := - 2046;
        ELSIF x =- 7827 THEN
            tanh_f := - 2046;
        ELSIF x =- 7826 THEN
            tanh_f := - 2046;
        ELSIF x =- 7825 THEN
            tanh_f := - 2046;
        ELSIF x =- 7824 THEN
            tanh_f := - 2046;
        ELSIF x =- 7823 THEN
            tanh_f := - 2046;
        ELSIF x =- 7822 THEN
            tanh_f := - 2046;
        ELSIF x =- 7821 THEN
            tanh_f := - 2046;
        ELSIF x =- 7820 THEN
            tanh_f := - 2046;
        ELSIF x =- 7819 THEN
            tanh_f := - 2046;
        ELSIF x =- 7818 THEN
            tanh_f := - 2046;
        ELSIF x =- 7817 THEN
            tanh_f := - 2046;
        ELSIF x =- 7816 THEN
            tanh_f := - 2046;
        ELSIF x =- 7815 THEN
            tanh_f := - 2046;
        ELSIF x =- 7814 THEN
            tanh_f := - 2046;
        ELSIF x =- 7813 THEN
            tanh_f := - 2046;
        ELSIF x =- 7812 THEN
            tanh_f := - 2046;
        ELSIF x =- 7811 THEN
            tanh_f := - 2046;
        ELSIF x =- 7810 THEN
            tanh_f := - 2046;
        ELSIF x =- 7809 THEN
            tanh_f := - 2046;
        ELSIF x =- 7808 THEN
            tanh_f := - 2046;
        ELSIF x =- 7807 THEN
            tanh_f := - 2046;
        ELSIF x =- 7806 THEN
            tanh_f := - 2046;
        ELSIF x =- 7805 THEN
            tanh_f := - 2046;
        ELSIF x =- 7804 THEN
            tanh_f := - 2046;
        ELSIF x =- 7803 THEN
            tanh_f := - 2046;
        ELSIF x =- 7802 THEN
            tanh_f := - 2046;
        ELSIF x =- 7801 THEN
            tanh_f := - 2046;
        ELSIF x =- 7800 THEN
            tanh_f := - 2046;
        ELSIF x =- 7799 THEN
            tanh_f := - 2046;
        ELSIF x =- 7798 THEN
            tanh_f := - 2046;
        ELSIF x =- 7797 THEN
            tanh_f := - 2046;
        ELSIF x =- 7796 THEN
            tanh_f := - 2046;
        ELSIF x =- 7795 THEN
            tanh_f := - 2046;
        ELSIF x =- 7794 THEN
            tanh_f := - 2046;
        ELSIF x =- 7793 THEN
            tanh_f := - 2046;
        ELSIF x =- 7792 THEN
            tanh_f := - 2046;
        ELSIF x =- 7791 THEN
            tanh_f := - 2046;
        ELSIF x =- 7790 THEN
            tanh_f := - 2046;
        ELSIF x =- 7789 THEN
            tanh_f := - 2046;
        ELSIF x =- 7788 THEN
            tanh_f := - 2046;
        ELSIF x =- 7787 THEN
            tanh_f := - 2046;
        ELSIF x =- 7786 THEN
            tanh_f := - 2046;
        ELSIF x =- 7785 THEN
            tanh_f := - 2046;
        ELSIF x =- 7784 THEN
            tanh_f := - 2046;
        ELSIF x =- 7783 THEN
            tanh_f := - 2046;
        ELSIF x =- 7782 THEN
            tanh_f := - 2046;
        ELSIF x =- 7781 THEN
            tanh_f := - 2046;
        ELSIF x =- 7780 THEN
            tanh_f := - 2046;
        ELSIF x =- 7779 THEN
            tanh_f := - 2046;
        ELSIF x =- 7778 THEN
            tanh_f := - 2046;
        ELSIF x =- 7777 THEN
            tanh_f := - 2046;
        ELSIF x =- 7776 THEN
            tanh_f := - 2046;
        ELSIF x =- 7775 THEN
            tanh_f := - 2046;
        ELSIF x =- 7774 THEN
            tanh_f := - 2046;
        ELSIF x =- 7773 THEN
            tanh_f := - 2046;
        ELSIF x =- 7772 THEN
            tanh_f := - 2046;
        ELSIF x =- 7771 THEN
            tanh_f := - 2046;
        ELSIF x =- 7770 THEN
            tanh_f := - 2046;
        ELSIF x =- 7769 THEN
            tanh_f := - 2046;
        ELSIF x =- 7768 THEN
            tanh_f := - 2046;
        ELSIF x =- 7767 THEN
            tanh_f := - 2046;
        ELSIF x =- 7766 THEN
            tanh_f := - 2046;
        ELSIF x =- 7765 THEN
            tanh_f := - 2046;
        ELSIF x =- 7764 THEN
            tanh_f := - 2046;
        ELSIF x =- 7763 THEN
            tanh_f := - 2046;
        ELSIF x =- 7762 THEN
            tanh_f := - 2046;
        ELSIF x =- 7761 THEN
            tanh_f := - 2046;
        ELSIF x =- 7760 THEN
            tanh_f := - 2046;
        ELSIF x =- 7759 THEN
            tanh_f := - 2046;
        ELSIF x =- 7758 THEN
            tanh_f := - 2046;
        ELSIF x =- 7757 THEN
            tanh_f := - 2046;
        ELSIF x =- 7756 THEN
            tanh_f := - 2046;
        ELSIF x =- 7755 THEN
            tanh_f := - 2046;
        ELSIF x =- 7754 THEN
            tanh_f := - 2046;
        ELSIF x =- 7753 THEN
            tanh_f := - 2046;
        ELSIF x =- 7752 THEN
            tanh_f := - 2046;
        ELSIF x =- 7751 THEN
            tanh_f := - 2046;
        ELSIF x =- 7750 THEN
            tanh_f := - 2046;
        ELSIF x =- 7749 THEN
            tanh_f := - 2046;
        ELSIF x =- 7748 THEN
            tanh_f := - 2046;
        ELSIF x =- 7747 THEN
            tanh_f := - 2046;
        ELSIF x =- 7746 THEN
            tanh_f := - 2046;
        ELSIF x =- 7745 THEN
            tanh_f := - 2046;
        ELSIF x =- 7744 THEN
            tanh_f := - 2046;
        ELSIF x =- 7743 THEN
            tanh_f := - 2046;
        ELSIF x =- 7742 THEN
            tanh_f := - 2046;
        ELSIF x =- 7741 THEN
            tanh_f := - 2046;
        ELSIF x =- 7740 THEN
            tanh_f := - 2046;
        ELSIF x =- 7739 THEN
            tanh_f := - 2046;
        ELSIF x =- 7738 THEN
            tanh_f := - 2046;
        ELSIF x =- 7737 THEN
            tanh_f := - 2046;
        ELSIF x =- 7736 THEN
            tanh_f := - 2046;
        ELSIF x =- 7735 THEN
            tanh_f := - 2046;
        ELSIF x =- 7734 THEN
            tanh_f := - 2046;
        ELSIF x =- 7733 THEN
            tanh_f := - 2046;
        ELSIF x =- 7732 THEN
            tanh_f := - 2046;
        ELSIF x =- 7731 THEN
            tanh_f := - 2046;
        ELSIF x =- 7730 THEN
            tanh_f := - 2046;
        ELSIF x =- 7729 THEN
            tanh_f := - 2046;
        ELSIF x =- 7728 THEN
            tanh_f := - 2046;
        ELSIF x =- 7727 THEN
            tanh_f := - 2046;
        ELSIF x =- 7726 THEN
            tanh_f := - 2046;
        ELSIF x =- 7725 THEN
            tanh_f := - 2046;
        ELSIF x =- 7724 THEN
            tanh_f := - 2046;
        ELSIF x =- 7723 THEN
            tanh_f := - 2046;
        ELSIF x =- 7722 THEN
            tanh_f := - 2046;
        ELSIF x =- 7721 THEN
            tanh_f := - 2046;
        ELSIF x =- 7720 THEN
            tanh_f := - 2046;
        ELSIF x =- 7719 THEN
            tanh_f := - 2046;
        ELSIF x =- 7718 THEN
            tanh_f := - 2046;
        ELSIF x =- 7717 THEN
            tanh_f := - 2046;
        ELSIF x =- 7716 THEN
            tanh_f := - 2046;
        ELSIF x =- 7715 THEN
            tanh_f := - 2046;
        ELSIF x =- 7714 THEN
            tanh_f := - 2046;
        ELSIF x =- 7713 THEN
            tanh_f := - 2046;
        ELSIF x =- 7712 THEN
            tanh_f := - 2046;
        ELSIF x =- 7711 THEN
            tanh_f := - 2046;
        ELSIF x =- 7710 THEN
            tanh_f := - 2046;
        ELSIF x =- 7709 THEN
            tanh_f := - 2046;
        ELSIF x =- 7708 THEN
            tanh_f := - 2046;
        ELSIF x =- 7707 THEN
            tanh_f := - 2046;
        ELSIF x =- 7706 THEN
            tanh_f := - 2046;
        ELSIF x =- 7705 THEN
            tanh_f := - 2046;
        ELSIF x =- 7704 THEN
            tanh_f := - 2046;
        ELSIF x =- 7703 THEN
            tanh_f := - 2046;
        ELSIF x =- 7702 THEN
            tanh_f := - 2046;
        ELSIF x =- 7701 THEN
            tanh_f := - 2046;
        ELSIF x =- 7700 THEN
            tanh_f := - 2046;
        ELSIF x =- 7699 THEN
            tanh_f := - 2046;
        ELSIF x =- 7698 THEN
            tanh_f := - 2046;
        ELSIF x =- 7697 THEN
            tanh_f := - 2046;
        ELSIF x =- 7696 THEN
            tanh_f := - 2046;
        ELSIF x =- 7695 THEN
            tanh_f := - 2046;
        ELSIF x =- 7694 THEN
            tanh_f := - 2046;
        ELSIF x =- 7693 THEN
            tanh_f := - 2046;
        ELSIF x =- 7692 THEN
            tanh_f := - 2046;
        ELSIF x =- 7691 THEN
            tanh_f := - 2046;
        ELSIF x =- 7690 THEN
            tanh_f := - 2046;
        ELSIF x =- 7689 THEN
            tanh_f := - 2046;
        ELSIF x =- 7688 THEN
            tanh_f := - 2046;
        ELSIF x =- 7687 THEN
            tanh_f := - 2046;
        ELSIF x =- 7686 THEN
            tanh_f := - 2046;
        ELSIF x =- 7685 THEN
            tanh_f := - 2046;
        ELSIF x =- 7684 THEN
            tanh_f := - 2046;
        ELSIF x =- 7683 THEN
            tanh_f := - 2046;
        ELSIF x =- 7682 THEN
            tanh_f := - 2046;
        ELSIF x =- 7681 THEN
            tanh_f := - 2046;
        ELSIF x =- 7680 THEN
            tanh_f := - 2046;
        ELSIF x =- 7679 THEN
            tanh_f := - 2046;
        ELSIF x =- 7678 THEN
            tanh_f := - 2046;
        ELSIF x =- 7677 THEN
            tanh_f := - 2046;
        ELSIF x =- 7676 THEN
            tanh_f := - 2046;
        ELSIF x =- 7675 THEN
            tanh_f := - 2046;
        ELSIF x =- 7674 THEN
            tanh_f := - 2046;
        ELSIF x =- 7673 THEN
            tanh_f := - 2046;
        ELSIF x =- 7672 THEN
            tanh_f := - 2046;
        ELSIF x =- 7671 THEN
            tanh_f := - 2046;
        ELSIF x =- 7670 THEN
            tanh_f := - 2046;
        ELSIF x =- 7669 THEN
            tanh_f := - 2046;
        ELSIF x =- 7668 THEN
            tanh_f := - 2046;
        ELSIF x =- 7667 THEN
            tanh_f := - 2046;
        ELSIF x =- 7666 THEN
            tanh_f := - 2046;
        ELSIF x =- 7665 THEN
            tanh_f := - 2046;
        ELSIF x =- 7664 THEN
            tanh_f := - 2046;
        ELSIF x =- 7663 THEN
            tanh_f := - 2046;
        ELSIF x =- 7662 THEN
            tanh_f := - 2046;
        ELSIF x =- 7661 THEN
            tanh_f := - 2046;
        ELSIF x =- 7660 THEN
            tanh_f := - 2046;
        ELSIF x =- 7659 THEN
            tanh_f := - 2046;
        ELSIF x =- 7658 THEN
            tanh_f := - 2046;
        ELSIF x =- 7657 THEN
            tanh_f := - 2046;
        ELSIF x =- 7656 THEN
            tanh_f := - 2046;
        ELSIF x =- 7655 THEN
            tanh_f := - 2046;
        ELSIF x =- 7654 THEN
            tanh_f := - 2046;
        ELSIF x =- 7653 THEN
            tanh_f := - 2046;
        ELSIF x =- 7652 THEN
            tanh_f := - 2046;
        ELSIF x =- 7651 THEN
            tanh_f := - 2046;
        ELSIF x =- 7650 THEN
            tanh_f := - 2046;
        ELSIF x =- 7649 THEN
            tanh_f := - 2046;
        ELSIF x =- 7648 THEN
            tanh_f := - 2046;
        ELSIF x =- 7647 THEN
            tanh_f := - 2046;
        ELSIF x =- 7646 THEN
            tanh_f := - 2046;
        ELSIF x =- 7645 THEN
            tanh_f := - 2046;
        ELSIF x =- 7644 THEN
            tanh_f := - 2046;
        ELSIF x =- 7643 THEN
            tanh_f := - 2046;
        ELSIF x =- 7642 THEN
            tanh_f := - 2046;
        ELSIF x =- 7641 THEN
            tanh_f := - 2046;
        ELSIF x =- 7640 THEN
            tanh_f := - 2046;
        ELSIF x =- 7639 THEN
            tanh_f := - 2046;
        ELSIF x =- 7638 THEN
            tanh_f := - 2046;
        ELSIF x =- 7637 THEN
            tanh_f := - 2046;
        ELSIF x =- 7636 THEN
            tanh_f := - 2046;
        ELSIF x =- 7635 THEN
            tanh_f := - 2046;
        ELSIF x =- 7634 THEN
            tanh_f := - 2046;
        ELSIF x =- 7633 THEN
            tanh_f := - 2046;
        ELSIF x =- 7632 THEN
            tanh_f := - 2046;
        ELSIF x =- 7631 THEN
            tanh_f := - 2046;
        ELSIF x =- 7630 THEN
            tanh_f := - 2046;
        ELSIF x =- 7629 THEN
            tanh_f := - 2046;
        ELSIF x =- 7628 THEN
            tanh_f := - 2046;
        ELSIF x =- 7627 THEN
            tanh_f := - 2046;
        ELSIF x =- 7626 THEN
            tanh_f := - 2046;
        ELSIF x =- 7625 THEN
            tanh_f := - 2046;
        ELSIF x =- 7624 THEN
            tanh_f := - 2046;
        ELSIF x =- 7623 THEN
            tanh_f := - 2046;
        ELSIF x =- 7622 THEN
            tanh_f := - 2046;
        ELSIF x =- 7621 THEN
            tanh_f := - 2046;
        ELSIF x =- 7620 THEN
            tanh_f := - 2046;
        ELSIF x =- 7619 THEN
            tanh_f := - 2046;
        ELSIF x =- 7618 THEN
            tanh_f := - 2046;
        ELSIF x =- 7617 THEN
            tanh_f := - 2046;
        ELSIF x =- 7616 THEN
            tanh_f := - 2046;
        ELSIF x =- 7615 THEN
            tanh_f := - 2046;
        ELSIF x =- 7614 THEN
            tanh_f := - 2046;
        ELSIF x =- 7613 THEN
            tanh_f := - 2046;
        ELSIF x =- 7612 THEN
            tanh_f := - 2046;
        ELSIF x =- 7611 THEN
            tanh_f := - 2046;
        ELSIF x =- 7610 THEN
            tanh_f := - 2046;
        ELSIF x =- 7609 THEN
            tanh_f := - 2046;
        ELSIF x =- 7608 THEN
            tanh_f := - 2046;
        ELSIF x =- 7607 THEN
            tanh_f := - 2046;
        ELSIF x =- 7606 THEN
            tanh_f := - 2046;
        ELSIF x =- 7605 THEN
            tanh_f := - 2046;
        ELSIF x =- 7604 THEN
            tanh_f := - 2046;
        ELSIF x =- 7603 THEN
            tanh_f := - 2046;
        ELSIF x =- 7602 THEN
            tanh_f := - 2046;
        ELSIF x =- 7601 THEN
            tanh_f := - 2046;
        ELSIF x =- 7600 THEN
            tanh_f := - 2046;
        ELSIF x =- 7599 THEN
            tanh_f := - 2046;
        ELSIF x =- 7598 THEN
            tanh_f := - 2046;
        ELSIF x =- 7597 THEN
            tanh_f := - 2046;
        ELSIF x =- 7596 THEN
            tanh_f := - 2046;
        ELSIF x =- 7595 THEN
            tanh_f := - 2046;
        ELSIF x =- 7594 THEN
            tanh_f := - 2046;
        ELSIF x =- 7593 THEN
            tanh_f := - 2046;
        ELSIF x =- 7592 THEN
            tanh_f := - 2046;
        ELSIF x =- 7591 THEN
            tanh_f := - 2046;
        ELSIF x =- 7590 THEN
            tanh_f := - 2046;
        ELSIF x =- 7589 THEN
            tanh_f := - 2046;
        ELSIF x =- 7588 THEN
            tanh_f := - 2046;
        ELSIF x =- 7587 THEN
            tanh_f := - 2046;
        ELSIF x =- 7586 THEN
            tanh_f := - 2046;
        ELSIF x =- 7585 THEN
            tanh_f := - 2046;
        ELSIF x =- 7584 THEN
            tanh_f := - 2046;
        ELSIF x =- 7583 THEN
            tanh_f := - 2046;
        ELSIF x =- 7582 THEN
            tanh_f := - 2046;
        ELSIF x =- 7581 THEN
            tanh_f := - 2046;
        ELSIF x =- 7580 THEN
            tanh_f := - 2046;
        ELSIF x =- 7579 THEN
            tanh_f := - 2046;
        ELSIF x =- 7578 THEN
            tanh_f := - 2046;
        ELSIF x =- 7577 THEN
            tanh_f := - 2046;
        ELSIF x =- 7576 THEN
            tanh_f := - 2046;
        ELSIF x =- 7575 THEN
            tanh_f := - 2046;
        ELSIF x =- 7574 THEN
            tanh_f := - 2046;
        ELSIF x =- 7573 THEN
            tanh_f := - 2046;
        ELSIF x =- 7572 THEN
            tanh_f := - 2046;
        ELSIF x =- 7571 THEN
            tanh_f := - 2046;
        ELSIF x =- 7570 THEN
            tanh_f := - 2046;
        ELSIF x =- 7569 THEN
            tanh_f := - 2046;
        ELSIF x =- 7568 THEN
            tanh_f := - 2046;
        ELSIF x =- 7567 THEN
            tanh_f := - 2046;
        ELSIF x =- 7566 THEN
            tanh_f := - 2046;
        ELSIF x =- 7565 THEN
            tanh_f := - 2046;
        ELSIF x =- 7564 THEN
            tanh_f := - 2046;
        ELSIF x =- 7563 THEN
            tanh_f := - 2046;
        ELSIF x =- 7562 THEN
            tanh_f := - 2046;
        ELSIF x =- 7561 THEN
            tanh_f := - 2046;
        ELSIF x =- 7560 THEN
            tanh_f := - 2046;
        ELSIF x =- 7559 THEN
            tanh_f := - 2046;
        ELSIF x =- 7558 THEN
            tanh_f := - 2046;
        ELSIF x =- 7557 THEN
            tanh_f := - 2046;
        ELSIF x =- 7556 THEN
            tanh_f := - 2046;
        ELSIF x =- 7555 THEN
            tanh_f := - 2046;
        ELSIF x =- 7554 THEN
            tanh_f := - 2046;
        ELSIF x =- 7553 THEN
            tanh_f := - 2046;
        ELSIF x =- 7552 THEN
            tanh_f := - 2046;
        ELSIF x =- 7551 THEN
            tanh_f := - 2046;
        ELSIF x =- 7550 THEN
            tanh_f := - 2046;
        ELSIF x =- 7549 THEN
            tanh_f := - 2046;
        ELSIF x =- 7548 THEN
            tanh_f := - 2046;
        ELSIF x =- 7547 THEN
            tanh_f := - 2046;
        ELSIF x =- 7546 THEN
            tanh_f := - 2046;
        ELSIF x =- 7545 THEN
            tanh_f := - 2046;
        ELSIF x =- 7544 THEN
            tanh_f := - 2046;
        ELSIF x =- 7543 THEN
            tanh_f := - 2046;
        ELSIF x =- 7542 THEN
            tanh_f := - 2046;
        ELSIF x =- 7541 THEN
            tanh_f := - 2046;
        ELSIF x =- 7540 THEN
            tanh_f := - 2046;
        ELSIF x =- 7539 THEN
            tanh_f := - 2046;
        ELSIF x =- 7538 THEN
            tanh_f := - 2046;
        ELSIF x =- 7537 THEN
            tanh_f := - 2046;
        ELSIF x =- 7536 THEN
            tanh_f := - 2046;
        ELSIF x =- 7535 THEN
            tanh_f := - 2046;
        ELSIF x =- 7534 THEN
            tanh_f := - 2046;
        ELSIF x =- 7533 THEN
            tanh_f := - 2046;
        ELSIF x =- 7532 THEN
            tanh_f := - 2046;
        ELSIF x =- 7531 THEN
            tanh_f := - 2046;
        ELSIF x =- 7530 THEN
            tanh_f := - 2046;
        ELSIF x =- 7529 THEN
            tanh_f := - 2046;
        ELSIF x =- 7528 THEN
            tanh_f := - 2046;
        ELSIF x =- 7527 THEN
            tanh_f := - 2046;
        ELSIF x =- 7526 THEN
            tanh_f := - 2046;
        ELSIF x =- 7525 THEN
            tanh_f := - 2046;
        ELSIF x =- 7524 THEN
            tanh_f := - 2046;
        ELSIF x =- 7523 THEN
            tanh_f := - 2046;
        ELSIF x =- 7522 THEN
            tanh_f := - 2046;
        ELSIF x =- 7521 THEN
            tanh_f := - 2046;
        ELSIF x =- 7520 THEN
            tanh_f := - 2046;
        ELSIF x =- 7519 THEN
            tanh_f := - 2046;
        ELSIF x =- 7518 THEN
            tanh_f := - 2046;
        ELSIF x =- 7517 THEN
            tanh_f := - 2046;
        ELSIF x =- 7516 THEN
            tanh_f := - 2046;
        ELSIF x =- 7515 THEN
            tanh_f := - 2046;
        ELSIF x =- 7514 THEN
            tanh_f := - 2046;
        ELSIF x =- 7513 THEN
            tanh_f := - 2046;
        ELSIF x =- 7512 THEN
            tanh_f := - 2046;
        ELSIF x =- 7511 THEN
            tanh_f := - 2046;
        ELSIF x =- 7510 THEN
            tanh_f := - 2046;
        ELSIF x =- 7509 THEN
            tanh_f := - 2046;
        ELSIF x =- 7508 THEN
            tanh_f := - 2046;
        ELSIF x =- 7507 THEN
            tanh_f := - 2046;
        ELSIF x =- 7506 THEN
            tanh_f := - 2046;
        ELSIF x =- 7505 THEN
            tanh_f := - 2046;
        ELSIF x =- 7504 THEN
            tanh_f := - 2046;
        ELSIF x =- 7503 THEN
            tanh_f := - 2046;
        ELSIF x =- 7502 THEN
            tanh_f := - 2046;
        ELSIF x =- 7501 THEN
            tanh_f := - 2046;
        ELSIF x =- 7500 THEN
            tanh_f := - 2046;
        ELSIF x =- 7499 THEN
            tanh_f := - 2046;
        ELSIF x =- 7498 THEN
            tanh_f := - 2046;
        ELSIF x =- 7497 THEN
            tanh_f := - 2046;
        ELSIF x =- 7496 THEN
            tanh_f := - 2046;
        ELSIF x =- 7495 THEN
            tanh_f := - 2046;
        ELSIF x =- 7494 THEN
            tanh_f := - 2046;
        ELSIF x =- 7493 THEN
            tanh_f := - 2046;
        ELSIF x =- 7492 THEN
            tanh_f := - 2046;
        ELSIF x =- 7491 THEN
            tanh_f := - 2046;
        ELSIF x =- 7490 THEN
            tanh_f := - 2046;
        ELSIF x =- 7489 THEN
            tanh_f := - 2046;
        ELSIF x =- 7488 THEN
            tanh_f := - 2046;
        ELSIF x =- 7487 THEN
            tanh_f := - 2046;
        ELSIF x =- 7486 THEN
            tanh_f := - 2046;
        ELSIF x =- 7485 THEN
            tanh_f := - 2046;
        ELSIF x =- 7484 THEN
            tanh_f := - 2046;
        ELSIF x =- 7483 THEN
            tanh_f := - 2046;
        ELSIF x =- 7482 THEN
            tanh_f := - 2046;
        ELSIF x =- 7481 THEN
            tanh_f := - 2046;
        ELSIF x =- 7480 THEN
            tanh_f := - 2046;
        ELSIF x =- 7479 THEN
            tanh_f := - 2046;
        ELSIF x =- 7478 THEN
            tanh_f := - 2046;
        ELSIF x =- 7477 THEN
            tanh_f := - 2046;
        ELSIF x =- 7476 THEN
            tanh_f := - 2046;
        ELSIF x =- 7475 THEN
            tanh_f := - 2046;
        ELSIF x =- 7474 THEN
            tanh_f := - 2046;
        ELSIF x =- 7473 THEN
            tanh_f := - 2046;
        ELSIF x =- 7472 THEN
            tanh_f := - 2046;
        ELSIF x =- 7471 THEN
            tanh_f := - 2046;
        ELSIF x =- 7470 THEN
            tanh_f := - 2046;
        ELSIF x =- 7469 THEN
            tanh_f := - 2046;
        ELSIF x =- 7468 THEN
            tanh_f := - 2046;
        ELSIF x =- 7467 THEN
            tanh_f := - 2046;
        ELSIF x =- 7466 THEN
            tanh_f := - 2046;
        ELSIF x =- 7465 THEN
            tanh_f := - 2046;
        ELSIF x =- 7464 THEN
            tanh_f := - 2046;
        ELSIF x =- 7463 THEN
            tanh_f := - 2046;
        ELSIF x =- 7462 THEN
            tanh_f := - 2046;
        ELSIF x =- 7461 THEN
            tanh_f := - 2046;
        ELSIF x =- 7460 THEN
            tanh_f := - 2046;
        ELSIF x =- 7459 THEN
            tanh_f := - 2046;
        ELSIF x =- 7458 THEN
            tanh_f := - 2046;
        ELSIF x =- 7457 THEN
            tanh_f := - 2046;
        ELSIF x =- 7456 THEN
            tanh_f := - 2046;
        ELSIF x =- 7455 THEN
            tanh_f := - 2046;
        ELSIF x =- 7454 THEN
            tanh_f := - 2046;
        ELSIF x =- 7453 THEN
            tanh_f := - 2046;
        ELSIF x =- 7452 THEN
            tanh_f := - 2046;
        ELSIF x =- 7451 THEN
            tanh_f := - 2046;
        ELSIF x =- 7450 THEN
            tanh_f := - 2046;
        ELSIF x =- 7449 THEN
            tanh_f := - 2046;
        ELSIF x =- 7448 THEN
            tanh_f := - 2046;
        ELSIF x =- 7447 THEN
            tanh_f := - 2046;
        ELSIF x =- 7446 THEN
            tanh_f := - 2046;
        ELSIF x =- 7445 THEN
            tanh_f := - 2046;
        ELSIF x =- 7444 THEN
            tanh_f := - 2046;
        ELSIF x =- 7443 THEN
            tanh_f := - 2046;
        ELSIF x =- 7442 THEN
            tanh_f := - 2046;
        ELSIF x =- 7441 THEN
            tanh_f := - 2046;
        ELSIF x =- 7440 THEN
            tanh_f := - 2046;
        ELSIF x =- 7439 THEN
            tanh_f := - 2046;
        ELSIF x =- 7438 THEN
            tanh_f := - 2046;
        ELSIF x =- 7437 THEN
            tanh_f := - 2046;
        ELSIF x =- 7436 THEN
            tanh_f := - 2046;
        ELSIF x =- 7435 THEN
            tanh_f := - 2046;
        ELSIF x =- 7434 THEN
            tanh_f := - 2046;
        ELSIF x =- 7433 THEN
            tanh_f := - 2046;
        ELSIF x =- 7432 THEN
            tanh_f := - 2046;
        ELSIF x =- 7431 THEN
            tanh_f := - 2046;
        ELSIF x =- 7430 THEN
            tanh_f := - 2046;
        ELSIF x =- 7429 THEN
            tanh_f := - 2046;
        ELSIF x =- 7428 THEN
            tanh_f := - 2046;
        ELSIF x =- 7427 THEN
            tanh_f := - 2046;
        ELSIF x =- 7426 THEN
            tanh_f := - 2046;
        ELSIF x =- 7425 THEN
            tanh_f := - 2046;
        ELSIF x =- 7424 THEN
            tanh_f := - 2046;
        ELSIF x =- 7423 THEN
            tanh_f := - 2044;
        ELSIF x =- 7422 THEN
            tanh_f := - 2044;
        ELSIF x =- 7421 THEN
            tanh_f := - 2044;
        ELSIF x =- 7420 THEN
            tanh_f := - 2044;
        ELSIF x =- 7419 THEN
            tanh_f := - 2044;
        ELSIF x =- 7418 THEN
            tanh_f := - 2044;
        ELSIF x =- 7417 THEN
            tanh_f := - 2044;
        ELSIF x =- 7416 THEN
            tanh_f := - 2044;
        ELSIF x =- 7415 THEN
            tanh_f := - 2044;
        ELSIF x =- 7414 THEN
            tanh_f := - 2044;
        ELSIF x =- 7413 THEN
            tanh_f := - 2044;
        ELSIF x =- 7412 THEN
            tanh_f := - 2044;
        ELSIF x =- 7411 THEN
            tanh_f := - 2044;
        ELSIF x =- 7410 THEN
            tanh_f := - 2044;
        ELSIF x =- 7409 THEN
            tanh_f := - 2044;
        ELSIF x =- 7408 THEN
            tanh_f := - 2044;
        ELSIF x =- 7407 THEN
            tanh_f := - 2044;
        ELSIF x =- 7406 THEN
            tanh_f := - 2044;
        ELSIF x =- 7405 THEN
            tanh_f := - 2044;
        ELSIF x =- 7404 THEN
            tanh_f := - 2044;
        ELSIF x =- 7403 THEN
            tanh_f := - 2044;
        ELSIF x =- 7402 THEN
            tanh_f := - 2044;
        ELSIF x =- 7401 THEN
            tanh_f := - 2044;
        ELSIF x =- 7400 THEN
            tanh_f := - 2044;
        ELSIF x =- 7399 THEN
            tanh_f := - 2044;
        ELSIF x =- 7398 THEN
            tanh_f := - 2044;
        ELSIF x =- 7397 THEN
            tanh_f := - 2044;
        ELSIF x =- 7396 THEN
            tanh_f := - 2044;
        ELSIF x =- 7395 THEN
            tanh_f := - 2044;
        ELSIF x =- 7394 THEN
            tanh_f := - 2044;
        ELSIF x =- 7393 THEN
            tanh_f := - 2044;
        ELSIF x =- 7392 THEN
            tanh_f := - 2044;
        ELSIF x =- 7391 THEN
            tanh_f := - 2044;
        ELSIF x =- 7390 THEN
            tanh_f := - 2044;
        ELSIF x =- 7389 THEN
            tanh_f := - 2044;
        ELSIF x =- 7388 THEN
            tanh_f := - 2044;
        ELSIF x =- 7387 THEN
            tanh_f := - 2044;
        ELSIF x =- 7386 THEN
            tanh_f := - 2044;
        ELSIF x =- 7385 THEN
            tanh_f := - 2044;
        ELSIF x =- 7384 THEN
            tanh_f := - 2044;
        ELSIF x =- 7383 THEN
            tanh_f := - 2044;
        ELSIF x =- 7382 THEN
            tanh_f := - 2044;
        ELSIF x =- 7381 THEN
            tanh_f := - 2044;
        ELSIF x =- 7380 THEN
            tanh_f := - 2044;
        ELSIF x =- 7379 THEN
            tanh_f := - 2044;
        ELSIF x =- 7378 THEN
            tanh_f := - 2044;
        ELSIF x =- 7377 THEN
            tanh_f := - 2044;
        ELSIF x =- 7376 THEN
            tanh_f := - 2044;
        ELSIF x =- 7375 THEN
            tanh_f := - 2044;
        ELSIF x =- 7374 THEN
            tanh_f := - 2044;
        ELSIF x =- 7373 THEN
            tanh_f := - 2044;
        ELSIF x =- 7372 THEN
            tanh_f := - 2044;
        ELSIF x =- 7371 THEN
            tanh_f := - 2044;
        ELSIF x =- 7370 THEN
            tanh_f := - 2044;
        ELSIF x =- 7369 THEN
            tanh_f := - 2044;
        ELSIF x =- 7368 THEN
            tanh_f := - 2044;
        ELSIF x =- 7367 THEN
            tanh_f := - 2044;
        ELSIF x =- 7366 THEN
            tanh_f := - 2044;
        ELSIF x =- 7365 THEN
            tanh_f := - 2044;
        ELSIF x =- 7364 THEN
            tanh_f := - 2044;
        ELSIF x =- 7363 THEN
            tanh_f := - 2044;
        ELSIF x =- 7362 THEN
            tanh_f := - 2044;
        ELSIF x =- 7361 THEN
            tanh_f := - 2044;
        ELSIF x =- 7360 THEN
            tanh_f := - 2044;
        ELSIF x =- 7359 THEN
            tanh_f := - 2044;
        ELSIF x =- 7358 THEN
            tanh_f := - 2044;
        ELSIF x =- 7357 THEN
            tanh_f := - 2044;
        ELSIF x =- 7356 THEN
            tanh_f := - 2044;
        ELSIF x =- 7355 THEN
            tanh_f := - 2044;
        ELSIF x =- 7354 THEN
            tanh_f := - 2044;
        ELSIF x =- 7353 THEN
            tanh_f := - 2044;
        ELSIF x =- 7352 THEN
            tanh_f := - 2044;
        ELSIF x =- 7351 THEN
            tanh_f := - 2044;
        ELSIF x =- 7350 THEN
            tanh_f := - 2044;
        ELSIF x =- 7349 THEN
            tanh_f := - 2044;
        ELSIF x =- 7348 THEN
            tanh_f := - 2044;
        ELSIF x =- 7347 THEN
            tanh_f := - 2044;
        ELSIF x =- 7346 THEN
            tanh_f := - 2044;
        ELSIF x =- 7345 THEN
            tanh_f := - 2044;
        ELSIF x =- 7344 THEN
            tanh_f := - 2044;
        ELSIF x =- 7343 THEN
            tanh_f := - 2044;
        ELSIF x =- 7342 THEN
            tanh_f := - 2044;
        ELSIF x =- 7341 THEN
            tanh_f := - 2044;
        ELSIF x =- 7340 THEN
            tanh_f := - 2044;
        ELSIF x =- 7339 THEN
            tanh_f := - 2044;
        ELSIF x =- 7338 THEN
            tanh_f := - 2044;
        ELSIF x =- 7337 THEN
            tanh_f := - 2044;
        ELSIF x =- 7336 THEN
            tanh_f := - 2044;
        ELSIF x =- 7335 THEN
            tanh_f := - 2044;
        ELSIF x =- 7334 THEN
            tanh_f := - 2044;
        ELSIF x =- 7333 THEN
            tanh_f := - 2044;
        ELSIF x =- 7332 THEN
            tanh_f := - 2044;
        ELSIF x =- 7331 THEN
            tanh_f := - 2044;
        ELSIF x =- 7330 THEN
            tanh_f := - 2044;
        ELSIF x =- 7329 THEN
            tanh_f := - 2044;
        ELSIF x =- 7328 THEN
            tanh_f := - 2044;
        ELSIF x =- 7327 THEN
            tanh_f := - 2044;
        ELSIF x =- 7326 THEN
            tanh_f := - 2044;
        ELSIF x =- 7325 THEN
            tanh_f := - 2044;
        ELSIF x =- 7324 THEN
            tanh_f := - 2044;
        ELSIF x =- 7323 THEN
            tanh_f := - 2044;
        ELSIF x =- 7322 THEN
            tanh_f := - 2044;
        ELSIF x =- 7321 THEN
            tanh_f := - 2044;
        ELSIF x =- 7320 THEN
            tanh_f := - 2044;
        ELSIF x =- 7319 THEN
            tanh_f := - 2044;
        ELSIF x =- 7318 THEN
            tanh_f := - 2044;
        ELSIF x =- 7317 THEN
            tanh_f := - 2044;
        ELSIF x =- 7316 THEN
            tanh_f := - 2044;
        ELSIF x =- 7315 THEN
            tanh_f := - 2044;
        ELSIF x =- 7314 THEN
            tanh_f := - 2044;
        ELSIF x =- 7313 THEN
            tanh_f := - 2044;
        ELSIF x =- 7312 THEN
            tanh_f := - 2044;
        ELSIF x =- 7311 THEN
            tanh_f := - 2044;
        ELSIF x =- 7310 THEN
            tanh_f := - 2044;
        ELSIF x =- 7309 THEN
            tanh_f := - 2044;
        ELSIF x =- 7308 THEN
            tanh_f := - 2044;
        ELSIF x =- 7307 THEN
            tanh_f := - 2044;
        ELSIF x =- 7306 THEN
            tanh_f := - 2044;
        ELSIF x =- 7305 THEN
            tanh_f := - 2044;
        ELSIF x =- 7304 THEN
            tanh_f := - 2044;
        ELSIF x =- 7303 THEN
            tanh_f := - 2044;
        ELSIF x =- 7302 THEN
            tanh_f := - 2044;
        ELSIF x =- 7301 THEN
            tanh_f := - 2044;
        ELSIF x =- 7300 THEN
            tanh_f := - 2044;
        ELSIF x =- 7299 THEN
            tanh_f := - 2044;
        ELSIF x =- 7298 THEN
            tanh_f := - 2044;
        ELSIF x =- 7297 THEN
            tanh_f := - 2044;
        ELSIF x =- 7296 THEN
            tanh_f := - 2044;
        ELSIF x =- 7295 THEN
            tanh_f := - 2044;
        ELSIF x =- 7294 THEN
            tanh_f := - 2044;
        ELSIF x =- 7293 THEN
            tanh_f := - 2044;
        ELSIF x =- 7292 THEN
            tanh_f := - 2044;
        ELSIF x =- 7291 THEN
            tanh_f := - 2044;
        ELSIF x =- 7290 THEN
            tanh_f := - 2044;
        ELSIF x =- 7289 THEN
            tanh_f := - 2044;
        ELSIF x =- 7288 THEN
            tanh_f := - 2044;
        ELSIF x =- 7287 THEN
            tanh_f := - 2044;
        ELSIF x =- 7286 THEN
            tanh_f := - 2044;
        ELSIF x =- 7285 THEN
            tanh_f := - 2044;
        ELSIF x =- 7284 THEN
            tanh_f := - 2044;
        ELSIF x =- 7283 THEN
            tanh_f := - 2044;
        ELSIF x =- 7282 THEN
            tanh_f := - 2044;
        ELSIF x =- 7281 THEN
            tanh_f := - 2044;
        ELSIF x =- 7280 THEN
            tanh_f := - 2044;
        ELSIF x =- 7279 THEN
            tanh_f := - 2044;
        ELSIF x =- 7278 THEN
            tanh_f := - 2044;
        ELSIF x =- 7277 THEN
            tanh_f := - 2044;
        ELSIF x =- 7276 THEN
            tanh_f := - 2044;
        ELSIF x =- 7275 THEN
            tanh_f := - 2044;
        ELSIF x =- 7274 THEN
            tanh_f := - 2044;
        ELSIF x =- 7273 THEN
            tanh_f := - 2044;
        ELSIF x =- 7272 THEN
            tanh_f := - 2044;
        ELSIF x =- 7271 THEN
            tanh_f := - 2044;
        ELSIF x =- 7270 THEN
            tanh_f := - 2044;
        ELSIF x =- 7269 THEN
            tanh_f := - 2044;
        ELSIF x =- 7268 THEN
            tanh_f := - 2044;
        ELSIF x =- 7267 THEN
            tanh_f := - 2044;
        ELSIF x =- 7266 THEN
            tanh_f := - 2044;
        ELSIF x =- 7265 THEN
            tanh_f := - 2044;
        ELSIF x =- 7264 THEN
            tanh_f := - 2044;
        ELSIF x =- 7263 THEN
            tanh_f := - 2044;
        ELSIF x =- 7262 THEN
            tanh_f := - 2044;
        ELSIF x =- 7261 THEN
            tanh_f := - 2044;
        ELSIF x =- 7260 THEN
            tanh_f := - 2044;
        ELSIF x =- 7259 THEN
            tanh_f := - 2044;
        ELSIF x =- 7258 THEN
            tanh_f := - 2044;
        ELSIF x =- 7257 THEN
            tanh_f := - 2044;
        ELSIF x =- 7256 THEN
            tanh_f := - 2044;
        ELSIF x =- 7255 THEN
            tanh_f := - 2044;
        ELSIF x =- 7254 THEN
            tanh_f := - 2044;
        ELSIF x =- 7253 THEN
            tanh_f := - 2044;
        ELSIF x =- 7252 THEN
            tanh_f := - 2044;
        ELSIF x =- 7251 THEN
            tanh_f := - 2044;
        ELSIF x =- 7250 THEN
            tanh_f := - 2044;
        ELSIF x =- 7249 THEN
            tanh_f := - 2044;
        ELSIF x =- 7248 THEN
            tanh_f := - 2044;
        ELSIF x =- 7247 THEN
            tanh_f := - 2044;
        ELSIF x =- 7246 THEN
            tanh_f := - 2044;
        ELSIF x =- 7245 THEN
            tanh_f := - 2044;
        ELSIF x =- 7244 THEN
            tanh_f := - 2044;
        ELSIF x =- 7243 THEN
            tanh_f := - 2044;
        ELSIF x =- 7242 THEN
            tanh_f := - 2044;
        ELSIF x =- 7241 THEN
            tanh_f := - 2044;
        ELSIF x =- 7240 THEN
            tanh_f := - 2044;
        ELSIF x =- 7239 THEN
            tanh_f := - 2044;
        ELSIF x =- 7238 THEN
            tanh_f := - 2044;
        ELSIF x =- 7237 THEN
            tanh_f := - 2044;
        ELSIF x =- 7236 THEN
            tanh_f := - 2044;
        ELSIF x =- 7235 THEN
            tanh_f := - 2044;
        ELSIF x =- 7234 THEN
            tanh_f := - 2044;
        ELSIF x =- 7233 THEN
            tanh_f := - 2044;
        ELSIF x =- 7232 THEN
            tanh_f := - 2044;
        ELSIF x =- 7231 THEN
            tanh_f := - 2044;
        ELSIF x =- 7230 THEN
            tanh_f := - 2044;
        ELSIF x =- 7229 THEN
            tanh_f := - 2044;
        ELSIF x =- 7228 THEN
            tanh_f := - 2044;
        ELSIF x =- 7227 THEN
            tanh_f := - 2044;
        ELSIF x =- 7226 THEN
            tanh_f := - 2044;
        ELSIF x =- 7225 THEN
            tanh_f := - 2044;
        ELSIF x =- 7224 THEN
            tanh_f := - 2044;
        ELSIF x =- 7223 THEN
            tanh_f := - 2044;
        ELSIF x =- 7222 THEN
            tanh_f := - 2044;
        ELSIF x =- 7221 THEN
            tanh_f := - 2044;
        ELSIF x =- 7220 THEN
            tanh_f := - 2044;
        ELSIF x =- 7219 THEN
            tanh_f := - 2044;
        ELSIF x =- 7218 THEN
            tanh_f := - 2044;
        ELSIF x =- 7217 THEN
            tanh_f := - 2044;
        ELSIF x =- 7216 THEN
            tanh_f := - 2044;
        ELSIF x =- 7215 THEN
            tanh_f := - 2044;
        ELSIF x =- 7214 THEN
            tanh_f := - 2044;
        ELSIF x =- 7213 THEN
            tanh_f := - 2044;
        ELSIF x =- 7212 THEN
            tanh_f := - 2044;
        ELSIF x =- 7211 THEN
            tanh_f := - 2044;
        ELSIF x =- 7210 THEN
            tanh_f := - 2044;
        ELSIF x =- 7209 THEN
            tanh_f := - 2044;
        ELSIF x =- 7208 THEN
            tanh_f := - 2044;
        ELSIF x =- 7207 THEN
            tanh_f := - 2044;
        ELSIF x =- 7206 THEN
            tanh_f := - 2044;
        ELSIF x =- 7205 THEN
            tanh_f := - 2044;
        ELSIF x =- 7204 THEN
            tanh_f := - 2044;
        ELSIF x =- 7203 THEN
            tanh_f := - 2044;
        ELSIF x =- 7202 THEN
            tanh_f := - 2044;
        ELSIF x =- 7201 THEN
            tanh_f := - 2044;
        ELSIF x =- 7200 THEN
            tanh_f := - 2044;
        ELSIF x =- 7199 THEN
            tanh_f := - 2044;
        ELSIF x =- 7198 THEN
            tanh_f := - 2044;
        ELSIF x =- 7197 THEN
            tanh_f := - 2044;
        ELSIF x =- 7196 THEN
            tanh_f := - 2044;
        ELSIF x =- 7195 THEN
            tanh_f := - 2044;
        ELSIF x =- 7194 THEN
            tanh_f := - 2044;
        ELSIF x =- 7193 THEN
            tanh_f := - 2044;
        ELSIF x =- 7192 THEN
            tanh_f := - 2044;
        ELSIF x =- 7191 THEN
            tanh_f := - 2044;
        ELSIF x =- 7190 THEN
            tanh_f := - 2044;
        ELSIF x =- 7189 THEN
            tanh_f := - 2044;
        ELSIF x =- 7188 THEN
            tanh_f := - 2044;
        ELSIF x =- 7187 THEN
            tanh_f := - 2044;
        ELSIF x =- 7186 THEN
            tanh_f := - 2044;
        ELSIF x =- 7185 THEN
            tanh_f := - 2044;
        ELSIF x =- 7184 THEN
            tanh_f := - 2044;
        ELSIF x =- 7183 THEN
            tanh_f := - 2044;
        ELSIF x =- 7182 THEN
            tanh_f := - 2044;
        ELSIF x =- 7181 THEN
            tanh_f := - 2044;
        ELSIF x =- 7180 THEN
            tanh_f := - 2044;
        ELSIF x =- 7179 THEN
            tanh_f := - 2044;
        ELSIF x =- 7178 THEN
            tanh_f := - 2044;
        ELSIF x =- 7177 THEN
            tanh_f := - 2044;
        ELSIF x =- 7176 THEN
            tanh_f := - 2044;
        ELSIF x =- 7175 THEN
            tanh_f := - 2044;
        ELSIF x =- 7174 THEN
            tanh_f := - 2044;
        ELSIF x =- 7173 THEN
            tanh_f := - 2044;
        ELSIF x =- 7172 THEN
            tanh_f := - 2044;
        ELSIF x =- 7171 THEN
            tanh_f := - 2044;
        ELSIF x =- 7170 THEN
            tanh_f := - 2044;
        ELSIF x =- 7169 THEN
            tanh_f := - 2044;
        ELSIF x =- 7168 THEN
            tanh_f := - 2044;
        ELSIF x =- 7167 THEN
            tanh_f := - 2044;
        ELSIF x =- 7166 THEN
            tanh_f := - 2044;
        ELSIF x =- 7165 THEN
            tanh_f := - 2044;
        ELSIF x =- 7164 THEN
            tanh_f := - 2044;
        ELSIF x =- 7163 THEN
            tanh_f := - 2044;
        ELSIF x =- 7162 THEN
            tanh_f := - 2044;
        ELSIF x =- 7161 THEN
            tanh_f := - 2044;
        ELSIF x =- 7160 THEN
            tanh_f := - 2044;
        ELSIF x =- 7159 THEN
            tanh_f := - 2044;
        ELSIF x =- 7158 THEN
            tanh_f := - 2044;
        ELSIF x =- 7157 THEN
            tanh_f := - 2044;
        ELSIF x =- 7156 THEN
            tanh_f := - 2044;
        ELSIF x =- 7155 THEN
            tanh_f := - 2044;
        ELSIF x =- 7154 THEN
            tanh_f := - 2044;
        ELSIF x =- 7153 THEN
            tanh_f := - 2044;
        ELSIF x =- 7152 THEN
            tanh_f := - 2044;
        ELSIF x =- 7151 THEN
            tanh_f := - 2044;
        ELSIF x =- 7150 THEN
            tanh_f := - 2044;
        ELSIF x =- 7149 THEN
            tanh_f := - 2044;
        ELSIF x =- 7148 THEN
            tanh_f := - 2044;
        ELSIF x =- 7147 THEN
            tanh_f := - 2044;
        ELSIF x =- 7146 THEN
            tanh_f := - 2044;
        ELSIF x =- 7145 THEN
            tanh_f := - 2044;
        ELSIF x =- 7144 THEN
            tanh_f := - 2044;
        ELSIF x =- 7143 THEN
            tanh_f := - 2044;
        ELSIF x =- 7142 THEN
            tanh_f := - 2044;
        ELSIF x =- 7141 THEN
            tanh_f := - 2044;
        ELSIF x =- 7140 THEN
            tanh_f := - 2044;
        ELSIF x =- 7139 THEN
            tanh_f := - 2044;
        ELSIF x =- 7138 THEN
            tanh_f := - 2044;
        ELSIF x =- 7137 THEN
            tanh_f := - 2044;
        ELSIF x =- 7136 THEN
            tanh_f := - 2044;
        ELSIF x =- 7135 THEN
            tanh_f := - 2044;
        ELSIF x =- 7134 THEN
            tanh_f := - 2044;
        ELSIF x =- 7133 THEN
            tanh_f := - 2044;
        ELSIF x =- 7132 THEN
            tanh_f := - 2044;
        ELSIF x =- 7131 THEN
            tanh_f := - 2044;
        ELSIF x =- 7130 THEN
            tanh_f := - 2044;
        ELSIF x =- 7129 THEN
            tanh_f := - 2044;
        ELSIF x =- 7128 THEN
            tanh_f := - 2044;
        ELSIF x =- 7127 THEN
            tanh_f := - 2044;
        ELSIF x =- 7126 THEN
            tanh_f := - 2044;
        ELSIF x =- 7125 THEN
            tanh_f := - 2044;
        ELSIF x =- 7124 THEN
            tanh_f := - 2044;
        ELSIF x =- 7123 THEN
            tanh_f := - 2044;
        ELSIF x =- 7122 THEN
            tanh_f := - 2044;
        ELSIF x =- 7121 THEN
            tanh_f := - 2044;
        ELSIF x =- 7120 THEN
            tanh_f := - 2044;
        ELSIF x =- 7119 THEN
            tanh_f := - 2044;
        ELSIF x =- 7118 THEN
            tanh_f := - 2044;
        ELSIF x =- 7117 THEN
            tanh_f := - 2044;
        ELSIF x =- 7116 THEN
            tanh_f := - 2044;
        ELSIF x =- 7115 THEN
            tanh_f := - 2044;
        ELSIF x =- 7114 THEN
            tanh_f := - 2044;
        ELSIF x =- 7113 THEN
            tanh_f := - 2044;
        ELSIF x =- 7112 THEN
            tanh_f := - 2044;
        ELSIF x =- 7111 THEN
            tanh_f := - 2044;
        ELSIF x =- 7110 THEN
            tanh_f := - 2044;
        ELSIF x =- 7109 THEN
            tanh_f := - 2044;
        ELSIF x =- 7108 THEN
            tanh_f := - 2044;
        ELSIF x =- 7107 THEN
            tanh_f := - 2044;
        ELSIF x =- 7106 THEN
            tanh_f := - 2044;
        ELSIF x =- 7105 THEN
            tanh_f := - 2044;
        ELSIF x =- 7104 THEN
            tanh_f := - 2044;
        ELSIF x =- 7103 THEN
            tanh_f := - 2044;
        ELSIF x =- 7102 THEN
            tanh_f := - 2044;
        ELSIF x =- 7101 THEN
            tanh_f := - 2044;
        ELSIF x =- 7100 THEN
            tanh_f := - 2044;
        ELSIF x =- 7099 THEN
            tanh_f := - 2044;
        ELSIF x =- 7098 THEN
            tanh_f := - 2044;
        ELSIF x =- 7097 THEN
            tanh_f := - 2044;
        ELSIF x =- 7096 THEN
            tanh_f := - 2044;
        ELSIF x =- 7095 THEN
            tanh_f := - 2044;
        ELSIF x =- 7094 THEN
            tanh_f := - 2044;
        ELSIF x =- 7093 THEN
            tanh_f := - 2044;
        ELSIF x =- 7092 THEN
            tanh_f := - 2044;
        ELSIF x =- 7091 THEN
            tanh_f := - 2044;
        ELSIF x =- 7090 THEN
            tanh_f := - 2044;
        ELSIF x =- 7089 THEN
            tanh_f := - 2044;
        ELSIF x =- 7088 THEN
            tanh_f := - 2044;
        ELSIF x =- 7087 THEN
            tanh_f := - 2044;
        ELSIF x =- 7086 THEN
            tanh_f := - 2044;
        ELSIF x =- 7085 THEN
            tanh_f := - 2044;
        ELSIF x =- 7084 THEN
            tanh_f := - 2044;
        ELSIF x =- 7083 THEN
            tanh_f := - 2044;
        ELSIF x =- 7082 THEN
            tanh_f := - 2044;
        ELSIF x =- 7081 THEN
            tanh_f := - 2044;
        ELSIF x =- 7080 THEN
            tanh_f := - 2044;
        ELSIF x =- 7079 THEN
            tanh_f := - 2044;
        ELSIF x =- 7078 THEN
            tanh_f := - 2044;
        ELSIF x =- 7077 THEN
            tanh_f := - 2044;
        ELSIF x =- 7076 THEN
            tanh_f := - 2044;
        ELSIF x =- 7075 THEN
            tanh_f := - 2044;
        ELSIF x =- 7074 THEN
            tanh_f := - 2044;
        ELSIF x =- 7073 THEN
            tanh_f := - 2044;
        ELSIF x =- 7072 THEN
            tanh_f := - 2044;
        ELSIF x =- 7071 THEN
            tanh_f := - 2044;
        ELSIF x =- 7070 THEN
            tanh_f := - 2044;
        ELSIF x =- 7069 THEN
            tanh_f := - 2044;
        ELSIF x =- 7068 THEN
            tanh_f := - 2044;
        ELSIF x =- 7067 THEN
            tanh_f := - 2044;
        ELSIF x =- 7066 THEN
            tanh_f := - 2044;
        ELSIF x =- 7065 THEN
            tanh_f := - 2044;
        ELSIF x =- 7064 THEN
            tanh_f := - 2044;
        ELSIF x =- 7063 THEN
            tanh_f := - 2044;
        ELSIF x =- 7062 THEN
            tanh_f := - 2044;
        ELSIF x =- 7061 THEN
            tanh_f := - 2044;
        ELSIF x =- 7060 THEN
            tanh_f := - 2044;
        ELSIF x =- 7059 THEN
            tanh_f := - 2044;
        ELSIF x =- 7058 THEN
            tanh_f := - 2044;
        ELSIF x =- 7057 THEN
            tanh_f := - 2044;
        ELSIF x =- 7056 THEN
            tanh_f := - 2044;
        ELSIF x =- 7055 THEN
            tanh_f := - 2044;
        ELSIF x =- 7054 THEN
            tanh_f := - 2044;
        ELSIF x =- 7053 THEN
            tanh_f := - 2044;
        ELSIF x =- 7052 THEN
            tanh_f := - 2044;
        ELSIF x =- 7051 THEN
            tanh_f := - 2044;
        ELSIF x =- 7050 THEN
            tanh_f := - 2044;
        ELSIF x =- 7049 THEN
            tanh_f := - 2044;
        ELSIF x =- 7048 THEN
            tanh_f := - 2044;
        ELSIF x =- 7047 THEN
            tanh_f := - 2044;
        ELSIF x =- 7046 THEN
            tanh_f := - 2044;
        ELSIF x =- 7045 THEN
            tanh_f := - 2044;
        ELSIF x =- 7044 THEN
            tanh_f := - 2044;
        ELSIF x =- 7043 THEN
            tanh_f := - 2044;
        ELSIF x =- 7042 THEN
            tanh_f := - 2044;
        ELSIF x =- 7041 THEN
            tanh_f := - 2044;
        ELSIF x =- 7040 THEN
            tanh_f := - 2044;
        ELSIF x =- 7039 THEN
            tanh_f := - 2044;
        ELSIF x =- 7038 THEN
            tanh_f := - 2044;
        ELSIF x =- 7037 THEN
            tanh_f := - 2044;
        ELSIF x =- 7036 THEN
            tanh_f := - 2044;
        ELSIF x =- 7035 THEN
            tanh_f := - 2044;
        ELSIF x =- 7034 THEN
            tanh_f := - 2044;
        ELSIF x =- 7033 THEN
            tanh_f := - 2044;
        ELSIF x =- 7032 THEN
            tanh_f := - 2044;
        ELSIF x =- 7031 THEN
            tanh_f := - 2044;
        ELSIF x =- 7030 THEN
            tanh_f := - 2044;
        ELSIF x =- 7029 THEN
            tanh_f := - 2044;
        ELSIF x =- 7028 THEN
            tanh_f := - 2044;
        ELSIF x =- 7027 THEN
            tanh_f := - 2044;
        ELSIF x =- 7026 THEN
            tanh_f := - 2044;
        ELSIF x =- 7025 THEN
            tanh_f := - 2044;
        ELSIF x =- 7024 THEN
            tanh_f := - 2044;
        ELSIF x =- 7023 THEN
            tanh_f := - 2044;
        ELSIF x =- 7022 THEN
            tanh_f := - 2044;
        ELSIF x =- 7021 THEN
            tanh_f := - 2044;
        ELSIF x =- 7020 THEN
            tanh_f := - 2044;
        ELSIF x =- 7019 THEN
            tanh_f := - 2044;
        ELSIF x =- 7018 THEN
            tanh_f := - 2044;
        ELSIF x =- 7017 THEN
            tanh_f := - 2044;
        ELSIF x =- 7016 THEN
            tanh_f := - 2044;
        ELSIF x =- 7015 THEN
            tanh_f := - 2044;
        ELSIF x =- 7014 THEN
            tanh_f := - 2044;
        ELSIF x =- 7013 THEN
            tanh_f := - 2044;
        ELSIF x =- 7012 THEN
            tanh_f := - 2044;
        ELSIF x =- 7011 THEN
            tanh_f := - 2044;
        ELSIF x =- 7010 THEN
            tanh_f := - 2044;
        ELSIF x =- 7009 THEN
            tanh_f := - 2044;
        ELSIF x =- 7008 THEN
            tanh_f := - 2044;
        ELSIF x =- 7007 THEN
            tanh_f := - 2044;
        ELSIF x =- 7006 THEN
            tanh_f := - 2044;
        ELSIF x =- 7005 THEN
            tanh_f := - 2044;
        ELSIF x =- 7004 THEN
            tanh_f := - 2044;
        ELSIF x =- 7003 THEN
            tanh_f := - 2044;
        ELSIF x =- 7002 THEN
            tanh_f := - 2044;
        ELSIF x =- 7001 THEN
            tanh_f := - 2044;
        ELSIF x =- 7000 THEN
            tanh_f := - 2044;
        ELSIF x =- 6999 THEN
            tanh_f := - 2044;
        ELSIF x =- 6998 THEN
            tanh_f := - 2044;
        ELSIF x =- 6997 THEN
            tanh_f := - 2044;
        ELSIF x =- 6996 THEN
            tanh_f := - 2044;
        ELSIF x =- 6995 THEN
            tanh_f := - 2044;
        ELSIF x =- 6994 THEN
            tanh_f := - 2044;
        ELSIF x =- 6993 THEN
            tanh_f := - 2044;
        ELSIF x =- 6992 THEN
            tanh_f := - 2044;
        ELSIF x =- 6991 THEN
            tanh_f := - 2044;
        ELSIF x =- 6990 THEN
            tanh_f := - 2044;
        ELSIF x =- 6989 THEN
            tanh_f := - 2044;
        ELSIF x =- 6988 THEN
            tanh_f := - 2044;
        ELSIF x =- 6987 THEN
            tanh_f := - 2044;
        ELSIF x =- 6986 THEN
            tanh_f := - 2044;
        ELSIF x =- 6985 THEN
            tanh_f := - 2044;
        ELSIF x =- 6984 THEN
            tanh_f := - 2044;
        ELSIF x =- 6983 THEN
            tanh_f := - 2044;
        ELSIF x =- 6982 THEN
            tanh_f := - 2044;
        ELSIF x =- 6981 THEN
            tanh_f := - 2044;
        ELSIF x =- 6980 THEN
            tanh_f := - 2044;
        ELSIF x =- 6979 THEN
            tanh_f := - 2044;
        ELSIF x =- 6978 THEN
            tanh_f := - 2044;
        ELSIF x =- 6977 THEN
            tanh_f := - 2044;
        ELSIF x =- 6976 THEN
            tanh_f := - 2044;
        ELSIF x =- 6975 THEN
            tanh_f := - 2044;
        ELSIF x =- 6974 THEN
            tanh_f := - 2044;
        ELSIF x =- 6973 THEN
            tanh_f := - 2044;
        ELSIF x =- 6972 THEN
            tanh_f := - 2044;
        ELSIF x =- 6971 THEN
            tanh_f := - 2044;
        ELSIF x =- 6970 THEN
            tanh_f := - 2044;
        ELSIF x =- 6969 THEN
            tanh_f := - 2044;
        ELSIF x =- 6968 THEN
            tanh_f := - 2044;
        ELSIF x =- 6967 THEN
            tanh_f := - 2044;
        ELSIF x =- 6966 THEN
            tanh_f := - 2044;
        ELSIF x =- 6965 THEN
            tanh_f := - 2044;
        ELSIF x =- 6964 THEN
            tanh_f := - 2044;
        ELSIF x =- 6963 THEN
            tanh_f := - 2044;
        ELSIF x =- 6962 THEN
            tanh_f := - 2044;
        ELSIF x =- 6961 THEN
            tanh_f := - 2044;
        ELSIF x =- 6960 THEN
            tanh_f := - 2044;
        ELSIF x =- 6959 THEN
            tanh_f := - 2044;
        ELSIF x =- 6958 THEN
            tanh_f := - 2044;
        ELSIF x =- 6957 THEN
            tanh_f := - 2044;
        ELSIF x =- 6956 THEN
            tanh_f := - 2044;
        ELSIF x =- 6955 THEN
            tanh_f := - 2044;
        ELSIF x =- 6954 THEN
            tanh_f := - 2044;
        ELSIF x =- 6953 THEN
            tanh_f := - 2044;
        ELSIF x =- 6952 THEN
            tanh_f := - 2044;
        ELSIF x =- 6951 THEN
            tanh_f := - 2044;
        ELSIF x =- 6950 THEN
            tanh_f := - 2044;
        ELSIF x =- 6949 THEN
            tanh_f := - 2044;
        ELSIF x =- 6948 THEN
            tanh_f := - 2044;
        ELSIF x =- 6947 THEN
            tanh_f := - 2044;
        ELSIF x =- 6946 THEN
            tanh_f := - 2044;
        ELSIF x =- 6945 THEN
            tanh_f := - 2044;
        ELSIF x =- 6944 THEN
            tanh_f := - 2044;
        ELSIF x =- 6943 THEN
            tanh_f := - 2044;
        ELSIF x =- 6942 THEN
            tanh_f := - 2044;
        ELSIF x =- 6941 THEN
            tanh_f := - 2044;
        ELSIF x =- 6940 THEN
            tanh_f := - 2044;
        ELSIF x =- 6939 THEN
            tanh_f := - 2044;
        ELSIF x =- 6938 THEN
            tanh_f := - 2044;
        ELSIF x =- 6937 THEN
            tanh_f := - 2044;
        ELSIF x =- 6936 THEN
            tanh_f := - 2044;
        ELSIF x =- 6935 THEN
            tanh_f := - 2044;
        ELSIF x =- 6934 THEN
            tanh_f := - 2044;
        ELSIF x =- 6933 THEN
            tanh_f := - 2044;
        ELSIF x =- 6932 THEN
            tanh_f := - 2044;
        ELSIF x =- 6931 THEN
            tanh_f := - 2044;
        ELSIF x =- 6930 THEN
            tanh_f := - 2044;
        ELSIF x =- 6929 THEN
            tanh_f := - 2044;
        ELSIF x =- 6928 THEN
            tanh_f := - 2044;
        ELSIF x =- 6927 THEN
            tanh_f := - 2044;
        ELSIF x =- 6926 THEN
            tanh_f := - 2044;
        ELSIF x =- 6925 THEN
            tanh_f := - 2044;
        ELSIF x =- 6924 THEN
            tanh_f := - 2044;
        ELSIF x =- 6923 THEN
            tanh_f := - 2044;
        ELSIF x =- 6922 THEN
            tanh_f := - 2044;
        ELSIF x =- 6921 THEN
            tanh_f := - 2044;
        ELSIF x =- 6920 THEN
            tanh_f := - 2044;
        ELSIF x =- 6919 THEN
            tanh_f := - 2044;
        ELSIF x =- 6918 THEN
            tanh_f := - 2044;
        ELSIF x =- 6917 THEN
            tanh_f := - 2044;
        ELSIF x =- 6916 THEN
            tanh_f := - 2044;
        ELSIF x =- 6915 THEN
            tanh_f := - 2044;
        ELSIF x =- 6914 THEN
            tanh_f := - 2044;
        ELSIF x =- 6913 THEN
            tanh_f := - 2044;
        ELSIF x =- 6912 THEN
            tanh_f := - 2044;
        ELSIF x =- 6911 THEN
            tanh_f := - 2042;
        ELSIF x =- 6910 THEN
            tanh_f := - 2042;
        ELSIF x =- 6909 THEN
            tanh_f := - 2042;
        ELSIF x =- 6908 THEN
            tanh_f := - 2042;
        ELSIF x =- 6907 THEN
            tanh_f := - 2042;
        ELSIF x =- 6906 THEN
            tanh_f := - 2042;
        ELSIF x =- 6905 THEN
            tanh_f := - 2042;
        ELSIF x =- 6904 THEN
            tanh_f := - 2042;
        ELSIF x =- 6903 THEN
            tanh_f := - 2042;
        ELSIF x =- 6902 THEN
            tanh_f := - 2042;
        ELSIF x =- 6901 THEN
            tanh_f := - 2042;
        ELSIF x =- 6900 THEN
            tanh_f := - 2042;
        ELSIF x =- 6899 THEN
            tanh_f := - 2042;
        ELSIF x =- 6898 THEN
            tanh_f := - 2042;
        ELSIF x =- 6897 THEN
            tanh_f := - 2042;
        ELSIF x =- 6896 THEN
            tanh_f := - 2042;
        ELSIF x =- 6895 THEN
            tanh_f := - 2042;
        ELSIF x =- 6894 THEN
            tanh_f := - 2042;
        ELSIF x =- 6893 THEN
            tanh_f := - 2042;
        ELSIF x =- 6892 THEN
            tanh_f := - 2042;
        ELSIF x =- 6891 THEN
            tanh_f := - 2042;
        ELSIF x =- 6890 THEN
            tanh_f := - 2042;
        ELSIF x =- 6889 THEN
            tanh_f := - 2042;
        ELSIF x =- 6888 THEN
            tanh_f := - 2042;
        ELSIF x =- 6887 THEN
            tanh_f := - 2042;
        ELSIF x =- 6886 THEN
            tanh_f := - 2042;
        ELSIF x =- 6885 THEN
            tanh_f := - 2042;
        ELSIF x =- 6884 THEN
            tanh_f := - 2042;
        ELSIF x =- 6883 THEN
            tanh_f := - 2042;
        ELSIF x =- 6882 THEN
            tanh_f := - 2042;
        ELSIF x =- 6881 THEN
            tanh_f := - 2042;
        ELSIF x =- 6880 THEN
            tanh_f := - 2042;
        ELSIF x =- 6879 THEN
            tanh_f := - 2042;
        ELSIF x =- 6878 THEN
            tanh_f := - 2042;
        ELSIF x =- 6877 THEN
            tanh_f := - 2042;
        ELSIF x =- 6876 THEN
            tanh_f := - 2042;
        ELSIF x =- 6875 THEN
            tanh_f := - 2042;
        ELSIF x =- 6874 THEN
            tanh_f := - 2042;
        ELSIF x =- 6873 THEN
            tanh_f := - 2042;
        ELSIF x =- 6872 THEN
            tanh_f := - 2042;
        ELSIF x =- 6871 THEN
            tanh_f := - 2042;
        ELSIF x =- 6870 THEN
            tanh_f := - 2042;
        ELSIF x =- 6869 THEN
            tanh_f := - 2042;
        ELSIF x =- 6868 THEN
            tanh_f := - 2042;
        ELSIF x =- 6867 THEN
            tanh_f := - 2042;
        ELSIF x =- 6866 THEN
            tanh_f := - 2042;
        ELSIF x =- 6865 THEN
            tanh_f := - 2042;
        ELSIF x =- 6864 THEN
            tanh_f := - 2042;
        ELSIF x =- 6863 THEN
            tanh_f := - 2042;
        ELSIF x =- 6862 THEN
            tanh_f := - 2042;
        ELSIF x =- 6861 THEN
            tanh_f := - 2042;
        ELSIF x =- 6860 THEN
            tanh_f := - 2042;
        ELSIF x =- 6859 THEN
            tanh_f := - 2042;
        ELSIF x =- 6858 THEN
            tanh_f := - 2042;
        ELSIF x =- 6857 THEN
            tanh_f := - 2042;
        ELSIF x =- 6856 THEN
            tanh_f := - 2042;
        ELSIF x =- 6855 THEN
            tanh_f := - 2042;
        ELSIF x =- 6854 THEN
            tanh_f := - 2042;
        ELSIF x =- 6853 THEN
            tanh_f := - 2042;
        ELSIF x =- 6852 THEN
            tanh_f := - 2042;
        ELSIF x =- 6851 THEN
            tanh_f := - 2042;
        ELSIF x =- 6850 THEN
            tanh_f := - 2042;
        ELSIF x =- 6849 THEN
            tanh_f := - 2042;
        ELSIF x =- 6848 THEN
            tanh_f := - 2042;
        ELSIF x =- 6847 THEN
            tanh_f := - 2042;
        ELSIF x =- 6846 THEN
            tanh_f := - 2042;
        ELSIF x =- 6845 THEN
            tanh_f := - 2042;
        ELSIF x =- 6844 THEN
            tanh_f := - 2042;
        ELSIF x =- 6843 THEN
            tanh_f := - 2042;
        ELSIF x =- 6842 THEN
            tanh_f := - 2042;
        ELSIF x =- 6841 THEN
            tanh_f := - 2042;
        ELSIF x =- 6840 THEN
            tanh_f := - 2042;
        ELSIF x =- 6839 THEN
            tanh_f := - 2042;
        ELSIF x =- 6838 THEN
            tanh_f := - 2042;
        ELSIF x =- 6837 THEN
            tanh_f := - 2042;
        ELSIF x =- 6836 THEN
            tanh_f := - 2042;
        ELSIF x =- 6835 THEN
            tanh_f := - 2042;
        ELSIF x =- 6834 THEN
            tanh_f := - 2042;
        ELSIF x =- 6833 THEN
            tanh_f := - 2042;
        ELSIF x =- 6832 THEN
            tanh_f := - 2042;
        ELSIF x =- 6831 THEN
            tanh_f := - 2042;
        ELSIF x =- 6830 THEN
            tanh_f := - 2042;
        ELSIF x =- 6829 THEN
            tanh_f := - 2042;
        ELSIF x =- 6828 THEN
            tanh_f := - 2042;
        ELSIF x =- 6827 THEN
            tanh_f := - 2042;
        ELSIF x =- 6826 THEN
            tanh_f := - 2042;
        ELSIF x =- 6825 THEN
            tanh_f := - 2042;
        ELSIF x =- 6824 THEN
            tanh_f := - 2042;
        ELSIF x =- 6823 THEN
            tanh_f := - 2042;
        ELSIF x =- 6822 THEN
            tanh_f := - 2042;
        ELSIF x =- 6821 THEN
            tanh_f := - 2042;
        ELSIF x =- 6820 THEN
            tanh_f := - 2042;
        ELSIF x =- 6819 THEN
            tanh_f := - 2042;
        ELSIF x =- 6818 THEN
            tanh_f := - 2042;
        ELSIF x =- 6817 THEN
            tanh_f := - 2042;
        ELSIF x =- 6816 THEN
            tanh_f := - 2042;
        ELSIF x =- 6815 THEN
            tanh_f := - 2042;
        ELSIF x =- 6814 THEN
            tanh_f := - 2042;
        ELSIF x =- 6813 THEN
            tanh_f := - 2042;
        ELSIF x =- 6812 THEN
            tanh_f := - 2042;
        ELSIF x =- 6811 THEN
            tanh_f := - 2042;
        ELSIF x =- 6810 THEN
            tanh_f := - 2042;
        ELSIF x =- 6809 THEN
            tanh_f := - 2042;
        ELSIF x =- 6808 THEN
            tanh_f := - 2042;
        ELSIF x =- 6807 THEN
            tanh_f := - 2042;
        ELSIF x =- 6806 THEN
            tanh_f := - 2042;
        ELSIF x =- 6805 THEN
            tanh_f := - 2042;
        ELSIF x =- 6804 THEN
            tanh_f := - 2042;
        ELSIF x =- 6803 THEN
            tanh_f := - 2042;
        ELSIF x =- 6802 THEN
            tanh_f := - 2042;
        ELSIF x =- 6801 THEN
            tanh_f := - 2042;
        ELSIF x =- 6800 THEN
            tanh_f := - 2042;
        ELSIF x =- 6799 THEN
            tanh_f := - 2042;
        ELSIF x =- 6798 THEN
            tanh_f := - 2042;
        ELSIF x =- 6797 THEN
            tanh_f := - 2042;
        ELSIF x =- 6796 THEN
            tanh_f := - 2042;
        ELSIF x =- 6795 THEN
            tanh_f := - 2042;
        ELSIF x =- 6794 THEN
            tanh_f := - 2042;
        ELSIF x =- 6793 THEN
            tanh_f := - 2042;
        ELSIF x =- 6792 THEN
            tanh_f := - 2042;
        ELSIF x =- 6791 THEN
            tanh_f := - 2042;
        ELSIF x =- 6790 THEN
            tanh_f := - 2042;
        ELSIF x =- 6789 THEN
            tanh_f := - 2042;
        ELSIF x =- 6788 THEN
            tanh_f := - 2042;
        ELSIF x =- 6787 THEN
            tanh_f := - 2042;
        ELSIF x =- 6786 THEN
            tanh_f := - 2042;
        ELSIF x =- 6785 THEN
            tanh_f := - 2042;
        ELSIF x =- 6784 THEN
            tanh_f := - 2042;
        ELSIF x =- 6783 THEN
            tanh_f := - 2042;
        ELSIF x =- 6782 THEN
            tanh_f := - 2042;
        ELSIF x =- 6781 THEN
            tanh_f := - 2042;
        ELSIF x =- 6780 THEN
            tanh_f := - 2042;
        ELSIF x =- 6779 THEN
            tanh_f := - 2042;
        ELSIF x =- 6778 THEN
            tanh_f := - 2042;
        ELSIF x =- 6777 THEN
            tanh_f := - 2042;
        ELSIF x =- 6776 THEN
            tanh_f := - 2042;
        ELSIF x =- 6775 THEN
            tanh_f := - 2042;
        ELSIF x =- 6774 THEN
            tanh_f := - 2042;
        ELSIF x =- 6773 THEN
            tanh_f := - 2042;
        ELSIF x =- 6772 THEN
            tanh_f := - 2042;
        ELSIF x =- 6771 THEN
            tanh_f := - 2042;
        ELSIF x =- 6770 THEN
            tanh_f := - 2042;
        ELSIF x =- 6769 THEN
            tanh_f := - 2042;
        ELSIF x =- 6768 THEN
            tanh_f := - 2042;
        ELSIF x =- 6767 THEN
            tanh_f := - 2042;
        ELSIF x =- 6766 THEN
            tanh_f := - 2042;
        ELSIF x =- 6765 THEN
            tanh_f := - 2042;
        ELSIF x =- 6764 THEN
            tanh_f := - 2042;
        ELSIF x =- 6763 THEN
            tanh_f := - 2042;
        ELSIF x =- 6762 THEN
            tanh_f := - 2042;
        ELSIF x =- 6761 THEN
            tanh_f := - 2042;
        ELSIF x =- 6760 THEN
            tanh_f := - 2042;
        ELSIF x =- 6759 THEN
            tanh_f := - 2042;
        ELSIF x =- 6758 THEN
            tanh_f := - 2042;
        ELSIF x =- 6757 THEN
            tanh_f := - 2042;
        ELSIF x =- 6756 THEN
            tanh_f := - 2042;
        ELSIF x =- 6755 THEN
            tanh_f := - 2042;
        ELSIF x =- 6754 THEN
            tanh_f := - 2042;
        ELSIF x =- 6753 THEN
            tanh_f := - 2042;
        ELSIF x =- 6752 THEN
            tanh_f := - 2042;
        ELSIF x =- 6751 THEN
            tanh_f := - 2042;
        ELSIF x =- 6750 THEN
            tanh_f := - 2042;
        ELSIF x =- 6749 THEN
            tanh_f := - 2042;
        ELSIF x =- 6748 THEN
            tanh_f := - 2042;
        ELSIF x =- 6747 THEN
            tanh_f := - 2042;
        ELSIF x =- 6746 THEN
            tanh_f := - 2042;
        ELSIF x =- 6745 THEN
            tanh_f := - 2042;
        ELSIF x =- 6744 THEN
            tanh_f := - 2042;
        ELSIF x =- 6743 THEN
            tanh_f := - 2042;
        ELSIF x =- 6742 THEN
            tanh_f := - 2042;
        ELSIF x =- 6741 THEN
            tanh_f := - 2042;
        ELSIF x =- 6740 THEN
            tanh_f := - 2042;
        ELSIF x =- 6739 THEN
            tanh_f := - 2042;
        ELSIF x =- 6738 THEN
            tanh_f := - 2042;
        ELSIF x =- 6737 THEN
            tanh_f := - 2042;
        ELSIF x =- 6736 THEN
            tanh_f := - 2042;
        ELSIF x =- 6735 THEN
            tanh_f := - 2042;
        ELSIF x =- 6734 THEN
            tanh_f := - 2042;
        ELSIF x =- 6733 THEN
            tanh_f := - 2042;
        ELSIF x =- 6732 THEN
            tanh_f := - 2042;
        ELSIF x =- 6731 THEN
            tanh_f := - 2042;
        ELSIF x =- 6730 THEN
            tanh_f := - 2042;
        ELSIF x =- 6729 THEN
            tanh_f := - 2042;
        ELSIF x =- 6728 THEN
            tanh_f := - 2042;
        ELSIF x =- 6727 THEN
            tanh_f := - 2042;
        ELSIF x =- 6726 THEN
            tanh_f := - 2042;
        ELSIF x =- 6725 THEN
            tanh_f := - 2042;
        ELSIF x =- 6724 THEN
            tanh_f := - 2042;
        ELSIF x =- 6723 THEN
            tanh_f := - 2042;
        ELSIF x =- 6722 THEN
            tanh_f := - 2042;
        ELSIF x =- 6721 THEN
            tanh_f := - 2042;
        ELSIF x =- 6720 THEN
            tanh_f := - 2042;
        ELSIF x =- 6719 THEN
            tanh_f := - 2042;
        ELSIF x =- 6718 THEN
            tanh_f := - 2042;
        ELSIF x =- 6717 THEN
            tanh_f := - 2042;
        ELSIF x =- 6716 THEN
            tanh_f := - 2042;
        ELSIF x =- 6715 THEN
            tanh_f := - 2042;
        ELSIF x =- 6714 THEN
            tanh_f := - 2042;
        ELSIF x =- 6713 THEN
            tanh_f := - 2042;
        ELSIF x =- 6712 THEN
            tanh_f := - 2042;
        ELSIF x =- 6711 THEN
            tanh_f := - 2042;
        ELSIF x =- 6710 THEN
            tanh_f := - 2042;
        ELSIF x =- 6709 THEN
            tanh_f := - 2042;
        ELSIF x =- 6708 THEN
            tanh_f := - 2042;
        ELSIF x =- 6707 THEN
            tanh_f := - 2042;
        ELSIF x =- 6706 THEN
            tanh_f := - 2042;
        ELSIF x =- 6705 THEN
            tanh_f := - 2042;
        ELSIF x =- 6704 THEN
            tanh_f := - 2042;
        ELSIF x =- 6703 THEN
            tanh_f := - 2042;
        ELSIF x =- 6702 THEN
            tanh_f := - 2042;
        ELSIF x =- 6701 THEN
            tanh_f := - 2042;
        ELSIF x =- 6700 THEN
            tanh_f := - 2042;
        ELSIF x =- 6699 THEN
            tanh_f := - 2042;
        ELSIF x =- 6698 THEN
            tanh_f := - 2042;
        ELSIF x =- 6697 THEN
            tanh_f := - 2042;
        ELSIF x =- 6696 THEN
            tanh_f := - 2042;
        ELSIF x =- 6695 THEN
            tanh_f := - 2042;
        ELSIF x =- 6694 THEN
            tanh_f := - 2042;
        ELSIF x =- 6693 THEN
            tanh_f := - 2042;
        ELSIF x =- 6692 THEN
            tanh_f := - 2042;
        ELSIF x =- 6691 THEN
            tanh_f := - 2042;
        ELSIF x =- 6690 THEN
            tanh_f := - 2042;
        ELSIF x =- 6689 THEN
            tanh_f := - 2042;
        ELSIF x =- 6688 THEN
            tanh_f := - 2042;
        ELSIF x =- 6687 THEN
            tanh_f := - 2042;
        ELSIF x =- 6686 THEN
            tanh_f := - 2042;
        ELSIF x =- 6685 THEN
            tanh_f := - 2042;
        ELSIF x =- 6684 THEN
            tanh_f := - 2042;
        ELSIF x =- 6683 THEN
            tanh_f := - 2042;
        ELSIF x =- 6682 THEN
            tanh_f := - 2042;
        ELSIF x =- 6681 THEN
            tanh_f := - 2042;
        ELSIF x =- 6680 THEN
            tanh_f := - 2042;
        ELSIF x =- 6679 THEN
            tanh_f := - 2042;
        ELSIF x =- 6678 THEN
            tanh_f := - 2042;
        ELSIF x =- 6677 THEN
            tanh_f := - 2042;
        ELSIF x =- 6676 THEN
            tanh_f := - 2042;
        ELSIF x =- 6675 THEN
            tanh_f := - 2042;
        ELSIF x =- 6674 THEN
            tanh_f := - 2042;
        ELSIF x =- 6673 THEN
            tanh_f := - 2042;
        ELSIF x =- 6672 THEN
            tanh_f := - 2042;
        ELSIF x =- 6671 THEN
            tanh_f := - 2042;
        ELSIF x =- 6670 THEN
            tanh_f := - 2042;
        ELSIF x =- 6669 THEN
            tanh_f := - 2042;
        ELSIF x =- 6668 THEN
            tanh_f := - 2042;
        ELSIF x =- 6667 THEN
            tanh_f := - 2042;
        ELSIF x =- 6666 THEN
            tanh_f := - 2042;
        ELSIF x =- 6665 THEN
            tanh_f := - 2042;
        ELSIF x =- 6664 THEN
            tanh_f := - 2042;
        ELSIF x =- 6663 THEN
            tanh_f := - 2042;
        ELSIF x =- 6662 THEN
            tanh_f := - 2042;
        ELSIF x =- 6661 THEN
            tanh_f := - 2042;
        ELSIF x =- 6660 THEN
            tanh_f := - 2042;
        ELSIF x =- 6659 THEN
            tanh_f := - 2042;
        ELSIF x =- 6658 THEN
            tanh_f := - 2042;
        ELSIF x =- 6657 THEN
            tanh_f := - 2042;
        ELSIF x =- 6656 THEN
            tanh_f := - 2042;
        ELSIF x =- 6655 THEN
            tanh_f := - 2042;
        ELSIF x =- 6654 THEN
            tanh_f := - 2042;
        ELSIF x =- 6653 THEN
            tanh_f := - 2042;
        ELSIF x =- 6652 THEN
            tanh_f := - 2042;
        ELSIF x =- 6651 THEN
            tanh_f := - 2042;
        ELSIF x =- 6650 THEN
            tanh_f := - 2042;
        ELSIF x =- 6649 THEN
            tanh_f := - 2042;
        ELSIF x =- 6648 THEN
            tanh_f := - 2042;
        ELSIF x =- 6647 THEN
            tanh_f := - 2042;
        ELSIF x =- 6646 THEN
            tanh_f := - 2042;
        ELSIF x =- 6645 THEN
            tanh_f := - 2042;
        ELSIF x =- 6644 THEN
            tanh_f := - 2042;
        ELSIF x =- 6643 THEN
            tanh_f := - 2042;
        ELSIF x =- 6642 THEN
            tanh_f := - 2042;
        ELSIF x =- 6641 THEN
            tanh_f := - 2042;
        ELSIF x =- 6640 THEN
            tanh_f := - 2042;
        ELSIF x =- 6639 THEN
            tanh_f := - 2042;
        ELSIF x =- 6638 THEN
            tanh_f := - 2042;
        ELSIF x =- 6637 THEN
            tanh_f := - 2042;
        ELSIF x =- 6636 THEN
            tanh_f := - 2042;
        ELSIF x =- 6635 THEN
            tanh_f := - 2042;
        ELSIF x =- 6634 THEN
            tanh_f := - 2042;
        ELSIF x =- 6633 THEN
            tanh_f := - 2042;
        ELSIF x =- 6632 THEN
            tanh_f := - 2042;
        ELSIF x =- 6631 THEN
            tanh_f := - 2042;
        ELSIF x =- 6630 THEN
            tanh_f := - 2042;
        ELSIF x =- 6629 THEN
            tanh_f := - 2042;
        ELSIF x =- 6628 THEN
            tanh_f := - 2042;
        ELSIF x =- 6627 THEN
            tanh_f := - 2042;
        ELSIF x =- 6626 THEN
            tanh_f := - 2042;
        ELSIF x =- 6625 THEN
            tanh_f := - 2042;
        ELSIF x =- 6624 THEN
            tanh_f := - 2042;
        ELSIF x =- 6623 THEN
            tanh_f := - 2042;
        ELSIF x =- 6622 THEN
            tanh_f := - 2042;
        ELSIF x =- 6621 THEN
            tanh_f := - 2042;
        ELSIF x =- 6620 THEN
            tanh_f := - 2042;
        ELSIF x =- 6619 THEN
            tanh_f := - 2042;
        ELSIF x =- 6618 THEN
            tanh_f := - 2042;
        ELSIF x =- 6617 THEN
            tanh_f := - 2042;
        ELSIF x =- 6616 THEN
            tanh_f := - 2042;
        ELSIF x =- 6615 THEN
            tanh_f := - 2042;
        ELSIF x =- 6614 THEN
            tanh_f := - 2042;
        ELSIF x =- 6613 THEN
            tanh_f := - 2042;
        ELSIF x =- 6612 THEN
            tanh_f := - 2042;
        ELSIF x =- 6611 THEN
            tanh_f := - 2042;
        ELSIF x =- 6610 THEN
            tanh_f := - 2042;
        ELSIF x =- 6609 THEN
            tanh_f := - 2042;
        ELSIF x =- 6608 THEN
            tanh_f := - 2042;
        ELSIF x =- 6607 THEN
            tanh_f := - 2042;
        ELSIF x =- 6606 THEN
            tanh_f := - 2042;
        ELSIF x =- 6605 THEN
            tanh_f := - 2042;
        ELSIF x =- 6604 THEN
            tanh_f := - 2042;
        ELSIF x =- 6603 THEN
            tanh_f := - 2042;
        ELSIF x =- 6602 THEN
            tanh_f := - 2042;
        ELSIF x =- 6601 THEN
            tanh_f := - 2042;
        ELSIF x =- 6600 THEN
            tanh_f := - 2042;
        ELSIF x =- 6599 THEN
            tanh_f := - 2042;
        ELSIF x =- 6598 THEN
            tanh_f := - 2042;
        ELSIF x =- 6597 THEN
            tanh_f := - 2042;
        ELSIF x =- 6596 THEN
            tanh_f := - 2042;
        ELSIF x =- 6595 THEN
            tanh_f := - 2042;
        ELSIF x =- 6594 THEN
            tanh_f := - 2042;
        ELSIF x =- 6593 THEN
            tanh_f := - 2042;
        ELSIF x =- 6592 THEN
            tanh_f := - 2042;
        ELSIF x =- 6591 THEN
            tanh_f := - 2042;
        ELSIF x =- 6590 THEN
            tanh_f := - 2042;
        ELSIF x =- 6589 THEN
            tanh_f := - 2042;
        ELSIF x =- 6588 THEN
            tanh_f := - 2042;
        ELSIF x =- 6587 THEN
            tanh_f := - 2042;
        ELSIF x =- 6586 THEN
            tanh_f := - 2042;
        ELSIF x =- 6585 THEN
            tanh_f := - 2042;
        ELSIF x =- 6584 THEN
            tanh_f := - 2042;
        ELSIF x =- 6583 THEN
            tanh_f := - 2042;
        ELSIF x =- 6582 THEN
            tanh_f := - 2042;
        ELSIF x =- 6581 THEN
            tanh_f := - 2042;
        ELSIF x =- 6580 THEN
            tanh_f := - 2042;
        ELSIF x =- 6579 THEN
            tanh_f := - 2042;
        ELSIF x =- 6578 THEN
            tanh_f := - 2042;
        ELSIF x =- 6577 THEN
            tanh_f := - 2042;
        ELSIF x =- 6576 THEN
            tanh_f := - 2042;
        ELSIF x =- 6575 THEN
            tanh_f := - 2042;
        ELSIF x =- 6574 THEN
            tanh_f := - 2042;
        ELSIF x =- 6573 THEN
            tanh_f := - 2042;
        ELSIF x =- 6572 THEN
            tanh_f := - 2042;
        ELSIF x =- 6571 THEN
            tanh_f := - 2042;
        ELSIF x =- 6570 THEN
            tanh_f := - 2042;
        ELSIF x =- 6569 THEN
            tanh_f := - 2042;
        ELSIF x =- 6568 THEN
            tanh_f := - 2042;
        ELSIF x =- 6567 THEN
            tanh_f := - 2042;
        ELSIF x =- 6566 THEN
            tanh_f := - 2042;
        ELSIF x =- 6565 THEN
            tanh_f := - 2042;
        ELSIF x =- 6564 THEN
            tanh_f := - 2042;
        ELSIF x =- 6563 THEN
            tanh_f := - 2042;
        ELSIF x =- 6562 THEN
            tanh_f := - 2042;
        ELSIF x =- 6561 THEN
            tanh_f := - 2042;
        ELSIF x =- 6560 THEN
            tanh_f := - 2042;
        ELSIF x =- 6559 THEN
            tanh_f := - 2042;
        ELSIF x =- 6558 THEN
            tanh_f := - 2042;
        ELSIF x =- 6557 THEN
            tanh_f := - 2042;
        ELSIF x =- 6556 THEN
            tanh_f := - 2042;
        ELSIF x =- 6555 THEN
            tanh_f := - 2042;
        ELSIF x =- 6554 THEN
            tanh_f := - 2042;
        ELSIF x =- 6553 THEN
            tanh_f := - 2042;
        ELSIF x =- 6552 THEN
            tanh_f := - 2042;
        ELSIF x =- 6551 THEN
            tanh_f := - 2042;
        ELSIF x =- 6550 THEN
            tanh_f := - 2042;
        ELSIF x =- 6549 THEN
            tanh_f := - 2042;
        ELSIF x =- 6548 THEN
            tanh_f := - 2042;
        ELSIF x =- 6547 THEN
            tanh_f := - 2042;
        ELSIF x =- 6546 THEN
            tanh_f := - 2042;
        ELSIF x =- 6545 THEN
            tanh_f := - 2042;
        ELSIF x =- 6544 THEN
            tanh_f := - 2042;
        ELSIF x =- 6543 THEN
            tanh_f := - 2042;
        ELSIF x =- 6542 THEN
            tanh_f := - 2042;
        ELSIF x =- 6541 THEN
            tanh_f := - 2042;
        ELSIF x =- 6540 THEN
            tanh_f := - 2042;
        ELSIF x =- 6539 THEN
            tanh_f := - 2042;
        ELSIF x =- 6538 THEN
            tanh_f := - 2042;
        ELSIF x =- 6537 THEN
            tanh_f := - 2042;
        ELSIF x =- 6536 THEN
            tanh_f := - 2042;
        ELSIF x =- 6535 THEN
            tanh_f := - 2042;
        ELSIF x =- 6534 THEN
            tanh_f := - 2042;
        ELSIF x =- 6533 THEN
            tanh_f := - 2042;
        ELSIF x =- 6532 THEN
            tanh_f := - 2042;
        ELSIF x =- 6531 THEN
            tanh_f := - 2042;
        ELSIF x =- 6530 THEN
            tanh_f := - 2042;
        ELSIF x =- 6529 THEN
            tanh_f := - 2042;
        ELSIF x =- 6528 THEN
            tanh_f := - 2042;
        ELSIF x =- 6527 THEN
            tanh_f := - 2042;
        ELSIF x =- 6526 THEN
            tanh_f := - 2042;
        ELSIF x =- 6525 THEN
            tanh_f := - 2042;
        ELSIF x =- 6524 THEN
            tanh_f := - 2042;
        ELSIF x =- 6523 THEN
            tanh_f := - 2042;
        ELSIF x =- 6522 THEN
            tanh_f := - 2042;
        ELSIF x =- 6521 THEN
            tanh_f := - 2042;
        ELSIF x =- 6520 THEN
            tanh_f := - 2042;
        ELSIF x =- 6519 THEN
            tanh_f := - 2042;
        ELSIF x =- 6518 THEN
            tanh_f := - 2042;
        ELSIF x =- 6517 THEN
            tanh_f := - 2042;
        ELSIF x =- 6516 THEN
            tanh_f := - 2042;
        ELSIF x =- 6515 THEN
            tanh_f := - 2042;
        ELSIF x =- 6514 THEN
            tanh_f := - 2042;
        ELSIF x =- 6513 THEN
            tanh_f := - 2042;
        ELSIF x =- 6512 THEN
            tanh_f := - 2042;
        ELSIF x =- 6511 THEN
            tanh_f := - 2042;
        ELSIF x =- 6510 THEN
            tanh_f := - 2042;
        ELSIF x =- 6509 THEN
            tanh_f := - 2042;
        ELSIF x =- 6508 THEN
            tanh_f := - 2042;
        ELSIF x =- 6507 THEN
            tanh_f := - 2042;
        ELSIF x =- 6506 THEN
            tanh_f := - 2042;
        ELSIF x =- 6505 THEN
            tanh_f := - 2042;
        ELSIF x =- 6504 THEN
            tanh_f := - 2042;
        ELSIF x =- 6503 THEN
            tanh_f := - 2042;
        ELSIF x =- 6502 THEN
            tanh_f := - 2042;
        ELSIF x =- 6501 THEN
            tanh_f := - 2042;
        ELSIF x =- 6500 THEN
            tanh_f := - 2042;
        ELSIF x =- 6499 THEN
            tanh_f := - 2042;
        ELSIF x =- 6498 THEN
            tanh_f := - 2042;
        ELSIF x =- 6497 THEN
            tanh_f := - 2042;
        ELSIF x =- 6496 THEN
            tanh_f := - 2042;
        ELSIF x =- 6495 THEN
            tanh_f := - 2042;
        ELSIF x =- 6494 THEN
            tanh_f := - 2042;
        ELSIF x =- 6493 THEN
            tanh_f := - 2042;
        ELSIF x =- 6492 THEN
            tanh_f := - 2042;
        ELSIF x =- 6491 THEN
            tanh_f := - 2042;
        ELSIF x =- 6490 THEN
            tanh_f := - 2042;
        ELSIF x =- 6489 THEN
            tanh_f := - 2042;
        ELSIF x =- 6488 THEN
            tanh_f := - 2042;
        ELSIF x =- 6487 THEN
            tanh_f := - 2042;
        ELSIF x =- 6486 THEN
            tanh_f := - 2042;
        ELSIF x =- 6485 THEN
            tanh_f := - 2042;
        ELSIF x =- 6484 THEN
            tanh_f := - 2042;
        ELSIF x =- 6483 THEN
            tanh_f := - 2042;
        ELSIF x =- 6482 THEN
            tanh_f := - 2042;
        ELSIF x =- 6481 THEN
            tanh_f := - 2042;
        ELSIF x =- 6480 THEN
            tanh_f := - 2042;
        ELSIF x =- 6479 THEN
            tanh_f := - 2042;
        ELSIF x =- 6478 THEN
            tanh_f := - 2042;
        ELSIF x =- 6477 THEN
            tanh_f := - 2042;
        ELSIF x =- 6476 THEN
            tanh_f := - 2042;
        ELSIF x =- 6475 THEN
            tanh_f := - 2042;
        ELSIF x =- 6474 THEN
            tanh_f := - 2042;
        ELSIF x =- 6473 THEN
            tanh_f := - 2042;
        ELSIF x =- 6472 THEN
            tanh_f := - 2042;
        ELSIF x =- 6471 THEN
            tanh_f := - 2042;
        ELSIF x =- 6470 THEN
            tanh_f := - 2042;
        ELSIF x =- 6469 THEN
            tanh_f := - 2042;
        ELSIF x =- 6468 THEN
            tanh_f := - 2042;
        ELSIF x =- 6467 THEN
            tanh_f := - 2042;
        ELSIF x =- 6466 THEN
            tanh_f := - 2042;
        ELSIF x =- 6465 THEN
            tanh_f := - 2042;
        ELSIF x =- 6464 THEN
            tanh_f := - 2042;
        ELSIF x =- 6463 THEN
            tanh_f := - 2042;
        ELSIF x =- 6462 THEN
            tanh_f := - 2042;
        ELSIF x =- 6461 THEN
            tanh_f := - 2042;
        ELSIF x =- 6460 THEN
            tanh_f := - 2042;
        ELSIF x =- 6459 THEN
            tanh_f := - 2042;
        ELSIF x =- 6458 THEN
            tanh_f := - 2042;
        ELSIF x =- 6457 THEN
            tanh_f := - 2042;
        ELSIF x =- 6456 THEN
            tanh_f := - 2042;
        ELSIF x =- 6455 THEN
            tanh_f := - 2042;
        ELSIF x =- 6454 THEN
            tanh_f := - 2042;
        ELSIF x =- 6453 THEN
            tanh_f := - 2042;
        ELSIF x =- 6452 THEN
            tanh_f := - 2042;
        ELSIF x =- 6451 THEN
            tanh_f := - 2042;
        ELSIF x =- 6450 THEN
            tanh_f := - 2042;
        ELSIF x =- 6449 THEN
            tanh_f := - 2042;
        ELSIF x =- 6448 THEN
            tanh_f := - 2042;
        ELSIF x =- 6447 THEN
            tanh_f := - 2042;
        ELSIF x =- 6446 THEN
            tanh_f := - 2042;
        ELSIF x =- 6445 THEN
            tanh_f := - 2042;
        ELSIF x =- 6444 THEN
            tanh_f := - 2042;
        ELSIF x =- 6443 THEN
            tanh_f := - 2042;
        ELSIF x =- 6442 THEN
            tanh_f := - 2042;
        ELSIF x =- 6441 THEN
            tanh_f := - 2042;
        ELSIF x =- 6440 THEN
            tanh_f := - 2042;
        ELSIF x =- 6439 THEN
            tanh_f := - 2042;
        ELSIF x =- 6438 THEN
            tanh_f := - 2042;
        ELSIF x =- 6437 THEN
            tanh_f := - 2042;
        ELSIF x =- 6436 THEN
            tanh_f := - 2042;
        ELSIF x =- 6435 THEN
            tanh_f := - 2042;
        ELSIF x =- 6434 THEN
            tanh_f := - 2042;
        ELSIF x =- 6433 THEN
            tanh_f := - 2042;
        ELSIF x =- 6432 THEN
            tanh_f := - 2042;
        ELSIF x =- 6431 THEN
            tanh_f := - 2042;
        ELSIF x =- 6430 THEN
            tanh_f := - 2042;
        ELSIF x =- 6429 THEN
            tanh_f := - 2042;
        ELSIF x =- 6428 THEN
            tanh_f := - 2042;
        ELSIF x =- 6427 THEN
            tanh_f := - 2042;
        ELSIF x =- 6426 THEN
            tanh_f := - 2042;
        ELSIF x =- 6425 THEN
            tanh_f := - 2042;
        ELSIF x =- 6424 THEN
            tanh_f := - 2042;
        ELSIF x =- 6423 THEN
            tanh_f := - 2042;
        ELSIF x =- 6422 THEN
            tanh_f := - 2042;
        ELSIF x =- 6421 THEN
            tanh_f := - 2042;
        ELSIF x =- 6420 THEN
            tanh_f := - 2042;
        ELSIF x =- 6419 THEN
            tanh_f := - 2042;
        ELSIF x =- 6418 THEN
            tanh_f := - 2042;
        ELSIF x =- 6417 THEN
            tanh_f := - 2042;
        ELSIF x =- 6416 THEN
            tanh_f := - 2042;
        ELSIF x =- 6415 THEN
            tanh_f := - 2042;
        ELSIF x =- 6414 THEN
            tanh_f := - 2042;
        ELSIF x =- 6413 THEN
            tanh_f := - 2042;
        ELSIF x =- 6412 THEN
            tanh_f := - 2042;
        ELSIF x =- 6411 THEN
            tanh_f := - 2042;
        ELSIF x =- 6410 THEN
            tanh_f := - 2042;
        ELSIF x =- 6409 THEN
            tanh_f := - 2042;
        ELSIF x =- 6408 THEN
            tanh_f := - 2042;
        ELSIF x =- 6407 THEN
            tanh_f := - 2042;
        ELSIF x =- 6406 THEN
            tanh_f := - 2042;
        ELSIF x =- 6405 THEN
            tanh_f := - 2042;
        ELSIF x =- 6404 THEN
            tanh_f := - 2042;
        ELSIF x =- 6403 THEN
            tanh_f := - 2042;
        ELSIF x =- 6402 THEN
            tanh_f := - 2042;
        ELSIF x =- 6401 THEN
            tanh_f := - 2042;
        ELSIF x =- 6400 THEN
            tanh_f := - 2042;
        ELSIF x =- 6399 THEN
            tanh_f := - 2040;
        ELSIF x =- 6398 THEN
            tanh_f := - 2040;
        ELSIF x =- 6397 THEN
            tanh_f := - 2040;
        ELSIF x =- 6396 THEN
            tanh_f := - 2040;
        ELSIF x =- 6395 THEN
            tanh_f := - 2040;
        ELSIF x =- 6394 THEN
            tanh_f := - 2040;
        ELSIF x =- 6393 THEN
            tanh_f := - 2040;
        ELSIF x =- 6392 THEN
            tanh_f := - 2040;
        ELSIF x =- 6391 THEN
            tanh_f := - 2040;
        ELSIF x =- 6390 THEN
            tanh_f := - 2040;
        ELSIF x =- 6389 THEN
            tanh_f := - 2040;
        ELSIF x =- 6388 THEN
            tanh_f := - 2040;
        ELSIF x =- 6387 THEN
            tanh_f := - 2040;
        ELSIF x =- 6386 THEN
            tanh_f := - 2040;
        ELSIF x =- 6385 THEN
            tanh_f := - 2040;
        ELSIF x =- 6384 THEN
            tanh_f := - 2040;
        ELSIF x =- 6383 THEN
            tanh_f := - 2040;
        ELSIF x =- 6382 THEN
            tanh_f := - 2040;
        ELSIF x =- 6381 THEN
            tanh_f := - 2040;
        ELSIF x =- 6380 THEN
            tanh_f := - 2040;
        ELSIF x =- 6379 THEN
            tanh_f := - 2040;
        ELSIF x =- 6378 THEN
            tanh_f := - 2040;
        ELSIF x =- 6377 THEN
            tanh_f := - 2040;
        ELSIF x =- 6376 THEN
            tanh_f := - 2040;
        ELSIF x =- 6375 THEN
            tanh_f := - 2040;
        ELSIF x =- 6374 THEN
            tanh_f := - 2040;
        ELSIF x =- 6373 THEN
            tanh_f := - 2040;
        ELSIF x =- 6372 THEN
            tanh_f := - 2040;
        ELSIF x =- 6371 THEN
            tanh_f := - 2040;
        ELSIF x =- 6370 THEN
            tanh_f := - 2040;
        ELSIF x =- 6369 THEN
            tanh_f := - 2040;
        ELSIF x =- 6368 THEN
            tanh_f := - 2040;
        ELSIF x =- 6367 THEN
            tanh_f := - 2040;
        ELSIF x =- 6366 THEN
            tanh_f := - 2040;
        ELSIF x =- 6365 THEN
            tanh_f := - 2040;
        ELSIF x =- 6364 THEN
            tanh_f := - 2040;
        ELSIF x =- 6363 THEN
            tanh_f := - 2040;
        ELSIF x =- 6362 THEN
            tanh_f := - 2040;
        ELSIF x =- 6361 THEN
            tanh_f := - 2040;
        ELSIF x =- 6360 THEN
            tanh_f := - 2040;
        ELSIF x =- 6359 THEN
            tanh_f := - 2040;
        ELSIF x =- 6358 THEN
            tanh_f := - 2040;
        ELSIF x =- 6357 THEN
            tanh_f := - 2040;
        ELSIF x =- 6356 THEN
            tanh_f := - 2040;
        ELSIF x =- 6355 THEN
            tanh_f := - 2040;
        ELSIF x =- 6354 THEN
            tanh_f := - 2040;
        ELSIF x =- 6353 THEN
            tanh_f := - 2040;
        ELSIF x =- 6352 THEN
            tanh_f := - 2040;
        ELSIF x =- 6351 THEN
            tanh_f := - 2040;
        ELSIF x =- 6350 THEN
            tanh_f := - 2040;
        ELSIF x =- 6349 THEN
            tanh_f := - 2040;
        ELSIF x =- 6348 THEN
            tanh_f := - 2040;
        ELSIF x =- 6347 THEN
            tanh_f := - 2040;
        ELSIF x =- 6346 THEN
            tanh_f := - 2040;
        ELSIF x =- 6345 THEN
            tanh_f := - 2040;
        ELSIF x =- 6344 THEN
            tanh_f := - 2040;
        ELSIF x =- 6343 THEN
            tanh_f := - 2040;
        ELSIF x =- 6342 THEN
            tanh_f := - 2040;
        ELSIF x =- 6341 THEN
            tanh_f := - 2040;
        ELSIF x =- 6340 THEN
            tanh_f := - 2040;
        ELSIF x =- 6339 THEN
            tanh_f := - 2040;
        ELSIF x =- 6338 THEN
            tanh_f := - 2040;
        ELSIF x =- 6337 THEN
            tanh_f := - 2040;
        ELSIF x =- 6336 THEN
            tanh_f := - 2040;
        ELSIF x =- 6335 THEN
            tanh_f := - 2040;
        ELSIF x =- 6334 THEN
            tanh_f := - 2040;
        ELSIF x =- 6333 THEN
            tanh_f := - 2040;
        ELSIF x =- 6332 THEN
            tanh_f := - 2040;
        ELSIF x =- 6331 THEN
            tanh_f := - 2040;
        ELSIF x =- 6330 THEN
            tanh_f := - 2040;
        ELSIF x =- 6329 THEN
            tanh_f := - 2040;
        ELSIF x =- 6328 THEN
            tanh_f := - 2040;
        ELSIF x =- 6327 THEN
            tanh_f := - 2040;
        ELSIF x =- 6326 THEN
            tanh_f := - 2040;
        ELSIF x =- 6325 THEN
            tanh_f := - 2040;
        ELSIF x =- 6324 THEN
            tanh_f := - 2040;
        ELSIF x =- 6323 THEN
            tanh_f := - 2040;
        ELSIF x =- 6322 THEN
            tanh_f := - 2040;
        ELSIF x =- 6321 THEN
            tanh_f := - 2040;
        ELSIF x =- 6320 THEN
            tanh_f := - 2040;
        ELSIF x =- 6319 THEN
            tanh_f := - 2040;
        ELSIF x =- 6318 THEN
            tanh_f := - 2040;
        ELSIF x =- 6317 THEN
            tanh_f := - 2040;
        ELSIF x =- 6316 THEN
            tanh_f := - 2040;
        ELSIF x =- 6315 THEN
            tanh_f := - 2040;
        ELSIF x =- 6314 THEN
            tanh_f := - 2040;
        ELSIF x =- 6313 THEN
            tanh_f := - 2040;
        ELSIF x =- 6312 THEN
            tanh_f := - 2040;
        ELSIF x =- 6311 THEN
            tanh_f := - 2040;
        ELSIF x =- 6310 THEN
            tanh_f := - 2040;
        ELSIF x =- 6309 THEN
            tanh_f := - 2040;
        ELSIF x =- 6308 THEN
            tanh_f := - 2040;
        ELSIF x =- 6307 THEN
            tanh_f := - 2040;
        ELSIF x =- 6306 THEN
            tanh_f := - 2040;
        ELSIF x =- 6305 THEN
            tanh_f := - 2040;
        ELSIF x =- 6304 THEN
            tanh_f := - 2040;
        ELSIF x =- 6303 THEN
            tanh_f := - 2040;
        ELSIF x =- 6302 THEN
            tanh_f := - 2040;
        ELSIF x =- 6301 THEN
            tanh_f := - 2040;
        ELSIF x =- 6300 THEN
            tanh_f := - 2040;
        ELSIF x =- 6299 THEN
            tanh_f := - 2040;
        ELSIF x =- 6298 THEN
            tanh_f := - 2040;
        ELSIF x =- 6297 THEN
            tanh_f := - 2040;
        ELSIF x =- 6296 THEN
            tanh_f := - 2040;
        ELSIF x =- 6295 THEN
            tanh_f := - 2040;
        ELSIF x =- 6294 THEN
            tanh_f := - 2040;
        ELSIF x =- 6293 THEN
            tanh_f := - 2040;
        ELSIF x =- 6292 THEN
            tanh_f := - 2040;
        ELSIF x =- 6291 THEN
            tanh_f := - 2040;
        ELSIF x =- 6290 THEN
            tanh_f := - 2040;
        ELSIF x =- 6289 THEN
            tanh_f := - 2040;
        ELSIF x =- 6288 THEN
            tanh_f := - 2040;
        ELSIF x =- 6287 THEN
            tanh_f := - 2040;
        ELSIF x =- 6286 THEN
            tanh_f := - 2040;
        ELSIF x =- 6285 THEN
            tanh_f := - 2040;
        ELSIF x =- 6284 THEN
            tanh_f := - 2040;
        ELSIF x =- 6283 THEN
            tanh_f := - 2040;
        ELSIF x =- 6282 THEN
            tanh_f := - 2040;
        ELSIF x =- 6281 THEN
            tanh_f := - 2040;
        ELSIF x =- 6280 THEN
            tanh_f := - 2040;
        ELSIF x =- 6279 THEN
            tanh_f := - 2040;
        ELSIF x =- 6278 THEN
            tanh_f := - 2040;
        ELSIF x =- 6277 THEN
            tanh_f := - 2040;
        ELSIF x =- 6276 THEN
            tanh_f := - 2040;
        ELSIF x =- 6275 THEN
            tanh_f := - 2040;
        ELSIF x =- 6274 THEN
            tanh_f := - 2040;
        ELSIF x =- 6273 THEN
            tanh_f := - 2040;
        ELSIF x =- 6272 THEN
            tanh_f := - 2040;
        ELSIF x =- 6271 THEN
            tanh_f := - 2040;
        ELSIF x =- 6270 THEN
            tanh_f := - 2040;
        ELSIF x =- 6269 THEN
            tanh_f := - 2040;
        ELSIF x =- 6268 THEN
            tanh_f := - 2040;
        ELSIF x =- 6267 THEN
            tanh_f := - 2040;
        ELSIF x =- 6266 THEN
            tanh_f := - 2040;
        ELSIF x =- 6265 THEN
            tanh_f := - 2040;
        ELSIF x =- 6264 THEN
            tanh_f := - 2040;
        ELSIF x =- 6263 THEN
            tanh_f := - 2040;
        ELSIF x =- 6262 THEN
            tanh_f := - 2040;
        ELSIF x =- 6261 THEN
            tanh_f := - 2040;
        ELSIF x =- 6260 THEN
            tanh_f := - 2040;
        ELSIF x =- 6259 THEN
            tanh_f := - 2040;
        ELSIF x =- 6258 THEN
            tanh_f := - 2040;
        ELSIF x =- 6257 THEN
            tanh_f := - 2040;
        ELSIF x =- 6256 THEN
            tanh_f := - 2040;
        ELSIF x =- 6255 THEN
            tanh_f := - 2040;
        ELSIF x =- 6254 THEN
            tanh_f := - 2040;
        ELSIF x =- 6253 THEN
            tanh_f := - 2040;
        ELSIF x =- 6252 THEN
            tanh_f := - 2040;
        ELSIF x =- 6251 THEN
            tanh_f := - 2040;
        ELSIF x =- 6250 THEN
            tanh_f := - 2040;
        ELSIF x =- 6249 THEN
            tanh_f := - 2040;
        ELSIF x =- 6248 THEN
            tanh_f := - 2040;
        ELSIF x =- 6247 THEN
            tanh_f := - 2040;
        ELSIF x =- 6246 THEN
            tanh_f := - 2040;
        ELSIF x =- 6245 THEN
            tanh_f := - 2040;
        ELSIF x =- 6244 THEN
            tanh_f := - 2040;
        ELSIF x =- 6243 THEN
            tanh_f := - 2040;
        ELSIF x =- 6242 THEN
            tanh_f := - 2040;
        ELSIF x =- 6241 THEN
            tanh_f := - 2040;
        ELSIF x =- 6240 THEN
            tanh_f := - 2040;
        ELSIF x =- 6239 THEN
            tanh_f := - 2040;
        ELSIF x =- 6238 THEN
            tanh_f := - 2040;
        ELSIF x =- 6237 THEN
            tanh_f := - 2040;
        ELSIF x =- 6236 THEN
            tanh_f := - 2040;
        ELSIF x =- 6235 THEN
            tanh_f := - 2040;
        ELSIF x =- 6234 THEN
            tanh_f := - 2040;
        ELSIF x =- 6233 THEN
            tanh_f := - 2040;
        ELSIF x =- 6232 THEN
            tanh_f := - 2040;
        ELSIF x =- 6231 THEN
            tanh_f := - 2040;
        ELSIF x =- 6230 THEN
            tanh_f := - 2040;
        ELSIF x =- 6229 THEN
            tanh_f := - 2040;
        ELSIF x =- 6228 THEN
            tanh_f := - 2040;
        ELSIF x =- 6227 THEN
            tanh_f := - 2040;
        ELSIF x =- 6226 THEN
            tanh_f := - 2040;
        ELSIF x =- 6225 THEN
            tanh_f := - 2040;
        ELSIF x =- 6224 THEN
            tanh_f := - 2040;
        ELSIF x =- 6223 THEN
            tanh_f := - 2040;
        ELSIF x =- 6222 THEN
            tanh_f := - 2040;
        ELSIF x =- 6221 THEN
            tanh_f := - 2040;
        ELSIF x =- 6220 THEN
            tanh_f := - 2040;
        ELSIF x =- 6219 THEN
            tanh_f := - 2040;
        ELSIF x =- 6218 THEN
            tanh_f := - 2040;
        ELSIF x =- 6217 THEN
            tanh_f := - 2040;
        ELSIF x =- 6216 THEN
            tanh_f := - 2040;
        ELSIF x =- 6215 THEN
            tanh_f := - 2040;
        ELSIF x =- 6214 THEN
            tanh_f := - 2040;
        ELSIF x =- 6213 THEN
            tanh_f := - 2040;
        ELSIF x =- 6212 THEN
            tanh_f := - 2040;
        ELSIF x =- 6211 THEN
            tanh_f := - 2040;
        ELSIF x =- 6210 THEN
            tanh_f := - 2040;
        ELSIF x =- 6209 THEN
            tanh_f := - 2040;
        ELSIF x =- 6208 THEN
            tanh_f := - 2040;
        ELSIF x =- 6207 THEN
            tanh_f := - 2040;
        ELSIF x =- 6206 THEN
            tanh_f := - 2040;
        ELSIF x =- 6205 THEN
            tanh_f := - 2040;
        ELSIF x =- 6204 THEN
            tanh_f := - 2040;
        ELSIF x =- 6203 THEN
            tanh_f := - 2040;
        ELSIF x =- 6202 THEN
            tanh_f := - 2040;
        ELSIF x =- 6201 THEN
            tanh_f := - 2040;
        ELSIF x =- 6200 THEN
            tanh_f := - 2040;
        ELSIF x =- 6199 THEN
            tanh_f := - 2040;
        ELSIF x =- 6198 THEN
            tanh_f := - 2040;
        ELSIF x =- 6197 THEN
            tanh_f := - 2040;
        ELSIF x =- 6196 THEN
            tanh_f := - 2040;
        ELSIF x =- 6195 THEN
            tanh_f := - 2040;
        ELSIF x =- 6194 THEN
            tanh_f := - 2040;
        ELSIF x =- 6193 THEN
            tanh_f := - 2040;
        ELSIF x =- 6192 THEN
            tanh_f := - 2040;
        ELSIF x =- 6191 THEN
            tanh_f := - 2040;
        ELSIF x =- 6190 THEN
            tanh_f := - 2040;
        ELSIF x =- 6189 THEN
            tanh_f := - 2040;
        ELSIF x =- 6188 THEN
            tanh_f := - 2040;
        ELSIF x =- 6187 THEN
            tanh_f := - 2040;
        ELSIF x =- 6186 THEN
            tanh_f := - 2040;
        ELSIF x =- 6185 THEN
            tanh_f := - 2040;
        ELSIF x =- 6184 THEN
            tanh_f := - 2040;
        ELSIF x =- 6183 THEN
            tanh_f := - 2040;
        ELSIF x =- 6182 THEN
            tanh_f := - 2040;
        ELSIF x =- 6181 THEN
            tanh_f := - 2040;
        ELSIF x =- 6180 THEN
            tanh_f := - 2040;
        ELSIF x =- 6179 THEN
            tanh_f := - 2040;
        ELSIF x =- 6178 THEN
            tanh_f := - 2040;
        ELSIF x =- 6177 THEN
            tanh_f := - 2040;
        ELSIF x =- 6176 THEN
            tanh_f := - 2040;
        ELSIF x =- 6175 THEN
            tanh_f := - 2040;
        ELSIF x =- 6174 THEN
            tanh_f := - 2040;
        ELSIF x =- 6173 THEN
            tanh_f := - 2040;
        ELSIF x =- 6172 THEN
            tanh_f := - 2040;
        ELSIF x =- 6171 THEN
            tanh_f := - 2040;
        ELSIF x =- 6170 THEN
            tanh_f := - 2040;
        ELSIF x =- 6169 THEN
            tanh_f := - 2040;
        ELSIF x =- 6168 THEN
            tanh_f := - 2040;
        ELSIF x =- 6167 THEN
            tanh_f := - 2040;
        ELSIF x =- 6166 THEN
            tanh_f := - 2040;
        ELSIF x =- 6165 THEN
            tanh_f := - 2040;
        ELSIF x =- 6164 THEN
            tanh_f := - 2040;
        ELSIF x =- 6163 THEN
            tanh_f := - 2040;
        ELSIF x =- 6162 THEN
            tanh_f := - 2040;
        ELSIF x =- 6161 THEN
            tanh_f := - 2040;
        ELSIF x =- 6160 THEN
            tanh_f := - 2040;
        ELSIF x =- 6159 THEN
            tanh_f := - 2040;
        ELSIF x =- 6158 THEN
            tanh_f := - 2040;
        ELSIF x =- 6157 THEN
            tanh_f := - 2040;
        ELSIF x =- 6156 THEN
            tanh_f := - 2040;
        ELSIF x =- 6155 THEN
            tanh_f := - 2040;
        ELSIF x =- 6154 THEN
            tanh_f := - 2040;
        ELSIF x =- 6153 THEN
            tanh_f := - 2040;
        ELSIF x =- 6152 THEN
            tanh_f := - 2040;
        ELSIF x =- 6151 THEN
            tanh_f := - 2040;
        ELSIF x =- 6150 THEN
            tanh_f := - 2040;
        ELSIF x =- 6149 THEN
            tanh_f := - 2040;
        ELSIF x =- 6148 THEN
            tanh_f := - 2040;
        ELSIF x =- 6147 THEN
            tanh_f := - 2040;
        ELSIF x =- 6146 THEN
            tanh_f := - 2040;
        ELSIF x =- 6145 THEN
            tanh_f := - 2040;
        ELSIF x =- 6144 THEN
            tanh_f := - 2040;
        ELSIF x =- 6143 THEN
            tanh_f := - 2036;
        ELSIF x =- 6142 THEN
            tanh_f := - 2036;
        ELSIF x =- 6141 THEN
            tanh_f := - 2036;
        ELSIF x =- 6140 THEN
            tanh_f := - 2036;
        ELSIF x =- 6139 THEN
            tanh_f := - 2036;
        ELSIF x =- 6138 THEN
            tanh_f := - 2036;
        ELSIF x =- 6137 THEN
            tanh_f := - 2036;
        ELSIF x =- 6136 THEN
            tanh_f := - 2036;
        ELSIF x =- 6135 THEN
            tanh_f := - 2036;
        ELSIF x =- 6134 THEN
            tanh_f := - 2036;
        ELSIF x =- 6133 THEN
            tanh_f := - 2036;
        ELSIF x =- 6132 THEN
            tanh_f := - 2036;
        ELSIF x =- 6131 THEN
            tanh_f := - 2036;
        ELSIF x =- 6130 THEN
            tanh_f := - 2036;
        ELSIF x =- 6129 THEN
            tanh_f := - 2036;
        ELSIF x =- 6128 THEN
            tanh_f := - 2036;
        ELSIF x =- 6127 THEN
            tanh_f := - 2036;
        ELSIF x =- 6126 THEN
            tanh_f := - 2036;
        ELSIF x =- 6125 THEN
            tanh_f := - 2036;
        ELSIF x =- 6124 THEN
            tanh_f := - 2036;
        ELSIF x =- 6123 THEN
            tanh_f := - 2036;
        ELSIF x =- 6122 THEN
            tanh_f := - 2036;
        ELSIF x =- 6121 THEN
            tanh_f := - 2036;
        ELSIF x =- 6120 THEN
            tanh_f := - 2036;
        ELSIF x =- 6119 THEN
            tanh_f := - 2036;
        ELSIF x =- 6118 THEN
            tanh_f := - 2036;
        ELSIF x =- 6117 THEN
            tanh_f := - 2036;
        ELSIF x =- 6116 THEN
            tanh_f := - 2036;
        ELSIF x =- 6115 THEN
            tanh_f := - 2036;
        ELSIF x =- 6114 THEN
            tanh_f := - 2036;
        ELSIF x =- 6113 THEN
            tanh_f := - 2036;
        ELSIF x =- 6112 THEN
            tanh_f := - 2036;
        ELSIF x =- 6111 THEN
            tanh_f := - 2036;
        ELSIF x =- 6110 THEN
            tanh_f := - 2036;
        ELSIF x =- 6109 THEN
            tanh_f := - 2036;
        ELSIF x =- 6108 THEN
            tanh_f := - 2036;
        ELSIF x =- 6107 THEN
            tanh_f := - 2036;
        ELSIF x =- 6106 THEN
            tanh_f := - 2036;
        ELSIF x =- 6105 THEN
            tanh_f := - 2036;
        ELSIF x =- 6104 THEN
            tanh_f := - 2036;
        ELSIF x =- 6103 THEN
            tanh_f := - 2036;
        ELSIF x =- 6102 THEN
            tanh_f := - 2036;
        ELSIF x =- 6101 THEN
            tanh_f := - 2036;
        ELSIF x =- 6100 THEN
            tanh_f := - 2036;
        ELSIF x =- 6099 THEN
            tanh_f := - 2036;
        ELSIF x =- 6098 THEN
            tanh_f := - 2036;
        ELSIF x =- 6097 THEN
            tanh_f := - 2036;
        ELSIF x =- 6096 THEN
            tanh_f := - 2036;
        ELSIF x =- 6095 THEN
            tanh_f := - 2036;
        ELSIF x =- 6094 THEN
            tanh_f := - 2036;
        ELSIF x =- 6093 THEN
            tanh_f := - 2036;
        ELSIF x =- 6092 THEN
            tanh_f := - 2036;
        ELSIF x =- 6091 THEN
            tanh_f := - 2036;
        ELSIF x =- 6090 THEN
            tanh_f := - 2036;
        ELSIF x =- 6089 THEN
            tanh_f := - 2036;
        ELSIF x =- 6088 THEN
            tanh_f := - 2036;
        ELSIF x =- 6087 THEN
            tanh_f := - 2036;
        ELSIF x =- 6086 THEN
            tanh_f := - 2036;
        ELSIF x =- 6085 THEN
            tanh_f := - 2036;
        ELSIF x =- 6084 THEN
            tanh_f := - 2036;
        ELSIF x =- 6083 THEN
            tanh_f := - 2036;
        ELSIF x =- 6082 THEN
            tanh_f := - 2036;
        ELSIF x =- 6081 THEN
            tanh_f := - 2036;
        ELSIF x =- 6080 THEN
            tanh_f := - 2036;
        ELSIF x =- 6079 THEN
            tanh_f := - 2036;
        ELSIF x =- 6078 THEN
            tanh_f := - 2036;
        ELSIF x =- 6077 THEN
            tanh_f := - 2036;
        ELSIF x =- 6076 THEN
            tanh_f := - 2036;
        ELSIF x =- 6075 THEN
            tanh_f := - 2036;
        ELSIF x =- 6074 THEN
            tanh_f := - 2036;
        ELSIF x =- 6073 THEN
            tanh_f := - 2036;
        ELSIF x =- 6072 THEN
            tanh_f := - 2036;
        ELSIF x =- 6071 THEN
            tanh_f := - 2036;
        ELSIF x =- 6070 THEN
            tanh_f := - 2036;
        ELSIF x =- 6069 THEN
            tanh_f := - 2036;
        ELSIF x =- 6068 THEN
            tanh_f := - 2036;
        ELSIF x =- 6067 THEN
            tanh_f := - 2036;
        ELSIF x =- 6066 THEN
            tanh_f := - 2036;
        ELSIF x =- 6065 THEN
            tanh_f := - 2036;
        ELSIF x =- 6064 THEN
            tanh_f := - 2036;
        ELSIF x =- 6063 THEN
            tanh_f := - 2036;
        ELSIF x =- 6062 THEN
            tanh_f := - 2036;
        ELSIF x =- 6061 THEN
            tanh_f := - 2036;
        ELSIF x =- 6060 THEN
            tanh_f := - 2036;
        ELSIF x =- 6059 THEN
            tanh_f := - 2036;
        ELSIF x =- 6058 THEN
            tanh_f := - 2036;
        ELSIF x =- 6057 THEN
            tanh_f := - 2036;
        ELSIF x =- 6056 THEN
            tanh_f := - 2036;
        ELSIF x =- 6055 THEN
            tanh_f := - 2036;
        ELSIF x =- 6054 THEN
            tanh_f := - 2036;
        ELSIF x =- 6053 THEN
            tanh_f := - 2036;
        ELSIF x =- 6052 THEN
            tanh_f := - 2036;
        ELSIF x =- 6051 THEN
            tanh_f := - 2036;
        ELSIF x =- 6050 THEN
            tanh_f := - 2036;
        ELSIF x =- 6049 THEN
            tanh_f := - 2036;
        ELSIF x =- 6048 THEN
            tanh_f := - 2036;
        ELSIF x =- 6047 THEN
            tanh_f := - 2036;
        ELSIF x =- 6046 THEN
            tanh_f := - 2036;
        ELSIF x =- 6045 THEN
            tanh_f := - 2036;
        ELSIF x =- 6044 THEN
            tanh_f := - 2036;
        ELSIF x =- 6043 THEN
            tanh_f := - 2036;
        ELSIF x =- 6042 THEN
            tanh_f := - 2036;
        ELSIF x =- 6041 THEN
            tanh_f := - 2036;
        ELSIF x =- 6040 THEN
            tanh_f := - 2036;
        ELSIF x =- 6039 THEN
            tanh_f := - 2036;
        ELSIF x =- 6038 THEN
            tanh_f := - 2036;
        ELSIF x =- 6037 THEN
            tanh_f := - 2036;
        ELSIF x =- 6036 THEN
            tanh_f := - 2036;
        ELSIF x =- 6035 THEN
            tanh_f := - 2036;
        ELSIF x =- 6034 THEN
            tanh_f := - 2036;
        ELSIF x =- 6033 THEN
            tanh_f := - 2036;
        ELSIF x =- 6032 THEN
            tanh_f := - 2036;
        ELSIF x =- 6031 THEN
            tanh_f := - 2036;
        ELSIF x =- 6030 THEN
            tanh_f := - 2036;
        ELSIF x =- 6029 THEN
            tanh_f := - 2036;
        ELSIF x =- 6028 THEN
            tanh_f := - 2036;
        ELSIF x =- 6027 THEN
            tanh_f := - 2036;
        ELSIF x =- 6026 THEN
            tanh_f := - 2036;
        ELSIF x =- 6025 THEN
            tanh_f := - 2036;
        ELSIF x =- 6024 THEN
            tanh_f := - 2036;
        ELSIF x =- 6023 THEN
            tanh_f := - 2036;
        ELSIF x =- 6022 THEN
            tanh_f := - 2036;
        ELSIF x =- 6021 THEN
            tanh_f := - 2036;
        ELSIF x =- 6020 THEN
            tanh_f := - 2036;
        ELSIF x =- 6019 THEN
            tanh_f := - 2036;
        ELSIF x =- 6018 THEN
            tanh_f := - 2036;
        ELSIF x =- 6017 THEN
            tanh_f := - 2036;
        ELSIF x =- 6016 THEN
            tanh_f := - 2036;
        ELSIF x =- 6015 THEN
            tanh_f := - 2036;
        ELSIF x =- 6014 THEN
            tanh_f := - 2036;
        ELSIF x =- 6013 THEN
            tanh_f := - 2036;
        ELSIF x =- 6012 THEN
            tanh_f := - 2036;
        ELSIF x =- 6011 THEN
            tanh_f := - 2036;
        ELSIF x =- 6010 THEN
            tanh_f := - 2036;
        ELSIF x =- 6009 THEN
            tanh_f := - 2036;
        ELSIF x =- 6008 THEN
            tanh_f := - 2036;
        ELSIF x =- 6007 THEN
            tanh_f := - 2036;
        ELSIF x =- 6006 THEN
            tanh_f := - 2036;
        ELSIF x =- 6005 THEN
            tanh_f := - 2036;
        ELSIF x =- 6004 THEN
            tanh_f := - 2036;
        ELSIF x =- 6003 THEN
            tanh_f := - 2036;
        ELSIF x =- 6002 THEN
            tanh_f := - 2036;
        ELSIF x =- 6001 THEN
            tanh_f := - 2036;
        ELSIF x =- 6000 THEN
            tanh_f := - 2036;
        ELSIF x =- 5999 THEN
            tanh_f := - 2036;
        ELSIF x =- 5998 THEN
            tanh_f := - 2036;
        ELSIF x =- 5997 THEN
            tanh_f := - 2036;
        ELSIF x =- 5996 THEN
            tanh_f := - 2036;
        ELSIF x =- 5995 THEN
            tanh_f := - 2036;
        ELSIF x =- 5994 THEN
            tanh_f := - 2036;
        ELSIF x =- 5993 THEN
            tanh_f := - 2036;
        ELSIF x =- 5992 THEN
            tanh_f := - 2036;
        ELSIF x =- 5991 THEN
            tanh_f := - 2036;
        ELSIF x =- 5990 THEN
            tanh_f := - 2036;
        ELSIF x =- 5989 THEN
            tanh_f := - 2036;
        ELSIF x =- 5988 THEN
            tanh_f := - 2036;
        ELSIF x =- 5987 THEN
            tanh_f := - 2036;
        ELSIF x =- 5986 THEN
            tanh_f := - 2036;
        ELSIF x =- 5985 THEN
            tanh_f := - 2036;
        ELSIF x =- 5984 THEN
            tanh_f := - 2036;
        ELSIF x =- 5983 THEN
            tanh_f := - 2036;
        ELSIF x =- 5982 THEN
            tanh_f := - 2036;
        ELSIF x =- 5981 THEN
            tanh_f := - 2036;
        ELSIF x =- 5980 THEN
            tanh_f := - 2036;
        ELSIF x =- 5979 THEN
            tanh_f := - 2036;
        ELSIF x =- 5978 THEN
            tanh_f := - 2036;
        ELSIF x =- 5977 THEN
            tanh_f := - 2036;
        ELSIF x =- 5976 THEN
            tanh_f := - 2036;
        ELSIF x =- 5975 THEN
            tanh_f := - 2036;
        ELSIF x =- 5974 THEN
            tanh_f := - 2036;
        ELSIF x =- 5973 THEN
            tanh_f := - 2036;
        ELSIF x =- 5972 THEN
            tanh_f := - 2036;
        ELSIF x =- 5971 THEN
            tanh_f := - 2036;
        ELSIF x =- 5970 THEN
            tanh_f := - 2036;
        ELSIF x =- 5969 THEN
            tanh_f := - 2036;
        ELSIF x =- 5968 THEN
            tanh_f := - 2036;
        ELSIF x =- 5967 THEN
            tanh_f := - 2036;
        ELSIF x =- 5966 THEN
            tanh_f := - 2036;
        ELSIF x =- 5965 THEN
            tanh_f := - 2036;
        ELSIF x =- 5964 THEN
            tanh_f := - 2036;
        ELSIF x =- 5963 THEN
            tanh_f := - 2036;
        ELSIF x =- 5962 THEN
            tanh_f := - 2036;
        ELSIF x =- 5961 THEN
            tanh_f := - 2036;
        ELSIF x =- 5960 THEN
            tanh_f := - 2036;
        ELSIF x =- 5959 THEN
            tanh_f := - 2036;
        ELSIF x =- 5958 THEN
            tanh_f := - 2036;
        ELSIF x =- 5957 THEN
            tanh_f := - 2036;
        ELSIF x =- 5956 THEN
            tanh_f := - 2036;
        ELSIF x =- 5955 THEN
            tanh_f := - 2036;
        ELSIF x =- 5954 THEN
            tanh_f := - 2036;
        ELSIF x =- 5953 THEN
            tanh_f := - 2036;
        ELSIF x =- 5952 THEN
            tanh_f := - 2036;
        ELSIF x =- 5951 THEN
            tanh_f := - 2036;
        ELSIF x =- 5950 THEN
            tanh_f := - 2036;
        ELSIF x =- 5949 THEN
            tanh_f := - 2036;
        ELSIF x =- 5948 THEN
            tanh_f := - 2036;
        ELSIF x =- 5947 THEN
            tanh_f := - 2036;
        ELSIF x =- 5946 THEN
            tanh_f := - 2036;
        ELSIF x =- 5945 THEN
            tanh_f := - 2036;
        ELSIF x =- 5944 THEN
            tanh_f := - 2036;
        ELSIF x =- 5943 THEN
            tanh_f := - 2036;
        ELSIF x =- 5942 THEN
            tanh_f := - 2036;
        ELSIF x =- 5941 THEN
            tanh_f := - 2036;
        ELSIF x =- 5940 THEN
            tanh_f := - 2036;
        ELSIF x =- 5939 THEN
            tanh_f := - 2036;
        ELSIF x =- 5938 THEN
            tanh_f := - 2036;
        ELSIF x =- 5937 THEN
            tanh_f := - 2036;
        ELSIF x =- 5936 THEN
            tanh_f := - 2036;
        ELSIF x =- 5935 THEN
            tanh_f := - 2036;
        ELSIF x =- 5934 THEN
            tanh_f := - 2036;
        ELSIF x =- 5933 THEN
            tanh_f := - 2036;
        ELSIF x =- 5932 THEN
            tanh_f := - 2036;
        ELSIF x =- 5931 THEN
            tanh_f := - 2036;
        ELSIF x =- 5930 THEN
            tanh_f := - 2036;
        ELSIF x =- 5929 THEN
            tanh_f := - 2036;
        ELSIF x =- 5928 THEN
            tanh_f := - 2036;
        ELSIF x =- 5927 THEN
            tanh_f := - 2036;
        ELSIF x =- 5926 THEN
            tanh_f := - 2036;
        ELSIF x =- 5925 THEN
            tanh_f := - 2036;
        ELSIF x =- 5924 THEN
            tanh_f := - 2036;
        ELSIF x =- 5923 THEN
            tanh_f := - 2036;
        ELSIF x =- 5922 THEN
            tanh_f := - 2036;
        ELSIF x =- 5921 THEN
            tanh_f := - 2036;
        ELSIF x =- 5920 THEN
            tanh_f := - 2036;
        ELSIF x =- 5919 THEN
            tanh_f := - 2036;
        ELSIF x =- 5918 THEN
            tanh_f := - 2036;
        ELSIF x =- 5917 THEN
            tanh_f := - 2036;
        ELSIF x =- 5916 THEN
            tanh_f := - 2036;
        ELSIF x =- 5915 THEN
            tanh_f := - 2036;
        ELSIF x =- 5914 THEN
            tanh_f := - 2036;
        ELSIF x =- 5913 THEN
            tanh_f := - 2036;
        ELSIF x =- 5912 THEN
            tanh_f := - 2036;
        ELSIF x =- 5911 THEN
            tanh_f := - 2036;
        ELSIF x =- 5910 THEN
            tanh_f := - 2036;
        ELSIF x =- 5909 THEN
            tanh_f := - 2036;
        ELSIF x =- 5908 THEN
            tanh_f := - 2036;
        ELSIF x =- 5907 THEN
            tanh_f := - 2036;
        ELSIF x =- 5906 THEN
            tanh_f := - 2036;
        ELSIF x =- 5905 THEN
            tanh_f := - 2036;
        ELSIF x =- 5904 THEN
            tanh_f := - 2036;
        ELSIF x =- 5903 THEN
            tanh_f := - 2036;
        ELSIF x =- 5902 THEN
            tanh_f := - 2036;
        ELSIF x =- 5901 THEN
            tanh_f := - 2036;
        ELSIF x =- 5900 THEN
            tanh_f := - 2036;
        ELSIF x =- 5899 THEN
            tanh_f := - 2036;
        ELSIF x =- 5898 THEN
            tanh_f := - 2036;
        ELSIF x =- 5897 THEN
            tanh_f := - 2036;
        ELSIF x =- 5896 THEN
            tanh_f := - 2036;
        ELSIF x =- 5895 THEN
            tanh_f := - 2036;
        ELSIF x =- 5894 THEN
            tanh_f := - 2036;
        ELSIF x =- 5893 THEN
            tanh_f := - 2036;
        ELSIF x =- 5892 THEN
            tanh_f := - 2036;
        ELSIF x =- 5891 THEN
            tanh_f := - 2036;
        ELSIF x =- 5890 THEN
            tanh_f := - 2036;
        ELSIF x =- 5889 THEN
            tanh_f := - 2036;
        ELSIF x =- 5888 THEN
            tanh_f := - 2036;
        ELSIF x =- 5887 THEN
            tanh_f := - 2036;
        ELSIF x =- 5886 THEN
            tanh_f := - 2036;
        ELSIF x =- 5885 THEN
            tanh_f := - 2036;
        ELSIF x =- 5884 THEN
            tanh_f := - 2036;
        ELSIF x =- 5883 THEN
            tanh_f := - 2036;
        ELSIF x =- 5882 THEN
            tanh_f := - 2036;
        ELSIF x =- 5881 THEN
            tanh_f := - 2036;
        ELSIF x =- 5880 THEN
            tanh_f := - 2036;
        ELSIF x =- 5879 THEN
            tanh_f := - 2036;
        ELSIF x =- 5878 THEN
            tanh_f := - 2036;
        ELSIF x =- 5877 THEN
            tanh_f := - 2036;
        ELSIF x =- 5876 THEN
            tanh_f := - 2036;
        ELSIF x =- 5875 THEN
            tanh_f := - 2036;
        ELSIF x =- 5874 THEN
            tanh_f := - 2036;
        ELSIF x =- 5873 THEN
            tanh_f := - 2036;
        ELSIF x =- 5872 THEN
            tanh_f := - 2036;
        ELSIF x =- 5871 THEN
            tanh_f := - 2036;
        ELSIF x =- 5870 THEN
            tanh_f := - 2036;
        ELSIF x =- 5869 THEN
            tanh_f := - 2036;
        ELSIF x =- 5868 THEN
            tanh_f := - 2036;
        ELSIF x =- 5867 THEN
            tanh_f := - 2036;
        ELSIF x =- 5866 THEN
            tanh_f := - 2036;
        ELSIF x =- 5865 THEN
            tanh_f := - 2036;
        ELSIF x =- 5864 THEN
            tanh_f := - 2036;
        ELSIF x =- 5863 THEN
            tanh_f := - 2036;
        ELSIF x =- 5862 THEN
            tanh_f := - 2036;
        ELSIF x =- 5861 THEN
            tanh_f := - 2036;
        ELSIF x =- 5860 THEN
            tanh_f := - 2036;
        ELSIF x =- 5859 THEN
            tanh_f := - 2035;
        ELSIF x =- 5858 THEN
            tanh_f := - 2035;
        ELSIF x =- 5857 THEN
            tanh_f := - 2035;
        ELSIF x =- 5856 THEN
            tanh_f := - 2035;
        ELSIF x =- 5855 THEN
            tanh_f := - 2035;
        ELSIF x =- 5854 THEN
            tanh_f := - 2035;
        ELSIF x =- 5853 THEN
            tanh_f := - 2035;
        ELSIF x =- 5852 THEN
            tanh_f := - 2035;
        ELSIF x =- 5851 THEN
            tanh_f := - 2035;
        ELSIF x =- 5850 THEN
            tanh_f := - 2035;
        ELSIF x =- 5849 THEN
            tanh_f := - 2035;
        ELSIF x =- 5848 THEN
            tanh_f := - 2035;
        ELSIF x =- 5847 THEN
            tanh_f := - 2035;
        ELSIF x =- 5846 THEN
            tanh_f := - 2035;
        ELSIF x =- 5845 THEN
            tanh_f := - 2035;
        ELSIF x =- 5844 THEN
            tanh_f := - 2035;
        ELSIF x =- 5843 THEN
            tanh_f := - 2035;
        ELSIF x =- 5842 THEN
            tanh_f := - 2035;
        ELSIF x =- 5841 THEN
            tanh_f := - 2035;
        ELSIF x =- 5840 THEN
            tanh_f := - 2035;
        ELSIF x =- 5839 THEN
            tanh_f := - 2035;
        ELSIF x =- 5838 THEN
            tanh_f := - 2035;
        ELSIF x =- 5837 THEN
            tanh_f := - 2035;
        ELSIF x =- 5836 THEN
            tanh_f := - 2035;
        ELSIF x =- 5835 THEN
            tanh_f := - 2035;
        ELSIF x =- 5834 THEN
            tanh_f := - 2035;
        ELSIF x =- 5833 THEN
            tanh_f := - 2035;
        ELSIF x =- 5832 THEN
            tanh_f := - 2035;
        ELSIF x =- 5831 THEN
            tanh_f := - 2035;
        ELSIF x =- 5830 THEN
            tanh_f := - 2035;
        ELSIF x =- 5829 THEN
            tanh_f := - 2035;
        ELSIF x =- 5828 THEN
            tanh_f := - 2035;
        ELSIF x =- 5827 THEN
            tanh_f := - 2035;
        ELSIF x =- 5826 THEN
            tanh_f := - 2035;
        ELSIF x =- 5825 THEN
            tanh_f := - 2035;
        ELSIF x =- 5824 THEN
            tanh_f := - 2035;
        ELSIF x =- 5823 THEN
            tanh_f := - 2035;
        ELSIF x =- 5822 THEN
            tanh_f := - 2035;
        ELSIF x =- 5821 THEN
            tanh_f := - 2035;
        ELSIF x =- 5820 THEN
            tanh_f := - 2035;
        ELSIF x =- 5819 THEN
            tanh_f := - 2035;
        ELSIF x =- 5818 THEN
            tanh_f := - 2035;
        ELSIF x =- 5817 THEN
            tanh_f := - 2035;
        ELSIF x =- 5816 THEN
            tanh_f := - 2035;
        ELSIF x =- 5815 THEN
            tanh_f := - 2035;
        ELSIF x =- 5814 THEN
            tanh_f := - 2035;
        ELSIF x =- 5813 THEN
            tanh_f := - 2035;
        ELSIF x =- 5812 THEN
            tanh_f := - 2035;
        ELSIF x =- 5811 THEN
            tanh_f := - 2035;
        ELSIF x =- 5810 THEN
            tanh_f := - 2035;
        ELSIF x =- 5809 THEN
            tanh_f := - 2035;
        ELSIF x =- 5808 THEN
            tanh_f := - 2035;
        ELSIF x =- 5807 THEN
            tanh_f := - 2035;
        ELSIF x =- 5806 THEN
            tanh_f := - 2035;
        ELSIF x =- 5805 THEN
            tanh_f := - 2035;
        ELSIF x =- 5804 THEN
            tanh_f := - 2035;
        ELSIF x =- 5803 THEN
            tanh_f := - 2035;
        ELSIF x =- 5802 THEN
            tanh_f := - 2034;
        ELSIF x =- 5801 THEN
            tanh_f := - 2034;
        ELSIF x =- 5800 THEN
            tanh_f := - 2034;
        ELSIF x =- 5799 THEN
            tanh_f := - 2034;
        ELSIF x =- 5798 THEN
            tanh_f := - 2034;
        ELSIF x =- 5797 THEN
            tanh_f := - 2034;
        ELSIF x =- 5796 THEN
            tanh_f := - 2034;
        ELSIF x =- 5795 THEN
            tanh_f := - 2034;
        ELSIF x =- 5794 THEN
            tanh_f := - 2034;
        ELSIF x =- 5793 THEN
            tanh_f := - 2034;
        ELSIF x =- 5792 THEN
            tanh_f := - 2034;
        ELSIF x =- 5791 THEN
            tanh_f := - 2034;
        ELSIF x =- 5790 THEN
            tanh_f := - 2034;
        ELSIF x =- 5789 THEN
            tanh_f := - 2034;
        ELSIF x =- 5788 THEN
            tanh_f := - 2034;
        ELSIF x =- 5787 THEN
            tanh_f := - 2034;
        ELSIF x =- 5786 THEN
            tanh_f := - 2034;
        ELSIF x =- 5785 THEN
            tanh_f := - 2034;
        ELSIF x =- 5784 THEN
            tanh_f := - 2034;
        ELSIF x =- 5783 THEN
            tanh_f := - 2034;
        ELSIF x =- 5782 THEN
            tanh_f := - 2034;
        ELSIF x =- 5781 THEN
            tanh_f := - 2034;
        ELSIF x =- 5780 THEN
            tanh_f := - 2034;
        ELSIF x =- 5779 THEN
            tanh_f := - 2034;
        ELSIF x =- 5778 THEN
            tanh_f := - 2034;
        ELSIF x =- 5777 THEN
            tanh_f := - 2034;
        ELSIF x =- 5776 THEN
            tanh_f := - 2034;
        ELSIF x =- 5775 THEN
            tanh_f := - 2034;
        ELSIF x =- 5774 THEN
            tanh_f := - 2034;
        ELSIF x =- 5773 THEN
            tanh_f := - 2034;
        ELSIF x =- 5772 THEN
            tanh_f := - 2034;
        ELSIF x =- 5771 THEN
            tanh_f := - 2034;
        ELSIF x =- 5770 THEN
            tanh_f := - 2034;
        ELSIF x =- 5769 THEN
            tanh_f := - 2034;
        ELSIF x =- 5768 THEN
            tanh_f := - 2034;
        ELSIF x =- 5767 THEN
            tanh_f := - 2034;
        ELSIF x =- 5766 THEN
            tanh_f := - 2034;
        ELSIF x =- 5765 THEN
            tanh_f := - 2034;
        ELSIF x =- 5764 THEN
            tanh_f := - 2034;
        ELSIF x =- 5763 THEN
            tanh_f := - 2034;
        ELSIF x =- 5762 THEN
            tanh_f := - 2034;
        ELSIF x =- 5761 THEN
            tanh_f := - 2034;
        ELSIF x =- 5760 THEN
            tanh_f := - 2034;
        ELSIF x =- 5759 THEN
            tanh_f := - 2034;
        ELSIF x =- 5758 THEN
            tanh_f := - 2034;
        ELSIF x =- 5757 THEN
            tanh_f := - 2034;
        ELSIF x =- 5756 THEN
            tanh_f := - 2034;
        ELSIF x =- 5755 THEN
            tanh_f := - 2034;
        ELSIF x =- 5754 THEN
            tanh_f := - 2034;
        ELSIF x =- 5753 THEN
            tanh_f := - 2034;
        ELSIF x =- 5752 THEN
            tanh_f := - 2034;
        ELSIF x =- 5751 THEN
            tanh_f := - 2034;
        ELSIF x =- 5750 THEN
            tanh_f := - 2034;
        ELSIF x =- 5749 THEN
            tanh_f := - 2034;
        ELSIF x =- 5748 THEN
            tanh_f := - 2034;
        ELSIF x =- 5747 THEN
            tanh_f := - 2034;
        ELSIF x =- 5746 THEN
            tanh_f := - 2034;
        ELSIF x =- 5745 THEN
            tanh_f := - 2033;
        ELSIF x =- 5744 THEN
            tanh_f := - 2033;
        ELSIF x =- 5743 THEN
            tanh_f := - 2033;
        ELSIF x =- 5742 THEN
            tanh_f := - 2033;
        ELSIF x =- 5741 THEN
            tanh_f := - 2033;
        ELSIF x =- 5740 THEN
            tanh_f := - 2033;
        ELSIF x =- 5739 THEN
            tanh_f := - 2033;
        ELSIF x =- 5738 THEN
            tanh_f := - 2033;
        ELSIF x =- 5737 THEN
            tanh_f := - 2033;
        ELSIF x =- 5736 THEN
            tanh_f := - 2033;
        ELSIF x =- 5735 THEN
            tanh_f := - 2033;
        ELSIF x =- 5734 THEN
            tanh_f := - 2033;
        ELSIF x =- 5733 THEN
            tanh_f := - 2033;
        ELSIF x =- 5732 THEN
            tanh_f := - 2033;
        ELSIF x =- 5731 THEN
            tanh_f := - 2033;
        ELSIF x =- 5730 THEN
            tanh_f := - 2033;
        ELSIF x =- 5729 THEN
            tanh_f := - 2033;
        ELSIF x =- 5728 THEN
            tanh_f := - 2033;
        ELSIF x =- 5727 THEN
            tanh_f := - 2033;
        ELSIF x =- 5726 THEN
            tanh_f := - 2033;
        ELSIF x =- 5725 THEN
            tanh_f := - 2033;
        ELSIF x =- 5724 THEN
            tanh_f := - 2033;
        ELSIF x =- 5723 THEN
            tanh_f := - 2033;
        ELSIF x =- 5722 THEN
            tanh_f := - 2033;
        ELSIF x =- 5721 THEN
            tanh_f := - 2033;
        ELSIF x =- 5720 THEN
            tanh_f := - 2033;
        ELSIF x =- 5719 THEN
            tanh_f := - 2033;
        ELSIF x =- 5718 THEN
            tanh_f := - 2033;
        ELSIF x =- 5717 THEN
            tanh_f := - 2033;
        ELSIF x =- 5716 THEN
            tanh_f := - 2033;
        ELSIF x =- 5715 THEN
            tanh_f := - 2033;
        ELSIF x =- 5714 THEN
            tanh_f := - 2033;
        ELSIF x =- 5713 THEN
            tanh_f := - 2033;
        ELSIF x =- 5712 THEN
            tanh_f := - 2033;
        ELSIF x =- 5711 THEN
            tanh_f := - 2033;
        ELSIF x =- 5710 THEN
            tanh_f := - 2033;
        ELSIF x =- 5709 THEN
            tanh_f := - 2033;
        ELSIF x =- 5708 THEN
            tanh_f := - 2033;
        ELSIF x =- 5707 THEN
            tanh_f := - 2033;
        ELSIF x =- 5706 THEN
            tanh_f := - 2033;
        ELSIF x =- 5705 THEN
            tanh_f := - 2033;
        ELSIF x =- 5704 THEN
            tanh_f := - 2033;
        ELSIF x =- 5703 THEN
            tanh_f := - 2033;
        ELSIF x =- 5702 THEN
            tanh_f := - 2033;
        ELSIF x =- 5701 THEN
            tanh_f := - 2033;
        ELSIF x =- 5700 THEN
            tanh_f := - 2033;
        ELSIF x =- 5699 THEN
            tanh_f := - 2033;
        ELSIF x =- 5698 THEN
            tanh_f := - 2033;
        ELSIF x =- 5697 THEN
            tanh_f := - 2033;
        ELSIF x =- 5696 THEN
            tanh_f := - 2033;
        ELSIF x =- 5695 THEN
            tanh_f := - 2033;
        ELSIF x =- 5694 THEN
            tanh_f := - 2033;
        ELSIF x =- 5693 THEN
            tanh_f := - 2033;
        ELSIF x =- 5692 THEN
            tanh_f := - 2033;
        ELSIF x =- 5691 THEN
            tanh_f := - 2033;
        ELSIF x =- 5690 THEN
            tanh_f := - 2033;
        ELSIF x =- 5689 THEN
            tanh_f := - 2033;
        ELSIF x =- 5688 THEN
            tanh_f := - 2032;
        ELSIF x =- 5687 THEN
            tanh_f := - 2032;
        ELSIF x =- 5686 THEN
            tanh_f := - 2032;
        ELSIF x =- 5685 THEN
            tanh_f := - 2032;
        ELSIF x =- 5684 THEN
            tanh_f := - 2032;
        ELSIF x =- 5683 THEN
            tanh_f := - 2032;
        ELSIF x =- 5682 THEN
            tanh_f := - 2032;
        ELSIF x =- 5681 THEN
            tanh_f := - 2032;
        ELSIF x =- 5680 THEN
            tanh_f := - 2032;
        ELSIF x =- 5679 THEN
            tanh_f := - 2032;
        ELSIF x =- 5678 THEN
            tanh_f := - 2032;
        ELSIF x =- 5677 THEN
            tanh_f := - 2032;
        ELSIF x =- 5676 THEN
            tanh_f := - 2032;
        ELSIF x =- 5675 THEN
            tanh_f := - 2032;
        ELSIF x =- 5674 THEN
            tanh_f := - 2032;
        ELSIF x =- 5673 THEN
            tanh_f := - 2032;
        ELSIF x =- 5672 THEN
            tanh_f := - 2032;
        ELSIF x =- 5671 THEN
            tanh_f := - 2032;
        ELSIF x =- 5670 THEN
            tanh_f := - 2032;
        ELSIF x =- 5669 THEN
            tanh_f := - 2032;
        ELSIF x =- 5668 THEN
            tanh_f := - 2032;
        ELSIF x =- 5667 THEN
            tanh_f := - 2032;
        ELSIF x =- 5666 THEN
            tanh_f := - 2032;
        ELSIF x =- 5665 THEN
            tanh_f := - 2032;
        ELSIF x =- 5664 THEN
            tanh_f := - 2032;
        ELSIF x =- 5663 THEN
            tanh_f := - 2032;
        ELSIF x =- 5662 THEN
            tanh_f := - 2032;
        ELSIF x =- 5661 THEN
            tanh_f := - 2032;
        ELSIF x =- 5660 THEN
            tanh_f := - 2032;
        ELSIF x =- 5659 THEN
            tanh_f := - 2032;
        ELSIF x =- 5658 THEN
            tanh_f := - 2032;
        ELSIF x =- 5657 THEN
            tanh_f := - 2032;
        ELSIF x =- 5656 THEN
            tanh_f := - 2032;
        ELSIF x =- 5655 THEN
            tanh_f := - 2032;
        ELSIF x =- 5654 THEN
            tanh_f := - 2032;
        ELSIF x =- 5653 THEN
            tanh_f := - 2032;
        ELSIF x =- 5652 THEN
            tanh_f := - 2032;
        ELSIF x =- 5651 THEN
            tanh_f := - 2032;
        ELSIF x =- 5650 THEN
            tanh_f := - 2032;
        ELSIF x =- 5649 THEN
            tanh_f := - 2032;
        ELSIF x =- 5648 THEN
            tanh_f := - 2032;
        ELSIF x =- 5647 THEN
            tanh_f := - 2032;
        ELSIF x =- 5646 THEN
            tanh_f := - 2032;
        ELSIF x =- 5645 THEN
            tanh_f := - 2032;
        ELSIF x =- 5644 THEN
            tanh_f := - 2032;
        ELSIF x =- 5643 THEN
            tanh_f := - 2032;
        ELSIF x =- 5642 THEN
            tanh_f := - 2032;
        ELSIF x =- 5641 THEN
            tanh_f := - 2032;
        ELSIF x =- 5640 THEN
            tanh_f := - 2032;
        ELSIF x =- 5639 THEN
            tanh_f := - 2032;
        ELSIF x =- 5638 THEN
            tanh_f := - 2032;
        ELSIF x =- 5637 THEN
            tanh_f := - 2032;
        ELSIF x =- 5636 THEN
            tanh_f := - 2032;
        ELSIF x =- 5635 THEN
            tanh_f := - 2032;
        ELSIF x =- 5634 THEN
            tanh_f := - 2032;
        ELSIF x =- 5633 THEN
            tanh_f := - 2032;
        ELSIF x =- 5632 THEN
            tanh_f := - 2031;
        ELSIF x =- 5631 THEN
            tanh_f := - 2032;
        ELSIF x =- 5630 THEN
            tanh_f := - 2032;
        ELSIF x =- 5629 THEN
            tanh_f := - 2032;
        ELSIF x =- 5628 THEN
            tanh_f := - 2032;
        ELSIF x =- 5627 THEN
            tanh_f := - 2032;
        ELSIF x =- 5626 THEN
            tanh_f := - 2032;
        ELSIF x =- 5625 THEN
            tanh_f := - 2032;
        ELSIF x =- 5624 THEN
            tanh_f := - 2032;
        ELSIF x =- 5623 THEN
            tanh_f := - 2032;
        ELSIF x =- 5622 THEN
            tanh_f := - 2032;
        ELSIF x =- 5621 THEN
            tanh_f := - 2032;
        ELSIF x =- 5620 THEN
            tanh_f := - 2032;
        ELSIF x =- 5619 THEN
            tanh_f := - 2032;
        ELSIF x =- 5618 THEN
            tanh_f := - 2032;
        ELSIF x =- 5617 THEN
            tanh_f := - 2032;
        ELSIF x =- 5616 THEN
            tanh_f := - 2032;
        ELSIF x =- 5615 THEN
            tanh_f := - 2032;
        ELSIF x =- 5614 THEN
            tanh_f := - 2032;
        ELSIF x =- 5613 THEN
            tanh_f := - 2032;
        ELSIF x =- 5612 THEN
            tanh_f := - 2032;
        ELSIF x =- 5611 THEN
            tanh_f := - 2032;
        ELSIF x =- 5610 THEN
            tanh_f := - 2032;
        ELSIF x =- 5609 THEN
            tanh_f := - 2032;
        ELSIF x =- 5608 THEN
            tanh_f := - 2032;
        ELSIF x =- 5607 THEN
            tanh_f := - 2032;
        ELSIF x =- 5606 THEN
            tanh_f := - 2032;
        ELSIF x =- 5605 THEN
            tanh_f := - 2032;
        ELSIF x =- 5604 THEN
            tanh_f := - 2032;
        ELSIF x =- 5603 THEN
            tanh_f := - 2032;
        ELSIF x =- 5602 THEN
            tanh_f := - 2032;
        ELSIF x =- 5601 THEN
            tanh_f := - 2032;
        ELSIF x =- 5600 THEN
            tanh_f := - 2032;
        ELSIF x =- 5599 THEN
            tanh_f := - 2032;
        ELSIF x =- 5598 THEN
            tanh_f := - 2032;
        ELSIF x =- 5597 THEN
            tanh_f := - 2032;
        ELSIF x =- 5596 THEN
            tanh_f := - 2032;
        ELSIF x =- 5595 THEN
            tanh_f := - 2032;
        ELSIF x =- 5594 THEN
            tanh_f := - 2032;
        ELSIF x =- 5593 THEN
            tanh_f := - 2032;
        ELSIF x =- 5592 THEN
            tanh_f := - 2032;
        ELSIF x =- 5591 THEN
            tanh_f := - 2032;
        ELSIF x =- 5590 THEN
            tanh_f := - 2032;
        ELSIF x =- 5589 THEN
            tanh_f := - 2031;
        ELSIF x =- 5588 THEN
            tanh_f := - 2031;
        ELSIF x =- 5587 THEN
            tanh_f := - 2031;
        ELSIF x =- 5586 THEN
            tanh_f := - 2031;
        ELSIF x =- 5585 THEN
            tanh_f := - 2031;
        ELSIF x =- 5584 THEN
            tanh_f := - 2031;
        ELSIF x =- 5583 THEN
            tanh_f := - 2031;
        ELSIF x =- 5582 THEN
            tanh_f := - 2031;
        ELSIF x =- 5581 THEN
            tanh_f := - 2031;
        ELSIF x =- 5580 THEN
            tanh_f := - 2031;
        ELSIF x =- 5579 THEN
            tanh_f := - 2031;
        ELSIF x =- 5578 THEN
            tanh_f := - 2031;
        ELSIF x =- 5577 THEN
            tanh_f := - 2031;
        ELSIF x =- 5576 THEN
            tanh_f := - 2031;
        ELSIF x =- 5575 THEN
            tanh_f := - 2031;
        ELSIF x =- 5574 THEN
            tanh_f := - 2031;
        ELSIF x =- 5573 THEN
            tanh_f := - 2031;
        ELSIF x =- 5572 THEN
            tanh_f := - 2031;
        ELSIF x =- 5571 THEN
            tanh_f := - 2031;
        ELSIF x =- 5570 THEN
            tanh_f := - 2031;
        ELSIF x =- 5569 THEN
            tanh_f := - 2031;
        ELSIF x =- 5568 THEN
            tanh_f := - 2031;
        ELSIF x =- 5567 THEN
            tanh_f := - 2031;
        ELSIF x =- 5566 THEN
            tanh_f := - 2031;
        ELSIF x =- 5565 THEN
            tanh_f := - 2031;
        ELSIF x =- 5564 THEN
            tanh_f := - 2031;
        ELSIF x =- 5563 THEN
            tanh_f := - 2031;
        ELSIF x =- 5562 THEN
            tanh_f := - 2031;
        ELSIF x =- 5561 THEN
            tanh_f := - 2031;
        ELSIF x =- 5560 THEN
            tanh_f := - 2031;
        ELSIF x =- 5559 THEN
            tanh_f := - 2031;
        ELSIF x =- 5558 THEN
            tanh_f := - 2031;
        ELSIF x =- 5557 THEN
            tanh_f := - 2031;
        ELSIF x =- 5556 THEN
            tanh_f := - 2031;
        ELSIF x =- 5555 THEN
            tanh_f := - 2031;
        ELSIF x =- 5554 THEN
            tanh_f := - 2031;
        ELSIF x =- 5553 THEN
            tanh_f := - 2031;
        ELSIF x =- 5552 THEN
            tanh_f := - 2031;
        ELSIF x =- 5551 THEN
            tanh_f := - 2031;
        ELSIF x =- 5550 THEN
            tanh_f := - 2031;
        ELSIF x =- 5549 THEN
            tanh_f := - 2031;
        ELSIF x =- 5548 THEN
            tanh_f := - 2031;
        ELSIF x =- 5547 THEN
            tanh_f := - 2031;
        ELSIF x =- 5546 THEN
            tanh_f := - 2030;
        ELSIF x =- 5545 THEN
            tanh_f := - 2030;
        ELSIF x =- 5544 THEN
            tanh_f := - 2030;
        ELSIF x =- 5543 THEN
            tanh_f := - 2030;
        ELSIF x =- 5542 THEN
            tanh_f := - 2030;
        ELSIF x =- 5541 THEN
            tanh_f := - 2030;
        ELSIF x =- 5540 THEN
            tanh_f := - 2030;
        ELSIF x =- 5539 THEN
            tanh_f := - 2030;
        ELSIF x =- 5538 THEN
            tanh_f := - 2030;
        ELSIF x =- 5537 THEN
            tanh_f := - 2030;
        ELSIF x =- 5536 THEN
            tanh_f := - 2030;
        ELSIF x =- 5535 THEN
            tanh_f := - 2030;
        ELSIF x =- 5534 THEN
            tanh_f := - 2030;
        ELSIF x =- 5533 THEN
            tanh_f := - 2030;
        ELSIF x =- 5532 THEN
            tanh_f := - 2030;
        ELSIF x =- 5531 THEN
            tanh_f := - 2030;
        ELSIF x =- 5530 THEN
            tanh_f := - 2030;
        ELSIF x =- 5529 THEN
            tanh_f := - 2030;
        ELSIF x =- 5528 THEN
            tanh_f := - 2030;
        ELSIF x =- 5527 THEN
            tanh_f := - 2030;
        ELSIF x =- 5526 THEN
            tanh_f := - 2030;
        ELSIF x =- 5525 THEN
            tanh_f := - 2030;
        ELSIF x =- 5524 THEN
            tanh_f := - 2030;
        ELSIF x =- 5523 THEN
            tanh_f := - 2030;
        ELSIF x =- 5522 THEN
            tanh_f := - 2030;
        ELSIF x =- 5521 THEN
            tanh_f := - 2030;
        ELSIF x =- 5520 THEN
            tanh_f := - 2030;
        ELSIF x =- 5519 THEN
            tanh_f := - 2030;
        ELSIF x =- 5518 THEN
            tanh_f := - 2030;
        ELSIF x =- 5517 THEN
            tanh_f := - 2030;
        ELSIF x =- 5516 THEN
            tanh_f := - 2030;
        ELSIF x =- 5515 THEN
            tanh_f := - 2030;
        ELSIF x =- 5514 THEN
            tanh_f := - 2030;
        ELSIF x =- 5513 THEN
            tanh_f := - 2030;
        ELSIF x =- 5512 THEN
            tanh_f := - 2030;
        ELSIF x =- 5511 THEN
            tanh_f := - 2030;
        ELSIF x =- 5510 THEN
            tanh_f := - 2030;
        ELSIF x =- 5509 THEN
            tanh_f := - 2030;
        ELSIF x =- 5508 THEN
            tanh_f := - 2030;
        ELSIF x =- 5507 THEN
            tanh_f := - 2030;
        ELSIF x =- 5506 THEN
            tanh_f := - 2030;
        ELSIF x =- 5505 THEN
            tanh_f := - 2030;
        ELSIF x =- 5504 THEN
            tanh_f := - 2029;
        ELSIF x =- 5503 THEN
            tanh_f := - 2029;
        ELSIF x =- 5502 THEN
            tanh_f := - 2029;
        ELSIF x =- 5501 THEN
            tanh_f := - 2029;
        ELSIF x =- 5500 THEN
            tanh_f := - 2029;
        ELSIF x =- 5499 THEN
            tanh_f := - 2029;
        ELSIF x =- 5498 THEN
            tanh_f := - 2029;
        ELSIF x =- 5497 THEN
            tanh_f := - 2029;
        ELSIF x =- 5496 THEN
            tanh_f := - 2029;
        ELSIF x =- 5495 THEN
            tanh_f := - 2029;
        ELSIF x =- 5494 THEN
            tanh_f := - 2029;
        ELSIF x =- 5493 THEN
            tanh_f := - 2029;
        ELSIF x =- 5492 THEN
            tanh_f := - 2029;
        ELSIF x =- 5491 THEN
            tanh_f := - 2029;
        ELSIF x =- 5490 THEN
            tanh_f := - 2029;
        ELSIF x =- 5489 THEN
            tanh_f := - 2029;
        ELSIF x =- 5488 THEN
            tanh_f := - 2029;
        ELSIF x =- 5487 THEN
            tanh_f := - 2029;
        ELSIF x =- 5486 THEN
            tanh_f := - 2029;
        ELSIF x =- 5485 THEN
            tanh_f := - 2029;
        ELSIF x =- 5484 THEN
            tanh_f := - 2029;
        ELSIF x =- 5483 THEN
            tanh_f := - 2029;
        ELSIF x =- 5482 THEN
            tanh_f := - 2029;
        ELSIF x =- 5481 THEN
            tanh_f := - 2029;
        ELSIF x =- 5480 THEN
            tanh_f := - 2029;
        ELSIF x =- 5479 THEN
            tanh_f := - 2029;
        ELSIF x =- 5478 THEN
            tanh_f := - 2029;
        ELSIF x =- 5477 THEN
            tanh_f := - 2029;
        ELSIF x =- 5476 THEN
            tanh_f := - 2029;
        ELSIF x =- 5475 THEN
            tanh_f := - 2029;
        ELSIF x =- 5474 THEN
            tanh_f := - 2029;
        ELSIF x =- 5473 THEN
            tanh_f := - 2029;
        ELSIF x =- 5472 THEN
            tanh_f := - 2029;
        ELSIF x =- 5471 THEN
            tanh_f := - 2029;
        ELSIF x =- 5470 THEN
            tanh_f := - 2029;
        ELSIF x =- 5469 THEN
            tanh_f := - 2029;
        ELSIF x =- 5468 THEN
            tanh_f := - 2029;
        ELSIF x =- 5467 THEN
            tanh_f := - 2029;
        ELSIF x =- 5466 THEN
            tanh_f := - 2029;
        ELSIF x =- 5465 THEN
            tanh_f := - 2029;
        ELSIF x =- 5464 THEN
            tanh_f := - 2029;
        ELSIF x =- 5463 THEN
            tanh_f := - 2029;
        ELSIF x =- 5462 THEN
            tanh_f := - 2029;
        ELSIF x =- 5461 THEN
            tanh_f := - 2028;
        ELSIF x =- 5460 THEN
            tanh_f := - 2028;
        ELSIF x =- 5459 THEN
            tanh_f := - 2028;
        ELSIF x =- 5458 THEN
            tanh_f := - 2028;
        ELSIF x =- 5457 THEN
            tanh_f := - 2028;
        ELSIF x =- 5456 THEN
            tanh_f := - 2028;
        ELSIF x =- 5455 THEN
            tanh_f := - 2028;
        ELSIF x =- 5454 THEN
            tanh_f := - 2028;
        ELSIF x =- 5453 THEN
            tanh_f := - 2028;
        ELSIF x =- 5452 THEN
            tanh_f := - 2028;
        ELSIF x =- 5451 THEN
            tanh_f := - 2028;
        ELSIF x =- 5450 THEN
            tanh_f := - 2028;
        ELSIF x =- 5449 THEN
            tanh_f := - 2028;
        ELSIF x =- 5448 THEN
            tanh_f := - 2028;
        ELSIF x =- 5447 THEN
            tanh_f := - 2028;
        ELSIF x =- 5446 THEN
            tanh_f := - 2028;
        ELSIF x =- 5445 THEN
            tanh_f := - 2028;
        ELSIF x =- 5444 THEN
            tanh_f := - 2028;
        ELSIF x =- 5443 THEN
            tanh_f := - 2028;
        ELSIF x =- 5442 THEN
            tanh_f := - 2028;
        ELSIF x =- 5441 THEN
            tanh_f := - 2028;
        ELSIF x =- 5440 THEN
            tanh_f := - 2028;
        ELSIF x =- 5439 THEN
            tanh_f := - 2028;
        ELSIF x =- 5438 THEN
            tanh_f := - 2028;
        ELSIF x =- 5437 THEN
            tanh_f := - 2028;
        ELSIF x =- 5436 THEN
            tanh_f := - 2028;
        ELSIF x =- 5435 THEN
            tanh_f := - 2028;
        ELSIF x =- 5434 THEN
            tanh_f := - 2028;
        ELSIF x =- 5433 THEN
            tanh_f := - 2028;
        ELSIF x =- 5432 THEN
            tanh_f := - 2028;
        ELSIF x =- 5431 THEN
            tanh_f := - 2028;
        ELSIF x =- 5430 THEN
            tanh_f := - 2028;
        ELSIF x =- 5429 THEN
            tanh_f := - 2028;
        ELSIF x =- 5428 THEN
            tanh_f := - 2028;
        ELSIF x =- 5427 THEN
            tanh_f := - 2028;
        ELSIF x =- 5426 THEN
            tanh_f := - 2028;
        ELSIF x =- 5425 THEN
            tanh_f := - 2028;
        ELSIF x =- 5424 THEN
            tanh_f := - 2028;
        ELSIF x =- 5423 THEN
            tanh_f := - 2028;
        ELSIF x =- 5422 THEN
            tanh_f := - 2028;
        ELSIF x =- 5421 THEN
            tanh_f := - 2028;
        ELSIF x =- 5420 THEN
            tanh_f := - 2028;
        ELSIF x =- 5419 THEN
            tanh_f := - 2028;
        ELSIF x =- 5418 THEN
            tanh_f := - 2027;
        ELSIF x =- 5417 THEN
            tanh_f := - 2027;
        ELSIF x =- 5416 THEN
            tanh_f := - 2027;
        ELSIF x =- 5415 THEN
            tanh_f := - 2027;
        ELSIF x =- 5414 THEN
            tanh_f := - 2027;
        ELSIF x =- 5413 THEN
            tanh_f := - 2027;
        ELSIF x =- 5412 THEN
            tanh_f := - 2027;
        ELSIF x =- 5411 THEN
            tanh_f := - 2027;
        ELSIF x =- 5410 THEN
            tanh_f := - 2027;
        ELSIF x =- 5409 THEN
            tanh_f := - 2027;
        ELSIF x =- 5408 THEN
            tanh_f := - 2027;
        ELSIF x =- 5407 THEN
            tanh_f := - 2027;
        ELSIF x =- 5406 THEN
            tanh_f := - 2027;
        ELSIF x =- 5405 THEN
            tanh_f := - 2027;
        ELSIF x =- 5404 THEN
            tanh_f := - 2027;
        ELSIF x =- 5403 THEN
            tanh_f := - 2027;
        ELSIF x =- 5402 THEN
            tanh_f := - 2027;
        ELSIF x =- 5401 THEN
            tanh_f := - 2027;
        ELSIF x =- 5400 THEN
            tanh_f := - 2027;
        ELSIF x =- 5399 THEN
            tanh_f := - 2027;
        ELSIF x =- 5398 THEN
            tanh_f := - 2027;
        ELSIF x =- 5397 THEN
            tanh_f := - 2027;
        ELSIF x =- 5396 THEN
            tanh_f := - 2027;
        ELSIF x =- 5395 THEN
            tanh_f := - 2027;
        ELSIF x =- 5394 THEN
            tanh_f := - 2027;
        ELSIF x =- 5393 THEN
            tanh_f := - 2027;
        ELSIF x =- 5392 THEN
            tanh_f := - 2027;
        ELSIF x =- 5391 THEN
            tanh_f := - 2027;
        ELSIF x =- 5390 THEN
            tanh_f := - 2027;
        ELSIF x =- 5389 THEN
            tanh_f := - 2027;
        ELSIF x =- 5388 THEN
            tanh_f := - 2027;
        ELSIF x =- 5387 THEN
            tanh_f := - 2027;
        ELSIF x =- 5386 THEN
            tanh_f := - 2027;
        ELSIF x =- 5385 THEN
            tanh_f := - 2027;
        ELSIF x =- 5384 THEN
            tanh_f := - 2027;
        ELSIF x =- 5383 THEN
            tanh_f := - 2027;
        ELSIF x =- 5382 THEN
            tanh_f := - 2027;
        ELSIF x =- 5381 THEN
            tanh_f := - 2027;
        ELSIF x =- 5380 THEN
            tanh_f := - 2027;
        ELSIF x =- 5379 THEN
            tanh_f := - 2027;
        ELSIF x =- 5378 THEN
            tanh_f := - 2027;
        ELSIF x =- 5377 THEN
            tanh_f := - 2027;
        ELSIF x =- 5376 THEN
            tanh_f := - 2026;
        ELSIF x =- 5375 THEN
            tanh_f := - 2027;
        ELSIF x =- 5374 THEN
            tanh_f := - 2027;
        ELSIF x =- 5373 THEN
            tanh_f := - 2027;
        ELSIF x =- 5372 THEN
            tanh_f := - 2027;
        ELSIF x =- 5371 THEN
            tanh_f := - 2027;
        ELSIF x =- 5370 THEN
            tanh_f := - 2027;
        ELSIF x =- 5369 THEN
            tanh_f := - 2027;
        ELSIF x =- 5368 THEN
            tanh_f := - 2027;
        ELSIF x =- 5367 THEN
            tanh_f := - 2027;
        ELSIF x =- 5366 THEN
            tanh_f := - 2027;
        ELSIF x =- 5365 THEN
            tanh_f := - 2027;
        ELSIF x =- 5364 THEN
            tanh_f := - 2027;
        ELSIF x =- 5363 THEN
            tanh_f := - 2027;
        ELSIF x =- 5362 THEN
            tanh_f := - 2027;
        ELSIF x =- 5361 THEN
            tanh_f := - 2027;
        ELSIF x =- 5360 THEN
            tanh_f := - 2027;
        ELSIF x =- 5359 THEN
            tanh_f := - 2027;
        ELSIF x =- 5358 THEN
            tanh_f := - 2027;
        ELSIF x =- 5357 THEN
            tanh_f := - 2027;
        ELSIF x =- 5356 THEN
            tanh_f := - 2027;
        ELSIF x =- 5355 THEN
            tanh_f := - 2027;
        ELSIF x =- 5354 THEN
            tanh_f := - 2027;
        ELSIF x =- 5353 THEN
            tanh_f := - 2027;
        ELSIF x =- 5352 THEN
            tanh_f := - 2027;
        ELSIF x =- 5351 THEN
            tanh_f := - 2027;
        ELSIF x =- 5350 THEN
            tanh_f := - 2027;
        ELSIF x =- 5349 THEN
            tanh_f := - 2027;
        ELSIF x =- 5348 THEN
            tanh_f := - 2027;
        ELSIF x =- 5347 THEN
            tanh_f := - 2027;
        ELSIF x =- 5346 THEN
            tanh_f := - 2027;
        ELSIF x =- 5345 THEN
            tanh_f := - 2027;
        ELSIF x =- 5344 THEN
            tanh_f := - 2027;
        ELSIF x =- 5343 THEN
            tanh_f := - 2027;
        ELSIF x =- 5342 THEN
            tanh_f := - 2027;
        ELSIF x =- 5341 THEN
            tanh_f := - 2027;
        ELSIF x =- 5340 THEN
            tanh_f := - 2027;
        ELSIF x =- 5339 THEN
            tanh_f := - 2026;
        ELSIF x =- 5338 THEN
            tanh_f := - 2026;
        ELSIF x =- 5337 THEN
            tanh_f := - 2026;
        ELSIF x =- 5336 THEN
            tanh_f := - 2026;
        ELSIF x =- 5335 THEN
            tanh_f := - 2026;
        ELSIF x =- 5334 THEN
            tanh_f := - 2026;
        ELSIF x =- 5333 THEN
            tanh_f := - 2026;
        ELSIF x =- 5332 THEN
            tanh_f := - 2026;
        ELSIF x =- 5331 THEN
            tanh_f := - 2026;
        ELSIF x =- 5330 THEN
            tanh_f := - 2026;
        ELSIF x =- 5329 THEN
            tanh_f := - 2026;
        ELSIF x =- 5328 THEN
            tanh_f := - 2026;
        ELSIF x =- 5327 THEN
            tanh_f := - 2026;
        ELSIF x =- 5326 THEN
            tanh_f := - 2026;
        ELSIF x =- 5325 THEN
            tanh_f := - 2026;
        ELSIF x =- 5324 THEN
            tanh_f := - 2026;
        ELSIF x =- 5323 THEN
            tanh_f := - 2026;
        ELSIF x =- 5322 THEN
            tanh_f := - 2026;
        ELSIF x =- 5321 THEN
            tanh_f := - 2026;
        ELSIF x =- 5320 THEN
            tanh_f := - 2026;
        ELSIF x =- 5319 THEN
            tanh_f := - 2026;
        ELSIF x =- 5318 THEN
            tanh_f := - 2026;
        ELSIF x =- 5317 THEN
            tanh_f := - 2026;
        ELSIF x =- 5316 THEN
            tanh_f := - 2026;
        ELSIF x =- 5315 THEN
            tanh_f := - 2026;
        ELSIF x =- 5314 THEN
            tanh_f := - 2026;
        ELSIF x =- 5313 THEN
            tanh_f := - 2026;
        ELSIF x =- 5312 THEN
            tanh_f := - 2026;
        ELSIF x =- 5311 THEN
            tanh_f := - 2026;
        ELSIF x =- 5310 THEN
            tanh_f := - 2026;
        ELSIF x =- 5309 THEN
            tanh_f := - 2026;
        ELSIF x =- 5308 THEN
            tanh_f := - 2026;
        ELSIF x =- 5307 THEN
            tanh_f := - 2026;
        ELSIF x =- 5306 THEN
            tanh_f := - 2026;
        ELSIF x =- 5305 THEN
            tanh_f := - 2026;
        ELSIF x =- 5304 THEN
            tanh_f := - 2026;
        ELSIF x =- 5303 THEN
            tanh_f := - 2026;
        ELSIF x =- 5302 THEN
            tanh_f := - 2025;
        ELSIF x =- 5301 THEN
            tanh_f := - 2025;
        ELSIF x =- 5300 THEN
            tanh_f := - 2025;
        ELSIF x =- 5299 THEN
            tanh_f := - 2025;
        ELSIF x =- 5298 THEN
            tanh_f := - 2025;
        ELSIF x =- 5297 THEN
            tanh_f := - 2025;
        ELSIF x =- 5296 THEN
            tanh_f := - 2025;
        ELSIF x =- 5295 THEN
            tanh_f := - 2025;
        ELSIF x =- 5294 THEN
            tanh_f := - 2025;
        ELSIF x =- 5293 THEN
            tanh_f := - 2025;
        ELSIF x =- 5292 THEN
            tanh_f := - 2025;
        ELSIF x =- 5291 THEN
            tanh_f := - 2025;
        ELSIF x =- 5290 THEN
            tanh_f := - 2025;
        ELSIF x =- 5289 THEN
            tanh_f := - 2025;
        ELSIF x =- 5288 THEN
            tanh_f := - 2025;
        ELSIF x =- 5287 THEN
            tanh_f := - 2025;
        ELSIF x =- 5286 THEN
            tanh_f := - 2025;
        ELSIF x =- 5285 THEN
            tanh_f := - 2025;
        ELSIF x =- 5284 THEN
            tanh_f := - 2025;
        ELSIF x =- 5283 THEN
            tanh_f := - 2025;
        ELSIF x =- 5282 THEN
            tanh_f := - 2025;
        ELSIF x =- 5281 THEN
            tanh_f := - 2025;
        ELSIF x =- 5280 THEN
            tanh_f := - 2025;
        ELSIF x =- 5279 THEN
            tanh_f := - 2025;
        ELSIF x =- 5278 THEN
            tanh_f := - 2025;
        ELSIF x =- 5277 THEN
            tanh_f := - 2025;
        ELSIF x =- 5276 THEN
            tanh_f := - 2025;
        ELSIF x =- 5275 THEN
            tanh_f := - 2025;
        ELSIF x =- 5274 THEN
            tanh_f := - 2025;
        ELSIF x =- 5273 THEN
            tanh_f := - 2025;
        ELSIF x =- 5272 THEN
            tanh_f := - 2025;
        ELSIF x =- 5271 THEN
            tanh_f := - 2025;
        ELSIF x =- 5270 THEN
            tanh_f := - 2025;
        ELSIF x =- 5269 THEN
            tanh_f := - 2025;
        ELSIF x =- 5268 THEN
            tanh_f := - 2025;
        ELSIF x =- 5267 THEN
            tanh_f := - 2025;
        ELSIF x =- 5266 THEN
            tanh_f := - 2024;
        ELSIF x =- 5265 THEN
            tanh_f := - 2024;
        ELSIF x =- 5264 THEN
            tanh_f := - 2024;
        ELSIF x =- 5263 THEN
            tanh_f := - 2024;
        ELSIF x =- 5262 THEN
            tanh_f := - 2024;
        ELSIF x =- 5261 THEN
            tanh_f := - 2024;
        ELSIF x =- 5260 THEN
            tanh_f := - 2024;
        ELSIF x =- 5259 THEN
            tanh_f := - 2024;
        ELSIF x =- 5258 THEN
            tanh_f := - 2024;
        ELSIF x =- 5257 THEN
            tanh_f := - 2024;
        ELSIF x =- 5256 THEN
            tanh_f := - 2024;
        ELSIF x =- 5255 THEN
            tanh_f := - 2024;
        ELSIF x =- 5254 THEN
            tanh_f := - 2024;
        ELSIF x =- 5253 THEN
            tanh_f := - 2024;
        ELSIF x =- 5252 THEN
            tanh_f := - 2024;
        ELSIF x =- 5251 THEN
            tanh_f := - 2024;
        ELSIF x =- 5250 THEN
            tanh_f := - 2024;
        ELSIF x =- 5249 THEN
            tanh_f := - 2024;
        ELSIF x =- 5248 THEN
            tanh_f := - 2024;
        ELSIF x =- 5247 THEN
            tanh_f := - 2024;
        ELSIF x =- 5246 THEN
            tanh_f := - 2024;
        ELSIF x =- 5245 THEN
            tanh_f := - 2024;
        ELSIF x =- 5244 THEN
            tanh_f := - 2024;
        ELSIF x =- 5243 THEN
            tanh_f := - 2024;
        ELSIF x =- 5242 THEN
            tanh_f := - 2024;
        ELSIF x =- 5241 THEN
            tanh_f := - 2024;
        ELSIF x =- 5240 THEN
            tanh_f := - 2024;
        ELSIF x =- 5239 THEN
            tanh_f := - 2024;
        ELSIF x =- 5238 THEN
            tanh_f := - 2024;
        ELSIF x =- 5237 THEN
            tanh_f := - 2024;
        ELSIF x =- 5236 THEN
            tanh_f := - 2024;
        ELSIF x =- 5235 THEN
            tanh_f := - 2024;
        ELSIF x =- 5234 THEN
            tanh_f := - 2024;
        ELSIF x =- 5233 THEN
            tanh_f := - 2024;
        ELSIF x =- 5232 THEN
            tanh_f := - 2024;
        ELSIF x =- 5231 THEN
            tanh_f := - 2024;
        ELSIF x =- 5230 THEN
            tanh_f := - 2024;
        ELSIF x =- 5229 THEN
            tanh_f := - 2023;
        ELSIF x =- 5228 THEN
            tanh_f := - 2023;
        ELSIF x =- 5227 THEN
            tanh_f := - 2023;
        ELSIF x =- 5226 THEN
            tanh_f := - 2023;
        ELSIF x =- 5225 THEN
            tanh_f := - 2023;
        ELSIF x =- 5224 THEN
            tanh_f := - 2023;
        ELSIF x =- 5223 THEN
            tanh_f := - 2023;
        ELSIF x =- 5222 THEN
            tanh_f := - 2023;
        ELSIF x =- 5221 THEN
            tanh_f := - 2023;
        ELSIF x =- 5220 THEN
            tanh_f := - 2023;
        ELSIF x =- 5219 THEN
            tanh_f := - 2023;
        ELSIF x =- 5218 THEN
            tanh_f := - 2023;
        ELSIF x =- 5217 THEN
            tanh_f := - 2023;
        ELSIF x =- 5216 THEN
            tanh_f := - 2023;
        ELSIF x =- 5215 THEN
            tanh_f := - 2023;
        ELSIF x =- 5214 THEN
            tanh_f := - 2023;
        ELSIF x =- 5213 THEN
            tanh_f := - 2023;
        ELSIF x =- 5212 THEN
            tanh_f := - 2023;
        ELSIF x =- 5211 THEN
            tanh_f := - 2023;
        ELSIF x =- 5210 THEN
            tanh_f := - 2023;
        ELSIF x =- 5209 THEN
            tanh_f := - 2023;
        ELSIF x =- 5208 THEN
            tanh_f := - 2023;
        ELSIF x =- 5207 THEN
            tanh_f := - 2023;
        ELSIF x =- 5206 THEN
            tanh_f := - 2023;
        ELSIF x =- 5205 THEN
            tanh_f := - 2023;
        ELSIF x =- 5204 THEN
            tanh_f := - 2023;
        ELSIF x =- 5203 THEN
            tanh_f := - 2023;
        ELSIF x =- 5202 THEN
            tanh_f := - 2023;
        ELSIF x =- 5201 THEN
            tanh_f := - 2023;
        ELSIF x =- 5200 THEN
            tanh_f := - 2023;
        ELSIF x =- 5199 THEN
            tanh_f := - 2023;
        ELSIF x =- 5198 THEN
            tanh_f := - 2023;
        ELSIF x =- 5197 THEN
            tanh_f := - 2023;
        ELSIF x =- 5196 THEN
            tanh_f := - 2023;
        ELSIF x =- 5195 THEN
            tanh_f := - 2023;
        ELSIF x =- 5194 THEN
            tanh_f := - 2023;
        ELSIF x =- 5193 THEN
            tanh_f := - 2022;
        ELSIF x =- 5192 THEN
            tanh_f := - 2022;
        ELSIF x =- 5191 THEN
            tanh_f := - 2022;
        ELSIF x =- 5190 THEN
            tanh_f := - 2022;
        ELSIF x =- 5189 THEN
            tanh_f := - 2022;
        ELSIF x =- 5188 THEN
            tanh_f := - 2022;
        ELSIF x =- 5187 THEN
            tanh_f := - 2022;
        ELSIF x =- 5186 THEN
            tanh_f := - 2022;
        ELSIF x =- 5185 THEN
            tanh_f := - 2022;
        ELSIF x =- 5184 THEN
            tanh_f := - 2022;
        ELSIF x =- 5183 THEN
            tanh_f := - 2022;
        ELSIF x =- 5182 THEN
            tanh_f := - 2022;
        ELSIF x =- 5181 THEN
            tanh_f := - 2022;
        ELSIF x =- 5180 THEN
            tanh_f := - 2022;
        ELSIF x =- 5179 THEN
            tanh_f := - 2022;
        ELSIF x =- 5178 THEN
            tanh_f := - 2022;
        ELSIF x =- 5177 THEN
            tanh_f := - 2022;
        ELSIF x =- 5176 THEN
            tanh_f := - 2022;
        ELSIF x =- 5175 THEN
            tanh_f := - 2022;
        ELSIF x =- 5174 THEN
            tanh_f := - 2022;
        ELSIF x =- 5173 THEN
            tanh_f := - 2022;
        ELSIF x =- 5172 THEN
            tanh_f := - 2022;
        ELSIF x =- 5171 THEN
            tanh_f := - 2022;
        ELSIF x =- 5170 THEN
            tanh_f := - 2022;
        ELSIF x =- 5169 THEN
            tanh_f := - 2022;
        ELSIF x =- 5168 THEN
            tanh_f := - 2022;
        ELSIF x =- 5167 THEN
            tanh_f := - 2022;
        ELSIF x =- 5166 THEN
            tanh_f := - 2022;
        ELSIF x =- 5165 THEN
            tanh_f := - 2022;
        ELSIF x =- 5164 THEN
            tanh_f := - 2022;
        ELSIF x =- 5163 THEN
            tanh_f := - 2022;
        ELSIF x =- 5162 THEN
            tanh_f := - 2022;
        ELSIF x =- 5161 THEN
            tanh_f := - 2022;
        ELSIF x =- 5160 THEN
            tanh_f := - 2022;
        ELSIF x =- 5159 THEN
            tanh_f := - 2022;
        ELSIF x =- 5158 THEN
            tanh_f := - 2022;
        ELSIF x =- 5157 THEN
            tanh_f := - 2022;
        ELSIF x =- 5156 THEN
            tanh_f := - 2021;
        ELSIF x =- 5155 THEN
            tanh_f := - 2021;
        ELSIF x =- 5154 THEN
            tanh_f := - 2021;
        ELSIF x =- 5153 THEN
            tanh_f := - 2021;
        ELSIF x =- 5152 THEN
            tanh_f := - 2021;
        ELSIF x =- 5151 THEN
            tanh_f := - 2021;
        ELSIF x =- 5150 THEN
            tanh_f := - 2021;
        ELSIF x =- 5149 THEN
            tanh_f := - 2021;
        ELSIF x =- 5148 THEN
            tanh_f := - 2021;
        ELSIF x =- 5147 THEN
            tanh_f := - 2021;
        ELSIF x =- 5146 THEN
            tanh_f := - 2021;
        ELSIF x =- 5145 THEN
            tanh_f := - 2021;
        ELSIF x =- 5144 THEN
            tanh_f := - 2021;
        ELSIF x =- 5143 THEN
            tanh_f := - 2021;
        ELSIF x =- 5142 THEN
            tanh_f := - 2021;
        ELSIF x =- 5141 THEN
            tanh_f := - 2021;
        ELSIF x =- 5140 THEN
            tanh_f := - 2021;
        ELSIF x =- 5139 THEN
            tanh_f := - 2021;
        ELSIF x =- 5138 THEN
            tanh_f := - 2021;
        ELSIF x =- 5137 THEN
            tanh_f := - 2021;
        ELSIF x =- 5136 THEN
            tanh_f := - 2021;
        ELSIF x =- 5135 THEN
            tanh_f := - 2021;
        ELSIF x =- 5134 THEN
            tanh_f := - 2021;
        ELSIF x =- 5133 THEN
            tanh_f := - 2021;
        ELSIF x =- 5132 THEN
            tanh_f := - 2021;
        ELSIF x =- 5131 THEN
            tanh_f := - 2021;
        ELSIF x =- 5130 THEN
            tanh_f := - 2021;
        ELSIF x =- 5129 THEN
            tanh_f := - 2021;
        ELSIF x =- 5128 THEN
            tanh_f := - 2021;
        ELSIF x =- 5127 THEN
            tanh_f := - 2021;
        ELSIF x =- 5126 THEN
            tanh_f := - 2021;
        ELSIF x =- 5125 THEN
            tanh_f := - 2021;
        ELSIF x =- 5124 THEN
            tanh_f := - 2021;
        ELSIF x =- 5123 THEN
            tanh_f := - 2021;
        ELSIF x =- 5122 THEN
            tanh_f := - 2021;
        ELSIF x =- 5121 THEN
            tanh_f := - 2021;
        ELSIF x =- 5120 THEN
            tanh_f := - 2020;
        ELSIF x =- 5119 THEN
            tanh_f := - 2020;
        ELSIF x =- 5118 THEN
            tanh_f := - 2020;
        ELSIF x =- 5117 THEN
            tanh_f := - 2020;
        ELSIF x =- 5116 THEN
            tanh_f := - 2020;
        ELSIF x =- 5115 THEN
            tanh_f := - 2020;
        ELSIF x =- 5114 THEN
            tanh_f := - 2020;
        ELSIF x =- 5113 THEN
            tanh_f := - 2020;
        ELSIF x =- 5112 THEN
            tanh_f := - 2020;
        ELSIF x =- 5111 THEN
            tanh_f := - 2020;
        ELSIF x =- 5110 THEN
            tanh_f := - 2020;
        ELSIF x =- 5109 THEN
            tanh_f := - 2020;
        ELSIF x =- 5108 THEN
            tanh_f := - 2020;
        ELSIF x =- 5107 THEN
            tanh_f := - 2020;
        ELSIF x =- 5106 THEN
            tanh_f := - 2020;
        ELSIF x =- 5105 THEN
            tanh_f := - 2020;
        ELSIF x =- 5104 THEN
            tanh_f := - 2020;
        ELSIF x =- 5103 THEN
            tanh_f := - 2020;
        ELSIF x =- 5102 THEN
            tanh_f := - 2020;
        ELSIF x =- 5101 THEN
            tanh_f := - 2020;
        ELSIF x =- 5100 THEN
            tanh_f := - 2020;
        ELSIF x =- 5099 THEN
            tanh_f := - 2020;
        ELSIF x =- 5098 THEN
            tanh_f := - 2020;
        ELSIF x =- 5097 THEN
            tanh_f := - 2020;
        ELSIF x =- 5096 THEN
            tanh_f := - 2020;
        ELSIF x =- 5095 THEN
            tanh_f := - 2020;
        ELSIF x =- 5094 THEN
            tanh_f := - 2020;
        ELSIF x =- 5093 THEN
            tanh_f := - 2020;
        ELSIF x =- 5092 THEN
            tanh_f := - 2020;
        ELSIF x =- 5091 THEN
            tanh_f := - 2020;
        ELSIF x =- 5090 THEN
            tanh_f := - 2020;
        ELSIF x =- 5089 THEN
            tanh_f := - 2020;
        ELSIF x =- 5088 THEN
            tanh_f := - 2020;
        ELSIF x =- 5087 THEN
            tanh_f := - 2020;
        ELSIF x =- 5086 THEN
            tanh_f := - 2020;
        ELSIF x =- 5085 THEN
            tanh_f := - 2020;
        ELSIF x =- 5084 THEN
            tanh_f := - 2020;
        ELSIF x =- 5083 THEN
            tanh_f := - 2020;
        ELSIF x =- 5082 THEN
            tanh_f := - 2020;
        ELSIF x =- 5081 THEN
            tanh_f := - 2020;
        ELSIF x =- 5080 THEN
            tanh_f := - 2019;
        ELSIF x =- 5079 THEN
            tanh_f := - 2019;
        ELSIF x =- 5078 THEN
            tanh_f := - 2019;
        ELSIF x =- 5077 THEN
            tanh_f := - 2019;
        ELSIF x =- 5076 THEN
            tanh_f := - 2019;
        ELSIF x =- 5075 THEN
            tanh_f := - 2019;
        ELSIF x =- 5074 THEN
            tanh_f := - 2019;
        ELSIF x =- 5073 THEN
            tanh_f := - 2019;
        ELSIF x =- 5072 THEN
            tanh_f := - 2019;
        ELSIF x =- 5071 THEN
            tanh_f := - 2019;
        ELSIF x =- 5070 THEN
            tanh_f := - 2019;
        ELSIF x =- 5069 THEN
            tanh_f := - 2019;
        ELSIF x =- 5068 THEN
            tanh_f := - 2019;
        ELSIF x =- 5067 THEN
            tanh_f := - 2019;
        ELSIF x =- 5066 THEN
            tanh_f := - 2019;
        ELSIF x =- 5065 THEN
            tanh_f := - 2019;
        ELSIF x =- 5064 THEN
            tanh_f := - 2019;
        ELSIF x =- 5063 THEN
            tanh_f := - 2019;
        ELSIF x =- 5062 THEN
            tanh_f := - 2019;
        ELSIF x =- 5061 THEN
            tanh_f := - 2019;
        ELSIF x =- 5060 THEN
            tanh_f := - 2019;
        ELSIF x =- 5059 THEN
            tanh_f := - 2019;
        ELSIF x =- 5058 THEN
            tanh_f := - 2019;
        ELSIF x =- 5057 THEN
            tanh_f := - 2019;
        ELSIF x =- 5056 THEN
            tanh_f := - 2019;
        ELSIF x =- 5055 THEN
            tanh_f := - 2019;
        ELSIF x =- 5054 THEN
            tanh_f := - 2019;
        ELSIF x =- 5053 THEN
            tanh_f := - 2019;
        ELSIF x =- 5052 THEN
            tanh_f := - 2019;
        ELSIF x =- 5051 THEN
            tanh_f := - 2019;
        ELSIF x =- 5050 THEN
            tanh_f := - 2019;
        ELSIF x =- 5049 THEN
            tanh_f := - 2019;
        ELSIF x =- 5048 THEN
            tanh_f := - 2019;
        ELSIF x =- 5047 THEN
            tanh_f := - 2019;
        ELSIF x =- 5046 THEN
            tanh_f := - 2019;
        ELSIF x =- 5045 THEN
            tanh_f := - 2019;
        ELSIF x =- 5044 THEN
            tanh_f := - 2019;
        ELSIF x =- 5043 THEN
            tanh_f := - 2019;
        ELSIF x =- 5042 THEN
            tanh_f := - 2019;
        ELSIF x =- 5041 THEN
            tanh_f := - 2018;
        ELSIF x =- 5040 THEN
            tanh_f := - 2018;
        ELSIF x =- 5039 THEN
            tanh_f := - 2018;
        ELSIF x =- 5038 THEN
            tanh_f := - 2018;
        ELSIF x =- 5037 THEN
            tanh_f := - 2018;
        ELSIF x =- 5036 THEN
            tanh_f := - 2018;
        ELSIF x =- 5035 THEN
            tanh_f := - 2018;
        ELSIF x =- 5034 THEN
            tanh_f := - 2018;
        ELSIF x =- 5033 THEN
            tanh_f := - 2018;
        ELSIF x =- 5032 THEN
            tanh_f := - 2018;
        ELSIF x =- 5031 THEN
            tanh_f := - 2018;
        ELSIF x =- 5030 THEN
            tanh_f := - 2018;
        ELSIF x =- 5029 THEN
            tanh_f := - 2018;
        ELSIF x =- 5028 THEN
            tanh_f := - 2018;
        ELSIF x =- 5027 THEN
            tanh_f := - 2018;
        ELSIF x =- 5026 THEN
            tanh_f := - 2018;
        ELSIF x =- 5025 THEN
            tanh_f := - 2018;
        ELSIF x =- 5024 THEN
            tanh_f := - 2018;
        ELSIF x =- 5023 THEN
            tanh_f := - 2018;
        ELSIF x =- 5022 THEN
            tanh_f := - 2018;
        ELSIF x =- 5021 THEN
            tanh_f := - 2018;
        ELSIF x =- 5020 THEN
            tanh_f := - 2018;
        ELSIF x =- 5019 THEN
            tanh_f := - 2018;
        ELSIF x =- 5018 THEN
            tanh_f := - 2018;
        ELSIF x =- 5017 THEN
            tanh_f := - 2018;
        ELSIF x =- 5016 THEN
            tanh_f := - 2018;
        ELSIF x =- 5015 THEN
            tanh_f := - 2018;
        ELSIF x =- 5014 THEN
            tanh_f := - 2018;
        ELSIF x =- 5013 THEN
            tanh_f := - 2018;
        ELSIF x =- 5012 THEN
            tanh_f := - 2018;
        ELSIF x =- 5011 THEN
            tanh_f := - 2018;
        ELSIF x =- 5010 THEN
            tanh_f := - 2018;
        ELSIF x =- 5009 THEN
            tanh_f := - 2018;
        ELSIF x =- 5008 THEN
            tanh_f := - 2018;
        ELSIF x =- 5007 THEN
            tanh_f := - 2018;
        ELSIF x =- 5006 THEN
            tanh_f := - 2018;
        ELSIF x =- 5005 THEN
            tanh_f := - 2018;
        ELSIF x =- 5004 THEN
            tanh_f := - 2018;
        ELSIF x =- 5003 THEN
            tanh_f := - 2018;
        ELSIF x =- 5002 THEN
            tanh_f := - 2018;
        ELSIF x =- 5001 THEN
            tanh_f := - 2017;
        ELSIF x =- 5000 THEN
            tanh_f := - 2017;
        ELSIF x =- 4999 THEN
            tanh_f := - 2017;
        ELSIF x =- 4998 THEN
            tanh_f := - 2017;
        ELSIF x =- 4997 THEN
            tanh_f := - 2017;
        ELSIF x =- 4996 THEN
            tanh_f := - 2017;
        ELSIF x =- 4995 THEN
            tanh_f := - 2017;
        ELSIF x =- 4994 THEN
            tanh_f := - 2017;
        ELSIF x =- 4993 THEN
            tanh_f := - 2017;
        ELSIF x =- 4992 THEN
            tanh_f := - 2017;
        ELSIF x =- 4991 THEN
            tanh_f := - 2017;
        ELSIF x =- 4990 THEN
            tanh_f := - 2017;
        ELSIF x =- 4989 THEN
            tanh_f := - 2017;
        ELSIF x =- 4988 THEN
            tanh_f := - 2017;
        ELSIF x =- 4987 THEN
            tanh_f := - 2017;
        ELSIF x =- 4986 THEN
            tanh_f := - 2017;
        ELSIF x =- 4985 THEN
            tanh_f := - 2017;
        ELSIF x =- 4984 THEN
            tanh_f := - 2017;
        ELSIF x =- 4983 THEN
            tanh_f := - 2017;
        ELSIF x =- 4982 THEN
            tanh_f := - 2017;
        ELSIF x =- 4981 THEN
            tanh_f := - 2017;
        ELSIF x =- 4980 THEN
            tanh_f := - 2017;
        ELSIF x =- 4979 THEN
            tanh_f := - 2017;
        ELSIF x =- 4978 THEN
            tanh_f := - 2017;
        ELSIF x =- 4977 THEN
            tanh_f := - 2017;
        ELSIF x =- 4976 THEN
            tanh_f := - 2017;
        ELSIF x =- 4975 THEN
            tanh_f := - 2017;
        ELSIF x =- 4974 THEN
            tanh_f := - 2017;
        ELSIF x =- 4973 THEN
            tanh_f := - 2017;
        ELSIF x =- 4972 THEN
            tanh_f := - 2017;
        ELSIF x =- 4971 THEN
            tanh_f := - 2017;
        ELSIF x =- 4970 THEN
            tanh_f := - 2017;
        ELSIF x =- 4969 THEN
            tanh_f := - 2017;
        ELSIF x =- 4968 THEN
            tanh_f := - 2017;
        ELSIF x =- 4967 THEN
            tanh_f := - 2017;
        ELSIF x =- 4966 THEN
            tanh_f := - 2017;
        ELSIF x =- 4965 THEN
            tanh_f := - 2017;
        ELSIF x =- 4964 THEN
            tanh_f := - 2017;
        ELSIF x =- 4963 THEN
            tanh_f := - 2017;
        ELSIF x =- 4962 THEN
            tanh_f := - 2016;
        ELSIF x =- 4961 THEN
            tanh_f := - 2016;
        ELSIF x =- 4960 THEN
            tanh_f := - 2016;
        ELSIF x =- 4959 THEN
            tanh_f := - 2016;
        ELSIF x =- 4958 THEN
            tanh_f := - 2016;
        ELSIF x =- 4957 THEN
            tanh_f := - 2016;
        ELSIF x =- 4956 THEN
            tanh_f := - 2016;
        ELSIF x =- 4955 THEN
            tanh_f := - 2016;
        ELSIF x =- 4954 THEN
            tanh_f := - 2016;
        ELSIF x =- 4953 THEN
            tanh_f := - 2016;
        ELSIF x =- 4952 THEN
            tanh_f := - 2016;
        ELSIF x =- 4951 THEN
            tanh_f := - 2016;
        ELSIF x =- 4950 THEN
            tanh_f := - 2016;
        ELSIF x =- 4949 THEN
            tanh_f := - 2016;
        ELSIF x =- 4948 THEN
            tanh_f := - 2016;
        ELSIF x =- 4947 THEN
            tanh_f := - 2016;
        ELSIF x =- 4946 THEN
            tanh_f := - 2016;
        ELSIF x =- 4945 THEN
            tanh_f := - 2016;
        ELSIF x =- 4944 THEN
            tanh_f := - 2016;
        ELSIF x =- 4943 THEN
            tanh_f := - 2016;
        ELSIF x =- 4942 THEN
            tanh_f := - 2016;
        ELSIF x =- 4941 THEN
            tanh_f := - 2016;
        ELSIF x =- 4940 THEN
            tanh_f := - 2016;
        ELSIF x =- 4939 THEN
            tanh_f := - 2016;
        ELSIF x =- 4938 THEN
            tanh_f := - 2016;
        ELSIF x =- 4937 THEN
            tanh_f := - 2016;
        ELSIF x =- 4936 THEN
            tanh_f := - 2016;
        ELSIF x =- 4935 THEN
            tanh_f := - 2016;
        ELSIF x =- 4934 THEN
            tanh_f := - 2016;
        ELSIF x =- 4933 THEN
            tanh_f := - 2016;
        ELSIF x =- 4932 THEN
            tanh_f := - 2016;
        ELSIF x =- 4931 THEN
            tanh_f := - 2016;
        ELSIF x =- 4930 THEN
            tanh_f := - 2016;
        ELSIF x =- 4929 THEN
            tanh_f := - 2016;
        ELSIF x =- 4928 THEN
            tanh_f := - 2016;
        ELSIF x =- 4927 THEN
            tanh_f := - 2016;
        ELSIF x =- 4926 THEN
            tanh_f := - 2016;
        ELSIF x =- 4925 THEN
            tanh_f := - 2016;
        ELSIF x =- 4924 THEN
            tanh_f := - 2016;
        ELSIF x =- 4923 THEN
            tanh_f := - 2015;
        ELSIF x =- 4922 THEN
            tanh_f := - 2015;
        ELSIF x =- 4921 THEN
            tanh_f := - 2015;
        ELSIF x =- 4920 THEN
            tanh_f := - 2015;
        ELSIF x =- 4919 THEN
            tanh_f := - 2015;
        ELSIF x =- 4918 THEN
            tanh_f := - 2015;
        ELSIF x =- 4917 THEN
            tanh_f := - 2015;
        ELSIF x =- 4916 THEN
            tanh_f := - 2015;
        ELSIF x =- 4915 THEN
            tanh_f := - 2015;
        ELSIF x =- 4914 THEN
            tanh_f := - 2015;
        ELSIF x =- 4913 THEN
            tanh_f := - 2015;
        ELSIF x =- 4912 THEN
            tanh_f := - 2015;
        ELSIF x =- 4911 THEN
            tanh_f := - 2015;
        ELSIF x =- 4910 THEN
            tanh_f := - 2015;
        ELSIF x =- 4909 THEN
            tanh_f := - 2015;
        ELSIF x =- 4908 THEN
            tanh_f := - 2015;
        ELSIF x =- 4907 THEN
            tanh_f := - 2015;
        ELSIF x =- 4906 THEN
            tanh_f := - 2015;
        ELSIF x =- 4905 THEN
            tanh_f := - 2015;
        ELSIF x =- 4904 THEN
            tanh_f := - 2015;
        ELSIF x =- 4903 THEN
            tanh_f := - 2015;
        ELSIF x =- 4902 THEN
            tanh_f := - 2015;
        ELSIF x =- 4901 THEN
            tanh_f := - 2015;
        ELSIF x =- 4900 THEN
            tanh_f := - 2015;
        ELSIF x =- 4899 THEN
            tanh_f := - 2015;
        ELSIF x =- 4898 THEN
            tanh_f := - 2015;
        ELSIF x =- 4897 THEN
            tanh_f := - 2015;
        ELSIF x =- 4896 THEN
            tanh_f := - 2015;
        ELSIF x =- 4895 THEN
            tanh_f := - 2015;
        ELSIF x =- 4894 THEN
            tanh_f := - 2015;
        ELSIF x =- 4893 THEN
            tanh_f := - 2015;
        ELSIF x =- 4892 THEN
            tanh_f := - 2015;
        ELSIF x =- 4891 THEN
            tanh_f := - 2015;
        ELSIF x =- 4890 THEN
            tanh_f := - 2015;
        ELSIF x =- 4889 THEN
            tanh_f := - 2015;
        ELSIF x =- 4888 THEN
            tanh_f := - 2015;
        ELSIF x =- 4887 THEN
            tanh_f := - 2015;
        ELSIF x =- 4886 THEN
            tanh_f := - 2015;
        ELSIF x =- 4885 THEN
            tanh_f := - 2015;
        ELSIF x =- 4884 THEN
            tanh_f := - 2015;
        ELSIF x =- 4883 THEN
            tanh_f := - 2014;
        ELSIF x =- 4882 THEN
            tanh_f := - 2014;
        ELSIF x =- 4881 THEN
            tanh_f := - 2014;
        ELSIF x =- 4880 THEN
            tanh_f := - 2014;
        ELSIF x =- 4879 THEN
            tanh_f := - 2014;
        ELSIF x =- 4878 THEN
            tanh_f := - 2014;
        ELSIF x =- 4877 THEN
            tanh_f := - 2014;
        ELSIF x =- 4876 THEN
            tanh_f := - 2014;
        ELSIF x =- 4875 THEN
            tanh_f := - 2014;
        ELSIF x =- 4874 THEN
            tanh_f := - 2014;
        ELSIF x =- 4873 THEN
            tanh_f := - 2014;
        ELSIF x =- 4872 THEN
            tanh_f := - 2014;
        ELSIF x =- 4871 THEN
            tanh_f := - 2014;
        ELSIF x =- 4870 THEN
            tanh_f := - 2014;
        ELSIF x =- 4869 THEN
            tanh_f := - 2014;
        ELSIF x =- 4868 THEN
            tanh_f := - 2014;
        ELSIF x =- 4867 THEN
            tanh_f := - 2014;
        ELSIF x =- 4866 THEN
            tanh_f := - 2014;
        ELSIF x =- 4865 THEN
            tanh_f := - 2014;
        ELSIF x =- 4864 THEN
            tanh_f := - 2014;
        ELSIF x =- 4863 THEN
            tanh_f := - 2014;
        ELSIF x =- 4862 THEN
            tanh_f := - 2014;
        ELSIF x =- 4861 THEN
            tanh_f := - 2014;
        ELSIF x =- 4860 THEN
            tanh_f := - 2014;
        ELSIF x =- 4859 THEN
            tanh_f := - 2014;
        ELSIF x =- 4858 THEN
            tanh_f := - 2014;
        ELSIF x =- 4857 THEN
            tanh_f := - 2014;
        ELSIF x =- 4856 THEN
            tanh_f := - 2014;
        ELSIF x =- 4855 THEN
            tanh_f := - 2014;
        ELSIF x =- 4854 THEN
            tanh_f := - 2014;
        ELSIF x =- 4853 THEN
            tanh_f := - 2014;
        ELSIF x =- 4852 THEN
            tanh_f := - 2014;
        ELSIF x =- 4851 THEN
            tanh_f := - 2013;
        ELSIF x =- 4850 THEN
            tanh_f := - 2013;
        ELSIF x =- 4849 THEN
            tanh_f := - 2013;
        ELSIF x =- 4848 THEN
            tanh_f := - 2013;
        ELSIF x =- 4847 THEN
            tanh_f := - 2013;
        ELSIF x =- 4846 THEN
            tanh_f := - 2013;
        ELSIF x =- 4845 THEN
            tanh_f := - 2013;
        ELSIF x =- 4844 THEN
            tanh_f := - 2013;
        ELSIF x =- 4843 THEN
            tanh_f := - 2013;
        ELSIF x =- 4842 THEN
            tanh_f := - 2013;
        ELSIF x =- 4841 THEN
            tanh_f := - 2013;
        ELSIF x =- 4840 THEN
            tanh_f := - 2013;
        ELSIF x =- 4839 THEN
            tanh_f := - 2013;
        ELSIF x =- 4838 THEN
            tanh_f := - 2013;
        ELSIF x =- 4837 THEN
            tanh_f := - 2013;
        ELSIF x =- 4836 THEN
            tanh_f := - 2013;
        ELSIF x =- 4835 THEN
            tanh_f := - 2013;
        ELSIF x =- 4834 THEN
            tanh_f := - 2013;
        ELSIF x =- 4833 THEN
            tanh_f := - 2013;
        ELSIF x =- 4832 THEN
            tanh_f := - 2013;
        ELSIF x =- 4831 THEN
            tanh_f := - 2013;
        ELSIF x =- 4830 THEN
            tanh_f := - 2013;
        ELSIF x =- 4829 THEN
            tanh_f := - 2013;
        ELSIF x =- 4828 THEN
            tanh_f := - 2013;
        ELSIF x =- 4827 THEN
            tanh_f := - 2012;
        ELSIF x =- 4826 THEN
            tanh_f := - 2012;
        ELSIF x =- 4825 THEN
            tanh_f := - 2012;
        ELSIF x =- 4824 THEN
            tanh_f := - 2012;
        ELSIF x =- 4823 THEN
            tanh_f := - 2012;
        ELSIF x =- 4822 THEN
            tanh_f := - 2012;
        ELSIF x =- 4821 THEN
            tanh_f := - 2012;
        ELSIF x =- 4820 THEN
            tanh_f := - 2012;
        ELSIF x =- 4819 THEN
            tanh_f := - 2012;
        ELSIF x =- 4818 THEN
            tanh_f := - 2012;
        ELSIF x =- 4817 THEN
            tanh_f := - 2012;
        ELSIF x =- 4816 THEN
            tanh_f := - 2012;
        ELSIF x =- 4815 THEN
            tanh_f := - 2012;
        ELSIF x =- 4814 THEN
            tanh_f := - 2012;
        ELSIF x =- 4813 THEN
            tanh_f := - 2012;
        ELSIF x =- 4812 THEN
            tanh_f := - 2012;
        ELSIF x =- 4811 THEN
            tanh_f := - 2012;
        ELSIF x =- 4810 THEN
            tanh_f := - 2012;
        ELSIF x =- 4809 THEN
            tanh_f := - 2012;
        ELSIF x =- 4808 THEN
            tanh_f := - 2012;
        ELSIF x =- 4807 THEN
            tanh_f := - 2012;
        ELSIF x =- 4806 THEN
            tanh_f := - 2012;
        ELSIF x =- 4805 THEN
            tanh_f := - 2012;
        ELSIF x =- 4804 THEN
            tanh_f := - 2012;
        ELSIF x =- 4803 THEN
            tanh_f := - 2011;
        ELSIF x =- 4802 THEN
            tanh_f := - 2011;
        ELSIF x =- 4801 THEN
            tanh_f := - 2011;
        ELSIF x =- 4800 THEN
            tanh_f := - 2011;
        ELSIF x =- 4799 THEN
            tanh_f := - 2011;
        ELSIF x =- 4798 THEN
            tanh_f := - 2011;
        ELSIF x =- 4797 THEN
            tanh_f := - 2011;
        ELSIF x =- 4796 THEN
            tanh_f := - 2011;
        ELSIF x =- 4795 THEN
            tanh_f := - 2011;
        ELSIF x =- 4794 THEN
            tanh_f := - 2011;
        ELSIF x =- 4793 THEN
            tanh_f := - 2011;
        ELSIF x =- 4792 THEN
            tanh_f := - 2011;
        ELSIF x =- 4791 THEN
            tanh_f := - 2011;
        ELSIF x =- 4790 THEN
            tanh_f := - 2011;
        ELSIF x =- 4789 THEN
            tanh_f := - 2011;
        ELSIF x =- 4788 THEN
            tanh_f := - 2011;
        ELSIF x =- 4787 THEN
            tanh_f := - 2011;
        ELSIF x =- 4786 THEN
            tanh_f := - 2011;
        ELSIF x =- 4785 THEN
            tanh_f := - 2011;
        ELSIF x =- 4784 THEN
            tanh_f := - 2011;
        ELSIF x =- 4783 THEN
            tanh_f := - 2011;
        ELSIF x =- 4782 THEN
            tanh_f := - 2011;
        ELSIF x =- 4781 THEN
            tanh_f := - 2011;
        ELSIF x =- 4780 THEN
            tanh_f := - 2011;
        ELSIF x =- 4779 THEN
            tanh_f := - 2011;
        ELSIF x =- 4778 THEN
            tanh_f := - 2010;
        ELSIF x =- 4777 THEN
            tanh_f := - 2010;
        ELSIF x =- 4776 THEN
            tanh_f := - 2010;
        ELSIF x =- 4775 THEN
            tanh_f := - 2010;
        ELSIF x =- 4774 THEN
            tanh_f := - 2010;
        ELSIF x =- 4773 THEN
            tanh_f := - 2010;
        ELSIF x =- 4772 THEN
            tanh_f := - 2010;
        ELSIF x =- 4771 THEN
            tanh_f := - 2010;
        ELSIF x =- 4770 THEN
            tanh_f := - 2010;
        ELSIF x =- 4769 THEN
            tanh_f := - 2010;
        ELSIF x =- 4768 THEN
            tanh_f := - 2010;
        ELSIF x =- 4767 THEN
            tanh_f := - 2010;
        ELSIF x =- 4766 THEN
            tanh_f := - 2010;
        ELSIF x =- 4765 THEN
            tanh_f := - 2010;
        ELSIF x =- 4764 THEN
            tanh_f := - 2010;
        ELSIF x =- 4763 THEN
            tanh_f := - 2010;
        ELSIF x =- 4762 THEN
            tanh_f := - 2010;
        ELSIF x =- 4761 THEN
            tanh_f := - 2010;
        ELSIF x =- 4760 THEN
            tanh_f := - 2010;
        ELSIF x =- 4759 THEN
            tanh_f := - 2010;
        ELSIF x =- 4758 THEN
            tanh_f := - 2010;
        ELSIF x =- 4757 THEN
            tanh_f := - 2010;
        ELSIF x =- 4756 THEN
            tanh_f := - 2010;
        ELSIF x =- 4755 THEN
            tanh_f := - 2010;
        ELSIF x =- 4754 THEN
            tanh_f := - 2009;
        ELSIF x =- 4753 THEN
            tanh_f := - 2009;
        ELSIF x =- 4752 THEN
            tanh_f := - 2009;
        ELSIF x =- 4751 THEN
            tanh_f := - 2009;
        ELSIF x =- 4750 THEN
            tanh_f := - 2009;
        ELSIF x =- 4749 THEN
            tanh_f := - 2009;
        ELSIF x =- 4748 THEN
            tanh_f := - 2009;
        ELSIF x =- 4747 THEN
            tanh_f := - 2009;
        ELSIF x =- 4746 THEN
            tanh_f := - 2009;
        ELSIF x =- 4745 THEN
            tanh_f := - 2009;
        ELSIF x =- 4744 THEN
            tanh_f := - 2009;
        ELSIF x =- 4743 THEN
            tanh_f := - 2009;
        ELSIF x =- 4742 THEN
            tanh_f := - 2009;
        ELSIF x =- 4741 THEN
            tanh_f := - 2009;
        ELSIF x =- 4740 THEN
            tanh_f := - 2009;
        ELSIF x =- 4739 THEN
            tanh_f := - 2009;
        ELSIF x =- 4738 THEN
            tanh_f := - 2009;
        ELSIF x =- 4737 THEN
            tanh_f := - 2009;
        ELSIF x =- 4736 THEN
            tanh_f := - 2009;
        ELSIF x =- 4735 THEN
            tanh_f := - 2009;
        ELSIF x =- 4734 THEN
            tanh_f := - 2009;
        ELSIF x =- 4733 THEN
            tanh_f := - 2009;
        ELSIF x =- 4732 THEN
            tanh_f := - 2009;
        ELSIF x =- 4731 THEN
            tanh_f := - 2009;
        ELSIF x =- 4730 THEN
            tanh_f := - 2009;
        ELSIF x =- 4729 THEN
            tanh_f := - 2008;
        ELSIF x =- 4728 THEN
            tanh_f := - 2008;
        ELSIF x =- 4727 THEN
            tanh_f := - 2008;
        ELSIF x =- 4726 THEN
            tanh_f := - 2008;
        ELSIF x =- 4725 THEN
            tanh_f := - 2008;
        ELSIF x =- 4724 THEN
            tanh_f := - 2008;
        ELSIF x =- 4723 THEN
            tanh_f := - 2008;
        ELSIF x =- 4722 THEN
            tanh_f := - 2008;
        ELSIF x =- 4721 THEN
            tanh_f := - 2008;
        ELSIF x =- 4720 THEN
            tanh_f := - 2008;
        ELSIF x =- 4719 THEN
            tanh_f := - 2008;
        ELSIF x =- 4718 THEN
            tanh_f := - 2008;
        ELSIF x =- 4717 THEN
            tanh_f := - 2008;
        ELSIF x =- 4716 THEN
            tanh_f := - 2008;
        ELSIF x =- 4715 THEN
            tanh_f := - 2008;
        ELSIF x =- 4714 THEN
            tanh_f := - 2008;
        ELSIF x =- 4713 THEN
            tanh_f := - 2008;
        ELSIF x =- 4712 THEN
            tanh_f := - 2008;
        ELSIF x =- 4711 THEN
            tanh_f := - 2008;
        ELSIF x =- 4710 THEN
            tanh_f := - 2008;
        ELSIF x =- 4709 THEN
            tanh_f := - 2008;
        ELSIF x =- 4708 THEN
            tanh_f := - 2008;
        ELSIF x =- 4707 THEN
            tanh_f := - 2008;
        ELSIF x =- 4706 THEN
            tanh_f := - 2008;
        ELSIF x =- 4705 THEN
            tanh_f := - 2007;
        ELSIF x =- 4704 THEN
            tanh_f := - 2007;
        ELSIF x =- 4703 THEN
            tanh_f := - 2007;
        ELSIF x =- 4702 THEN
            tanh_f := - 2007;
        ELSIF x =- 4701 THEN
            tanh_f := - 2007;
        ELSIF x =- 4700 THEN
            tanh_f := - 2007;
        ELSIF x =- 4699 THEN
            tanh_f := - 2007;
        ELSIF x =- 4698 THEN
            tanh_f := - 2007;
        ELSIF x =- 4697 THEN
            tanh_f := - 2007;
        ELSIF x =- 4696 THEN
            tanh_f := - 2007;
        ELSIF x =- 4695 THEN
            tanh_f := - 2007;
        ELSIF x =- 4694 THEN
            tanh_f := - 2007;
        ELSIF x =- 4693 THEN
            tanh_f := - 2007;
        ELSIF x =- 4692 THEN
            tanh_f := - 2007;
        ELSIF x =- 4691 THEN
            tanh_f := - 2007;
        ELSIF x =- 4690 THEN
            tanh_f := - 2007;
        ELSIF x =- 4689 THEN
            tanh_f := - 2007;
        ELSIF x =- 4688 THEN
            tanh_f := - 2007;
        ELSIF x =- 4687 THEN
            tanh_f := - 2007;
        ELSIF x =- 4686 THEN
            tanh_f := - 2007;
        ELSIF x =- 4685 THEN
            tanh_f := - 2007;
        ELSIF x =- 4684 THEN
            tanh_f := - 2007;
        ELSIF x =- 4683 THEN
            tanh_f := - 2007;
        ELSIF x =- 4682 THEN
            tanh_f := - 2007;
        ELSIF x =- 4681 THEN
            tanh_f := - 2006;
        ELSIF x =- 4680 THEN
            tanh_f := - 2006;
        ELSIF x =- 4679 THEN
            tanh_f := - 2006;
        ELSIF x =- 4678 THEN
            tanh_f := - 2006;
        ELSIF x =- 4677 THEN
            tanh_f := - 2006;
        ELSIF x =- 4676 THEN
            tanh_f := - 2006;
        ELSIF x =- 4675 THEN
            tanh_f := - 2006;
        ELSIF x =- 4674 THEN
            tanh_f := - 2006;
        ELSIF x =- 4673 THEN
            tanh_f := - 2006;
        ELSIF x =- 4672 THEN
            tanh_f := - 2006;
        ELSIF x =- 4671 THEN
            tanh_f := - 2006;
        ELSIF x =- 4670 THEN
            tanh_f := - 2006;
        ELSIF x =- 4669 THEN
            tanh_f := - 2006;
        ELSIF x =- 4668 THEN
            tanh_f := - 2006;
        ELSIF x =- 4667 THEN
            tanh_f := - 2006;
        ELSIF x =- 4666 THEN
            tanh_f := - 2006;
        ELSIF x =- 4665 THEN
            tanh_f := - 2006;
        ELSIF x =- 4664 THEN
            tanh_f := - 2006;
        ELSIF x =- 4663 THEN
            tanh_f := - 2006;
        ELSIF x =- 4662 THEN
            tanh_f := - 2006;
        ELSIF x =- 4661 THEN
            tanh_f := - 2006;
        ELSIF x =- 4660 THEN
            tanh_f := - 2006;
        ELSIF x =- 4659 THEN
            tanh_f := - 2006;
        ELSIF x =- 4658 THEN
            tanh_f := - 2006;
        ELSIF x =- 4657 THEN
            tanh_f := - 2006;
        ELSIF x =- 4656 THEN
            tanh_f := - 2005;
        ELSIF x =- 4655 THEN
            tanh_f := - 2005;
        ELSIF x =- 4654 THEN
            tanh_f := - 2005;
        ELSIF x =- 4653 THEN
            tanh_f := - 2005;
        ELSIF x =- 4652 THEN
            tanh_f := - 2005;
        ELSIF x =- 4651 THEN
            tanh_f := - 2005;
        ELSIF x =- 4650 THEN
            tanh_f := - 2005;
        ELSIF x =- 4649 THEN
            tanh_f := - 2005;
        ELSIF x =- 4648 THEN
            tanh_f := - 2005;
        ELSIF x =- 4647 THEN
            tanh_f := - 2005;
        ELSIF x =- 4646 THEN
            tanh_f := - 2005;
        ELSIF x =- 4645 THEN
            tanh_f := - 2005;
        ELSIF x =- 4644 THEN
            tanh_f := - 2005;
        ELSIF x =- 4643 THEN
            tanh_f := - 2005;
        ELSIF x =- 4642 THEN
            tanh_f := - 2005;
        ELSIF x =- 4641 THEN
            tanh_f := - 2005;
        ELSIF x =- 4640 THEN
            tanh_f := - 2005;
        ELSIF x =- 4639 THEN
            tanh_f := - 2005;
        ELSIF x =- 4638 THEN
            tanh_f := - 2005;
        ELSIF x =- 4637 THEN
            tanh_f := - 2005;
        ELSIF x =- 4636 THEN
            tanh_f := - 2005;
        ELSIF x =- 4635 THEN
            tanh_f := - 2005;
        ELSIF x =- 4634 THEN
            tanh_f := - 2005;
        ELSIF x =- 4633 THEN
            tanh_f := - 2005;
        ELSIF x =- 4632 THEN
            tanh_f := - 2004;
        ELSIF x =- 4631 THEN
            tanh_f := - 2004;
        ELSIF x =- 4630 THEN
            tanh_f := - 2004;
        ELSIF x =- 4629 THEN
            tanh_f := - 2004;
        ELSIF x =- 4628 THEN
            tanh_f := - 2004;
        ELSIF x =- 4627 THEN
            tanh_f := - 2004;
        ELSIF x =- 4626 THEN
            tanh_f := - 2004;
        ELSIF x =- 4625 THEN
            tanh_f := - 2004;
        ELSIF x =- 4624 THEN
            tanh_f := - 2004;
        ELSIF x =- 4623 THEN
            tanh_f := - 2004;
        ELSIF x =- 4622 THEN
            tanh_f := - 2004;
        ELSIF x =- 4621 THEN
            tanh_f := - 2004;
        ELSIF x =- 4620 THEN
            tanh_f := - 2004;
        ELSIF x =- 4619 THEN
            tanh_f := - 2004;
        ELSIF x =- 4618 THEN
            tanh_f := - 2004;
        ELSIF x =- 4617 THEN
            tanh_f := - 2004;
        ELSIF x =- 4616 THEN
            tanh_f := - 2004;
        ELSIF x =- 4615 THEN
            tanh_f := - 2004;
        ELSIF x =- 4614 THEN
            tanh_f := - 2004;
        ELSIF x =- 4613 THEN
            tanh_f := - 2004;
        ELSIF x =- 4612 THEN
            tanh_f := - 2004;
        ELSIF x =- 4611 THEN
            tanh_f := - 2004;
        ELSIF x =- 4610 THEN
            tanh_f := - 2004;
        ELSIF x =- 4609 THEN
            tanh_f := - 2004;
        ELSIF x =- 4608 THEN
            tanh_f := - 2003;
        ELSIF x =- 4607 THEN
            tanh_f := - 2003;
        ELSIF x =- 4606 THEN
            tanh_f := - 2003;
        ELSIF x =- 4605 THEN
            tanh_f := - 2003;
        ELSIF x =- 4604 THEN
            tanh_f := - 2003;
        ELSIF x =- 4603 THEN
            tanh_f := - 2003;
        ELSIF x =- 4602 THEN
            tanh_f := - 2003;
        ELSIF x =- 4601 THEN
            tanh_f := - 2003;
        ELSIF x =- 4600 THEN
            tanh_f := - 2003;
        ELSIF x =- 4599 THEN
            tanh_f := - 2003;
        ELSIF x =- 4598 THEN
            tanh_f := - 2003;
        ELSIF x =- 4597 THEN
            tanh_f := - 2003;
        ELSIF x =- 4596 THEN
            tanh_f := - 2003;
        ELSIF x =- 4595 THEN
            tanh_f := - 2003;
        ELSIF x =- 4594 THEN
            tanh_f := - 2003;
        ELSIF x =- 4593 THEN
            tanh_f := - 2003;
        ELSIF x =- 4592 THEN
            tanh_f := - 2003;
        ELSIF x =- 4591 THEN
            tanh_f := - 2003;
        ELSIF x =- 4590 THEN
            tanh_f := - 2003;
        ELSIF x =- 4589 THEN
            tanh_f := - 2003;
        ELSIF x =- 4588 THEN
            tanh_f := - 2003;
        ELSIF x =- 4587 THEN
            tanh_f := - 2002;
        ELSIF x =- 4586 THEN
            tanh_f := - 2002;
        ELSIF x =- 4585 THEN
            tanh_f := - 2002;
        ELSIF x =- 4584 THEN
            tanh_f := - 2002;
        ELSIF x =- 4583 THEN
            tanh_f := - 2002;
        ELSIF x =- 4582 THEN
            tanh_f := - 2002;
        ELSIF x =- 4581 THEN
            tanh_f := - 2002;
        ELSIF x =- 4580 THEN
            tanh_f := - 2002;
        ELSIF x =- 4579 THEN
            tanh_f := - 2002;
        ELSIF x =- 4578 THEN
            tanh_f := - 2002;
        ELSIF x =- 4577 THEN
            tanh_f := - 2002;
        ELSIF x =- 4576 THEN
            tanh_f := - 2002;
        ELSIF x =- 4575 THEN
            tanh_f := - 2002;
        ELSIF x =- 4574 THEN
            tanh_f := - 2002;
        ELSIF x =- 4573 THEN
            tanh_f := - 2002;
        ELSIF x =- 4572 THEN
            tanh_f := - 2002;
        ELSIF x =- 4571 THEN
            tanh_f := - 2002;
        ELSIF x =- 4570 THEN
            tanh_f := - 2002;
        ELSIF x =- 4569 THEN
            tanh_f := - 2002;
        ELSIF x =- 4568 THEN
            tanh_f := - 2002;
        ELSIF x =- 4567 THEN
            tanh_f := - 2001;
        ELSIF x =- 4566 THEN
            tanh_f := - 2001;
        ELSIF x =- 4565 THEN
            tanh_f := - 2001;
        ELSIF x =- 4564 THEN
            tanh_f := - 2001;
        ELSIF x =- 4563 THEN
            tanh_f := - 2001;
        ELSIF x =- 4562 THEN
            tanh_f := - 2001;
        ELSIF x =- 4561 THEN
            tanh_f := - 2001;
        ELSIF x =- 4560 THEN
            tanh_f := - 2001;
        ELSIF x =- 4559 THEN
            tanh_f := - 2001;
        ELSIF x =- 4558 THEN
            tanh_f := - 2001;
        ELSIF x =- 4557 THEN
            tanh_f := - 2001;
        ELSIF x =- 4556 THEN
            tanh_f := - 2001;
        ELSIF x =- 4555 THEN
            tanh_f := - 2001;
        ELSIF x =- 4554 THEN
            tanh_f := - 2001;
        ELSIF x =- 4553 THEN
            tanh_f := - 2001;
        ELSIF x =- 4552 THEN
            tanh_f := - 2001;
        ELSIF x =- 4551 THEN
            tanh_f := - 2001;
        ELSIF x =- 4550 THEN
            tanh_f := - 2001;
        ELSIF x =- 4549 THEN
            tanh_f := - 2001;
        ELSIF x =- 4548 THEN
            tanh_f := - 2001;
        ELSIF x =- 4547 THEN
            tanh_f := - 2001;
        ELSIF x =- 4546 THEN
            tanh_f := - 2000;
        ELSIF x =- 4545 THEN
            tanh_f := - 2000;
        ELSIF x =- 4544 THEN
            tanh_f := - 2000;
        ELSIF x =- 4543 THEN
            tanh_f := - 2000;
        ELSIF x =- 4542 THEN
            tanh_f := - 2000;
        ELSIF x =- 4541 THEN
            tanh_f := - 2000;
        ELSIF x =- 4540 THEN
            tanh_f := - 2000;
        ELSIF x =- 4539 THEN
            tanh_f := - 2000;
        ELSIF x =- 4538 THEN
            tanh_f := - 2000;
        ELSIF x =- 4537 THEN
            tanh_f := - 2000;
        ELSIF x =- 4536 THEN
            tanh_f := - 2000;
        ELSIF x =- 4535 THEN
            tanh_f := - 2000;
        ELSIF x =- 4534 THEN
            tanh_f := - 2000;
        ELSIF x =- 4533 THEN
            tanh_f := - 2000;
        ELSIF x =- 4532 THEN
            tanh_f := - 2000;
        ELSIF x =- 4531 THEN
            tanh_f := - 2000;
        ELSIF x =- 4530 THEN
            tanh_f := - 2000;
        ELSIF x =- 4529 THEN
            tanh_f := - 2000;
        ELSIF x =- 4528 THEN
            tanh_f := - 2000;
        ELSIF x =- 4527 THEN
            tanh_f := - 2000;
        ELSIF x =- 4526 THEN
            tanh_f := - 1999;
        ELSIF x =- 4525 THEN
            tanh_f := - 1999;
        ELSIF x =- 4524 THEN
            tanh_f := - 1999;
        ELSIF x =- 4523 THEN
            tanh_f := - 1999;
        ELSIF x =- 4522 THEN
            tanh_f := - 1999;
        ELSIF x =- 4521 THEN
            tanh_f := - 1999;
        ELSIF x =- 4520 THEN
            tanh_f := - 1999;
        ELSIF x =- 4519 THEN
            tanh_f := - 1999;
        ELSIF x =- 4518 THEN
            tanh_f := - 1999;
        ELSIF x =- 4517 THEN
            tanh_f := - 1999;
        ELSIF x =- 4516 THEN
            tanh_f := - 1999;
        ELSIF x =- 4515 THEN
            tanh_f := - 1999;
        ELSIF x =- 4514 THEN
            tanh_f := - 1999;
        ELSIF x =- 4513 THEN
            tanh_f := - 1999;
        ELSIF x =- 4512 THEN
            tanh_f := - 1999;
        ELSIF x =- 4511 THEN
            tanh_f := - 1999;
        ELSIF x =- 4510 THEN
            tanh_f := - 1999;
        ELSIF x =- 4509 THEN
            tanh_f := - 1999;
        ELSIF x =- 4508 THEN
            tanh_f := - 1999;
        ELSIF x =- 4507 THEN
            tanh_f := - 1999;
        ELSIF x =- 4506 THEN
            tanh_f := - 1999;
        ELSIF x =- 4505 THEN
            tanh_f := - 1998;
        ELSIF x =- 4504 THEN
            tanh_f := - 1998;
        ELSIF x =- 4503 THEN
            tanh_f := - 1998;
        ELSIF x =- 4502 THEN
            tanh_f := - 1998;
        ELSIF x =- 4501 THEN
            tanh_f := - 1998;
        ELSIF x =- 4500 THEN
            tanh_f := - 1998;
        ELSIF x =- 4499 THEN
            tanh_f := - 1998;
        ELSIF x =- 4498 THEN
            tanh_f := - 1998;
        ELSIF x =- 4497 THEN
            tanh_f := - 1998;
        ELSIF x =- 4496 THEN
            tanh_f := - 1998;
        ELSIF x =- 4495 THEN
            tanh_f := - 1998;
        ELSIF x =- 4494 THEN
            tanh_f := - 1998;
        ELSIF x =- 4493 THEN
            tanh_f := - 1998;
        ELSIF x =- 4492 THEN
            tanh_f := - 1998;
        ELSIF x =- 4491 THEN
            tanh_f := - 1998;
        ELSIF x =- 4490 THEN
            tanh_f := - 1998;
        ELSIF x =- 4489 THEN
            tanh_f := - 1998;
        ELSIF x =- 4488 THEN
            tanh_f := - 1998;
        ELSIF x =- 4487 THEN
            tanh_f := - 1998;
        ELSIF x =- 4486 THEN
            tanh_f := - 1998;
        ELSIF x =- 4485 THEN
            tanh_f := - 1997;
        ELSIF x =- 4484 THEN
            tanh_f := - 1997;
        ELSIF x =- 4483 THEN
            tanh_f := - 1997;
        ELSIF x =- 4482 THEN
            tanh_f := - 1997;
        ELSIF x =- 4481 THEN
            tanh_f := - 1997;
        ELSIF x =- 4480 THEN
            tanh_f := - 1997;
        ELSIF x =- 4479 THEN
            tanh_f := - 1997;
        ELSIF x =- 4478 THEN
            tanh_f := - 1997;
        ELSIF x =- 4477 THEN
            tanh_f := - 1997;
        ELSIF x =- 4476 THEN
            tanh_f := - 1997;
        ELSIF x =- 4475 THEN
            tanh_f := - 1997;
        ELSIF x =- 4474 THEN
            tanh_f := - 1997;
        ELSIF x =- 4473 THEN
            tanh_f := - 1997;
        ELSIF x =- 4472 THEN
            tanh_f := - 1997;
        ELSIF x =- 4471 THEN
            tanh_f := - 1997;
        ELSIF x =- 4470 THEN
            tanh_f := - 1997;
        ELSIF x =- 4469 THEN
            tanh_f := - 1997;
        ELSIF x =- 4468 THEN
            tanh_f := - 1997;
        ELSIF x =- 4467 THEN
            tanh_f := - 1997;
        ELSIF x =- 4466 THEN
            tanh_f := - 1997;
        ELSIF x =- 4465 THEN
            tanh_f := - 1997;
        ELSIF x =- 4464 THEN
            tanh_f := - 1996;
        ELSIF x =- 4463 THEN
            tanh_f := - 1996;
        ELSIF x =- 4462 THEN
            tanh_f := - 1996;
        ELSIF x =- 4461 THEN
            tanh_f := - 1996;
        ELSIF x =- 4460 THEN
            tanh_f := - 1996;
        ELSIF x =- 4459 THEN
            tanh_f := - 1996;
        ELSIF x =- 4458 THEN
            tanh_f := - 1996;
        ELSIF x =- 4457 THEN
            tanh_f := - 1996;
        ELSIF x =- 4456 THEN
            tanh_f := - 1996;
        ELSIF x =- 4455 THEN
            tanh_f := - 1996;
        ELSIF x =- 4454 THEN
            tanh_f := - 1996;
        ELSIF x =- 4453 THEN
            tanh_f := - 1996;
        ELSIF x =- 4452 THEN
            tanh_f := - 1996;
        ELSIF x =- 4451 THEN
            tanh_f := - 1996;
        ELSIF x =- 4450 THEN
            tanh_f := - 1996;
        ELSIF x =- 4449 THEN
            tanh_f := - 1996;
        ELSIF x =- 4448 THEN
            tanh_f := - 1996;
        ELSIF x =- 4447 THEN
            tanh_f := - 1996;
        ELSIF x =- 4446 THEN
            tanh_f := - 1996;
        ELSIF x =- 4445 THEN
            tanh_f := - 1996;
        ELSIF x =- 4444 THEN
            tanh_f := - 1995;
        ELSIF x =- 4443 THEN
            tanh_f := - 1995;
        ELSIF x =- 4442 THEN
            tanh_f := - 1995;
        ELSIF x =- 4441 THEN
            tanh_f := - 1995;
        ELSIF x =- 4440 THEN
            tanh_f := - 1995;
        ELSIF x =- 4439 THEN
            tanh_f := - 1995;
        ELSIF x =- 4438 THEN
            tanh_f := - 1995;
        ELSIF x =- 4437 THEN
            tanh_f := - 1995;
        ELSIF x =- 4436 THEN
            tanh_f := - 1995;
        ELSIF x =- 4435 THEN
            tanh_f := - 1995;
        ELSIF x =- 4434 THEN
            tanh_f := - 1995;
        ELSIF x =- 4433 THEN
            tanh_f := - 1995;
        ELSIF x =- 4432 THEN
            tanh_f := - 1995;
        ELSIF x =- 4431 THEN
            tanh_f := - 1995;
        ELSIF x =- 4430 THEN
            tanh_f := - 1995;
        ELSIF x =- 4429 THEN
            tanh_f := - 1995;
        ELSIF x =- 4428 THEN
            tanh_f := - 1995;
        ELSIF x =- 4427 THEN
            tanh_f := - 1995;
        ELSIF x =- 4426 THEN
            tanh_f := - 1995;
        ELSIF x =- 4425 THEN
            tanh_f := - 1995;
        ELSIF x =- 4424 THEN
            tanh_f := - 1995;
        ELSIF x =- 4423 THEN
            tanh_f := - 1994;
        ELSIF x =- 4422 THEN
            tanh_f := - 1994;
        ELSIF x =- 4421 THEN
            tanh_f := - 1994;
        ELSIF x =- 4420 THEN
            tanh_f := - 1994;
        ELSIF x =- 4419 THEN
            tanh_f := - 1994;
        ELSIF x =- 4418 THEN
            tanh_f := - 1994;
        ELSIF x =- 4417 THEN
            tanh_f := - 1994;
        ELSIF x =- 4416 THEN
            tanh_f := - 1994;
        ELSIF x =- 4415 THEN
            tanh_f := - 1994;
        ELSIF x =- 4414 THEN
            tanh_f := - 1994;
        ELSIF x =- 4413 THEN
            tanh_f := - 1994;
        ELSIF x =- 4412 THEN
            tanh_f := - 1994;
        ELSIF x =- 4411 THEN
            tanh_f := - 1994;
        ELSIF x =- 4410 THEN
            tanh_f := - 1994;
        ELSIF x =- 4409 THEN
            tanh_f := - 1994;
        ELSIF x =- 4408 THEN
            tanh_f := - 1994;
        ELSIF x =- 4407 THEN
            tanh_f := - 1994;
        ELSIF x =- 4406 THEN
            tanh_f := - 1994;
        ELSIF x =- 4405 THEN
            tanh_f := - 1994;
        ELSIF x =- 4404 THEN
            tanh_f := - 1994;
        ELSIF x =- 4403 THEN
            tanh_f := - 1993;
        ELSIF x =- 4402 THEN
            tanh_f := - 1993;
        ELSIF x =- 4401 THEN
            tanh_f := - 1993;
        ELSIF x =- 4400 THEN
            tanh_f := - 1993;
        ELSIF x =- 4399 THEN
            tanh_f := - 1993;
        ELSIF x =- 4398 THEN
            tanh_f := - 1993;
        ELSIF x =- 4397 THEN
            tanh_f := - 1993;
        ELSIF x =- 4396 THEN
            tanh_f := - 1993;
        ELSIF x =- 4395 THEN
            tanh_f := - 1993;
        ELSIF x =- 4394 THEN
            tanh_f := - 1993;
        ELSIF x =- 4393 THEN
            tanh_f := - 1993;
        ELSIF x =- 4392 THEN
            tanh_f := - 1993;
        ELSIF x =- 4391 THEN
            tanh_f := - 1993;
        ELSIF x =- 4390 THEN
            tanh_f := - 1993;
        ELSIF x =- 4389 THEN
            tanh_f := - 1993;
        ELSIF x =- 4388 THEN
            tanh_f := - 1993;
        ELSIF x =- 4387 THEN
            tanh_f := - 1993;
        ELSIF x =- 4386 THEN
            tanh_f := - 1993;
        ELSIF x =- 4385 THEN
            tanh_f := - 1993;
        ELSIF x =- 4384 THEN
            tanh_f := - 1993;
        ELSIF x =- 4383 THEN
            tanh_f := - 1993;
        ELSIF x =- 4382 THEN
            tanh_f := - 1992;
        ELSIF x =- 4381 THEN
            tanh_f := - 1992;
        ELSIF x =- 4380 THEN
            tanh_f := - 1992;
        ELSIF x =- 4379 THEN
            tanh_f := - 1992;
        ELSIF x =- 4378 THEN
            tanh_f := - 1992;
        ELSIF x =- 4377 THEN
            tanh_f := - 1992;
        ELSIF x =- 4376 THEN
            tanh_f := - 1992;
        ELSIF x =- 4375 THEN
            tanh_f := - 1992;
        ELSIF x =- 4374 THEN
            tanh_f := - 1992;
        ELSIF x =- 4373 THEN
            tanh_f := - 1992;
        ELSIF x =- 4372 THEN
            tanh_f := - 1992;
        ELSIF x =- 4371 THEN
            tanh_f := - 1992;
        ELSIF x =- 4370 THEN
            tanh_f := - 1992;
        ELSIF x =- 4369 THEN
            tanh_f := - 1992;
        ELSIF x =- 4368 THEN
            tanh_f := - 1992;
        ELSIF x =- 4367 THEN
            tanh_f := - 1992;
        ELSIF x =- 4366 THEN
            tanh_f := - 1992;
        ELSIF x =- 4365 THEN
            tanh_f := - 1992;
        ELSIF x =- 4364 THEN
            tanh_f := - 1992;
        ELSIF x =- 4363 THEN
            tanh_f := - 1992;
        ELSIF x =- 4362 THEN
            tanh_f := - 1991;
        ELSIF x =- 4361 THEN
            tanh_f := - 1991;
        ELSIF x =- 4360 THEN
            tanh_f := - 1991;
        ELSIF x =- 4359 THEN
            tanh_f := - 1991;
        ELSIF x =- 4358 THEN
            tanh_f := - 1991;
        ELSIF x =- 4357 THEN
            tanh_f := - 1991;
        ELSIF x =- 4356 THEN
            tanh_f := - 1991;
        ELSIF x =- 4355 THEN
            tanh_f := - 1991;
        ELSIF x =- 4354 THEN
            tanh_f := - 1991;
        ELSIF x =- 4353 THEN
            tanh_f := - 1991;
        ELSIF x =- 4352 THEN
            tanh_f := - 1991;
        ELSIF x =- 4351 THEN
            tanh_f := - 1991;
        ELSIF x =- 4350 THEN
            tanh_f := - 1991;
        ELSIF x =- 4349 THEN
            tanh_f := - 1991;
        ELSIF x =- 4348 THEN
            tanh_f := - 1991;
        ELSIF x =- 4347 THEN
            tanh_f := - 1991;
        ELSIF x =- 4346 THEN
            tanh_f := - 1991;
        ELSIF x =- 4345 THEN
            tanh_f := - 1991;
        ELSIF x =- 4344 THEN
            tanh_f := - 1991;
        ELSIF x =- 4343 THEN
            tanh_f := - 1991;
        ELSIF x =- 4342 THEN
            tanh_f := - 1991;
        ELSIF x =- 4341 THEN
            tanh_f := - 1991;
        ELSIF x =- 4340 THEN
            tanh_f := - 1991;
        ELSIF x =- 4339 THEN
            tanh_f := - 1991;
        ELSIF x =- 4338 THEN
            tanh_f := - 1991;
        ELSIF x =- 4337 THEN
            tanh_f := - 1991;
        ELSIF x =- 4336 THEN
            tanh_f := - 1990;
        ELSIF x =- 4335 THEN
            tanh_f := - 1990;
        ELSIF x =- 4334 THEN
            tanh_f := - 1990;
        ELSIF x =- 4333 THEN
            tanh_f := - 1990;
        ELSIF x =- 4332 THEN
            tanh_f := - 1990;
        ELSIF x =- 4331 THEN
            tanh_f := - 1990;
        ELSIF x =- 4330 THEN
            tanh_f := - 1990;
        ELSIF x =- 4329 THEN
            tanh_f := - 1990;
        ELSIF x =- 4328 THEN
            tanh_f := - 1990;
        ELSIF x =- 4327 THEN
            tanh_f := - 1990;
        ELSIF x =- 4326 THEN
            tanh_f := - 1990;
        ELSIF x =- 4325 THEN
            tanh_f := - 1990;
        ELSIF x =- 4324 THEN
            tanh_f := - 1990;
        ELSIF x =- 4323 THEN
            tanh_f := - 1990;
        ELSIF x =- 4322 THEN
            tanh_f := - 1990;
        ELSIF x =- 4321 THEN
            tanh_f := - 1989;
        ELSIF x =- 4320 THEN
            tanh_f := - 1989;
        ELSIF x =- 4319 THEN
            tanh_f := - 1989;
        ELSIF x =- 4318 THEN
            tanh_f := - 1989;
        ELSIF x =- 4317 THEN
            tanh_f := - 1989;
        ELSIF x =- 4316 THEN
            tanh_f := - 1989;
        ELSIF x =- 4315 THEN
            tanh_f := - 1989;
        ELSIF x =- 4314 THEN
            tanh_f := - 1989;
        ELSIF x =- 4313 THEN
            tanh_f := - 1989;
        ELSIF x =- 4312 THEN
            tanh_f := - 1989;
        ELSIF x =- 4311 THEN
            tanh_f := - 1989;
        ELSIF x =- 4310 THEN
            tanh_f := - 1989;
        ELSIF x =- 4309 THEN
            tanh_f := - 1989;
        ELSIF x =- 4308 THEN
            tanh_f := - 1989;
        ELSIF x =- 4307 THEN
            tanh_f := - 1989;
        ELSIF x =- 4306 THEN
            tanh_f := - 1988;
        ELSIF x =- 4305 THEN
            tanh_f := - 1988;
        ELSIF x =- 4304 THEN
            tanh_f := - 1988;
        ELSIF x =- 4303 THEN
            tanh_f := - 1988;
        ELSIF x =- 4302 THEN
            tanh_f := - 1988;
        ELSIF x =- 4301 THEN
            tanh_f := - 1988;
        ELSIF x =- 4300 THEN
            tanh_f := - 1988;
        ELSIF x =- 4299 THEN
            tanh_f := - 1988;
        ELSIF x =- 4298 THEN
            tanh_f := - 1988;
        ELSIF x =- 4297 THEN
            tanh_f := - 1988;
        ELSIF x =- 4296 THEN
            tanh_f := - 1988;
        ELSIF x =- 4295 THEN
            tanh_f := - 1988;
        ELSIF x =- 4294 THEN
            tanh_f := - 1988;
        ELSIF x =- 4293 THEN
            tanh_f := - 1988;
        ELSIF x =- 4292 THEN
            tanh_f := - 1988;
        ELSIF x =- 4291 THEN
            tanh_f := - 1987;
        ELSIF x =- 4290 THEN
            tanh_f := - 1987;
        ELSIF x =- 4289 THEN
            tanh_f := - 1987;
        ELSIF x =- 4288 THEN
            tanh_f := - 1987;
        ELSIF x =- 4287 THEN
            tanh_f := - 1987;
        ELSIF x =- 4286 THEN
            tanh_f := - 1987;
        ELSIF x =- 4285 THEN
            tanh_f := - 1987;
        ELSIF x =- 4284 THEN
            tanh_f := - 1987;
        ELSIF x =- 4283 THEN
            tanh_f := - 1987;
        ELSIF x =- 4282 THEN
            tanh_f := - 1987;
        ELSIF x =- 4281 THEN
            tanh_f := - 1987;
        ELSIF x =- 4280 THEN
            tanh_f := - 1987;
        ELSIF x =- 4279 THEN
            tanh_f := - 1987;
        ELSIF x =- 4278 THEN
            tanh_f := - 1987;
        ELSIF x =- 4277 THEN
            tanh_f := - 1987;
        ELSIF x =- 4276 THEN
            tanh_f := - 1986;
        ELSIF x =- 4275 THEN
            tanh_f := - 1986;
        ELSIF x =- 4274 THEN
            tanh_f := - 1986;
        ELSIF x =- 4273 THEN
            tanh_f := - 1986;
        ELSIF x =- 4272 THEN
            tanh_f := - 1986;
        ELSIF x =- 4271 THEN
            tanh_f := - 1986;
        ELSIF x =- 4270 THEN
            tanh_f := - 1986;
        ELSIF x =- 4269 THEN
            tanh_f := - 1986;
        ELSIF x =- 4268 THEN
            tanh_f := - 1986;
        ELSIF x =- 4267 THEN
            tanh_f := - 1986;
        ELSIF x =- 4266 THEN
            tanh_f := - 1986;
        ELSIF x =- 4265 THEN
            tanh_f := - 1986;
        ELSIF x =- 4264 THEN
            tanh_f := - 1986;
        ELSIF x =- 4263 THEN
            tanh_f := - 1986;
        ELSIF x =- 4262 THEN
            tanh_f := - 1986;
        ELSIF x =- 4261 THEN
            tanh_f := - 1985;
        ELSIF x =- 4260 THEN
            tanh_f := - 1985;
        ELSIF x =- 4259 THEN
            tanh_f := - 1985;
        ELSIF x =- 4258 THEN
            tanh_f := - 1985;
        ELSIF x =- 4257 THEN
            tanh_f := - 1985;
        ELSIF x =- 4256 THEN
            tanh_f := - 1985;
        ELSIF x =- 4255 THEN
            tanh_f := - 1985;
        ELSIF x =- 4254 THEN
            tanh_f := - 1985;
        ELSIF x =- 4253 THEN
            tanh_f := - 1985;
        ELSIF x =- 4252 THEN
            tanh_f := - 1985;
        ELSIF x =- 4251 THEN
            tanh_f := - 1985;
        ELSIF x =- 4250 THEN
            tanh_f := - 1985;
        ELSIF x =- 4249 THEN
            tanh_f := - 1985;
        ELSIF x =- 4248 THEN
            tanh_f := - 1985;
        ELSIF x =- 4247 THEN
            tanh_f := - 1985;
        ELSIF x =- 4246 THEN
            tanh_f := - 1984;
        ELSIF x =- 4245 THEN
            tanh_f := - 1984;
        ELSIF x =- 4244 THEN
            tanh_f := - 1984;
        ELSIF x =- 4243 THEN
            tanh_f := - 1984;
        ELSIF x =- 4242 THEN
            tanh_f := - 1984;
        ELSIF x =- 4241 THEN
            tanh_f := - 1984;
        ELSIF x =- 4240 THEN
            tanh_f := - 1984;
        ELSIF x =- 4239 THEN
            tanh_f := - 1984;
        ELSIF x =- 4238 THEN
            tanh_f := - 1984;
        ELSIF x =- 4237 THEN
            tanh_f := - 1984;
        ELSIF x =- 4236 THEN
            tanh_f := - 1984;
        ELSIF x =- 4235 THEN
            tanh_f := - 1984;
        ELSIF x =- 4234 THEN
            tanh_f := - 1984;
        ELSIF x =- 4233 THEN
            tanh_f := - 1984;
        ELSIF x =- 4232 THEN
            tanh_f := - 1984;
        ELSIF x =- 4231 THEN
            tanh_f := - 1983;
        ELSIF x =- 4230 THEN
            tanh_f := - 1983;
        ELSIF x =- 4229 THEN
            tanh_f := - 1983;
        ELSIF x =- 4228 THEN
            tanh_f := - 1983;
        ELSIF x =- 4227 THEN
            tanh_f := - 1983;
        ELSIF x =- 4226 THEN
            tanh_f := - 1983;
        ELSIF x =- 4225 THEN
            tanh_f := - 1983;
        ELSIF x =- 4224 THEN
            tanh_f := - 1983;
        ELSIF x =- 4223 THEN
            tanh_f := - 1983;
        ELSIF x =- 4222 THEN
            tanh_f := - 1983;
        ELSIF x =- 4221 THEN
            tanh_f := - 1983;
        ELSIF x =- 4220 THEN
            tanh_f := - 1983;
        ELSIF x =- 4219 THEN
            tanh_f := - 1983;
        ELSIF x =- 4218 THEN
            tanh_f := - 1983;
        ELSIF x =- 4217 THEN
            tanh_f := - 1983;
        ELSIF x =- 4216 THEN
            tanh_f := - 1982;
        ELSIF x =- 4215 THEN
            tanh_f := - 1982;
        ELSIF x =- 4214 THEN
            tanh_f := - 1982;
        ELSIF x =- 4213 THEN
            tanh_f := - 1982;
        ELSIF x =- 4212 THEN
            tanh_f := - 1982;
        ELSIF x =- 4211 THEN
            tanh_f := - 1982;
        ELSIF x =- 4210 THEN
            tanh_f := - 1982;
        ELSIF x =- 4209 THEN
            tanh_f := - 1982;
        ELSIF x =- 4208 THEN
            tanh_f := - 1982;
        ELSIF x =- 4207 THEN
            tanh_f := - 1982;
        ELSIF x =- 4206 THEN
            tanh_f := - 1982;
        ELSIF x =- 4205 THEN
            tanh_f := - 1982;
        ELSIF x =- 4204 THEN
            tanh_f := - 1982;
        ELSIF x =- 4203 THEN
            tanh_f := - 1982;
        ELSIF x =- 4202 THEN
            tanh_f := - 1982;
        ELSIF x =- 4201 THEN
            tanh_f := - 1981;
        ELSIF x =- 4200 THEN
            tanh_f := - 1981;
        ELSIF x =- 4199 THEN
            tanh_f := - 1981;
        ELSIF x =- 4198 THEN
            tanh_f := - 1981;
        ELSIF x =- 4197 THEN
            tanh_f := - 1981;
        ELSIF x =- 4196 THEN
            tanh_f := - 1981;
        ELSIF x =- 4195 THEN
            tanh_f := - 1981;
        ELSIF x =- 4194 THEN
            tanh_f := - 1981;
        ELSIF x =- 4193 THEN
            tanh_f := - 1981;
        ELSIF x =- 4192 THEN
            tanh_f := - 1981;
        ELSIF x =- 4191 THEN
            tanh_f := - 1981;
        ELSIF x =- 4190 THEN
            tanh_f := - 1981;
        ELSIF x =- 4189 THEN
            tanh_f := - 1981;
        ELSIF x =- 4188 THEN
            tanh_f := - 1981;
        ELSIF x =- 4187 THEN
            tanh_f := - 1981;
        ELSIF x =- 4186 THEN
            tanh_f := - 1980;
        ELSIF x =- 4185 THEN
            tanh_f := - 1980;
        ELSIF x =- 4184 THEN
            tanh_f := - 1980;
        ELSIF x =- 4183 THEN
            tanh_f := - 1980;
        ELSIF x =- 4182 THEN
            tanh_f := - 1980;
        ELSIF x =- 4181 THEN
            tanh_f := - 1980;
        ELSIF x =- 4180 THEN
            tanh_f := - 1980;
        ELSIF x =- 4179 THEN
            tanh_f := - 1980;
        ELSIF x =- 4178 THEN
            tanh_f := - 1980;
        ELSIF x =- 4177 THEN
            tanh_f := - 1980;
        ELSIF x =- 4176 THEN
            tanh_f := - 1980;
        ELSIF x =- 4175 THEN
            tanh_f := - 1980;
        ELSIF x =- 4174 THEN
            tanh_f := - 1980;
        ELSIF x =- 4173 THEN
            tanh_f := - 1980;
        ELSIF x =- 4172 THEN
            tanh_f := - 1980;
        ELSIF x =- 4171 THEN
            tanh_f := - 1979;
        ELSIF x =- 4170 THEN
            tanh_f := - 1979;
        ELSIF x =- 4169 THEN
            tanh_f := - 1979;
        ELSIF x =- 4168 THEN
            tanh_f := - 1979;
        ELSIF x =- 4167 THEN
            tanh_f := - 1979;
        ELSIF x =- 4166 THEN
            tanh_f := - 1979;
        ELSIF x =- 4165 THEN
            tanh_f := - 1979;
        ELSIF x =- 4164 THEN
            tanh_f := - 1979;
        ELSIF x =- 4163 THEN
            tanh_f := - 1979;
        ELSIF x =- 4162 THEN
            tanh_f := - 1979;
        ELSIF x =- 4161 THEN
            tanh_f := - 1979;
        ELSIF x =- 4160 THEN
            tanh_f := - 1979;
        ELSIF x =- 4159 THEN
            tanh_f := - 1979;
        ELSIF x =- 4158 THEN
            tanh_f := - 1979;
        ELSIF x =- 4157 THEN
            tanh_f := - 1979;
        ELSIF x =- 4156 THEN
            tanh_f := - 1978;
        ELSIF x =- 4155 THEN
            tanh_f := - 1978;
        ELSIF x =- 4154 THEN
            tanh_f := - 1978;
        ELSIF x =- 4153 THEN
            tanh_f := - 1978;
        ELSIF x =- 4152 THEN
            tanh_f := - 1978;
        ELSIF x =- 4151 THEN
            tanh_f := - 1978;
        ELSIF x =- 4150 THEN
            tanh_f := - 1978;
        ELSIF x =- 4149 THEN
            tanh_f := - 1978;
        ELSIF x =- 4148 THEN
            tanh_f := - 1978;
        ELSIF x =- 4147 THEN
            tanh_f := - 1978;
        ELSIF x =- 4146 THEN
            tanh_f := - 1978;
        ELSIF x =- 4145 THEN
            tanh_f := - 1978;
        ELSIF x =- 4144 THEN
            tanh_f := - 1978;
        ELSIF x =- 4143 THEN
            tanh_f := - 1978;
        ELSIF x =- 4142 THEN
            tanh_f := - 1978;
        ELSIF x =- 4141 THEN
            tanh_f := - 1977;
        ELSIF x =- 4140 THEN
            tanh_f := - 1977;
        ELSIF x =- 4139 THEN
            tanh_f := - 1977;
        ELSIF x =- 4138 THEN
            tanh_f := - 1977;
        ELSIF x =- 4137 THEN
            tanh_f := - 1977;
        ELSIF x =- 4136 THEN
            tanh_f := - 1977;
        ELSIF x =- 4135 THEN
            tanh_f := - 1977;
        ELSIF x =- 4134 THEN
            tanh_f := - 1977;
        ELSIF x =- 4133 THEN
            tanh_f := - 1977;
        ELSIF x =- 4132 THEN
            tanh_f := - 1977;
        ELSIF x =- 4131 THEN
            tanh_f := - 1977;
        ELSIF x =- 4130 THEN
            tanh_f := - 1977;
        ELSIF x =- 4129 THEN
            tanh_f := - 1977;
        ELSIF x =- 4128 THEN
            tanh_f := - 1977;
        ELSIF x =- 4127 THEN
            tanh_f := - 1977;
        ELSIF x =- 4126 THEN
            tanh_f := - 1976;
        ELSIF x =- 4125 THEN
            tanh_f := - 1976;
        ELSIF x =- 4124 THEN
            tanh_f := - 1976;
        ELSIF x =- 4123 THEN
            tanh_f := - 1976;
        ELSIF x =- 4122 THEN
            tanh_f := - 1976;
        ELSIF x =- 4121 THEN
            tanh_f := - 1976;
        ELSIF x =- 4120 THEN
            tanh_f := - 1976;
        ELSIF x =- 4119 THEN
            tanh_f := - 1976;
        ELSIF x =- 4118 THEN
            tanh_f := - 1976;
        ELSIF x =- 4117 THEN
            tanh_f := - 1976;
        ELSIF x =- 4116 THEN
            tanh_f := - 1976;
        ELSIF x =- 4115 THEN
            tanh_f := - 1976;
        ELSIF x =- 4114 THEN
            tanh_f := - 1976;
        ELSIF x =- 4113 THEN
            tanh_f := - 1976;
        ELSIF x =- 4112 THEN
            tanh_f := - 1976;
        ELSIF x =- 4111 THEN
            tanh_f := - 1975;
        ELSIF x =- 4110 THEN
            tanh_f := - 1975;
        ELSIF x =- 4109 THEN
            tanh_f := - 1975;
        ELSIF x =- 4108 THEN
            tanh_f := - 1975;
        ELSIF x =- 4107 THEN
            tanh_f := - 1975;
        ELSIF x =- 4106 THEN
            tanh_f := - 1975;
        ELSIF x =- 4105 THEN
            tanh_f := - 1975;
        ELSIF x =- 4104 THEN
            tanh_f := - 1975;
        ELSIF x =- 4103 THEN
            tanh_f := - 1975;
        ELSIF x =- 4102 THEN
            tanh_f := - 1975;
        ELSIF x =- 4101 THEN
            tanh_f := - 1975;
        ELSIF x =- 4100 THEN
            tanh_f := - 1975;
        ELSIF x =- 4099 THEN
            tanh_f := - 1975;
        ELSIF x =- 4098 THEN
            tanh_f := - 1975;
        ELSIF x =- 4097 THEN
            tanh_f := - 1975;
        ELSIF x =- 4096 THEN
            tanh_f := - 1974;
        ELSIF x =- 4095 THEN
            tanh_f := - 1974;
        ELSIF x =- 4094 THEN
            tanh_f := - 1974;
        ELSIF x =- 4093 THEN
            tanh_f := - 1974;
        ELSIF x =- 4092 THEN
            tanh_f := - 1974;
        ELSIF x =- 4091 THEN
            tanh_f := - 1974;
        ELSIF x =- 4090 THEN
            tanh_f := - 1974;
        ELSIF x =- 4089 THEN
            tanh_f := - 1974;
        ELSIF x =- 4088 THEN
            tanh_f := - 1974;
        ELSIF x =- 4087 THEN
            tanh_f := - 1974;
        ELSIF x =- 4086 THEN
            tanh_f := - 1974;
        ELSIF x =- 4085 THEN
            tanh_f := - 1974;
        ELSIF x =- 4084 THEN
            tanh_f := - 1974;
        ELSIF x =- 4083 THEN
            tanh_f := - 1974;
        ELSIF x =- 4082 THEN
            tanh_f := - 1973;
        ELSIF x =- 4081 THEN
            tanh_f := - 1973;
        ELSIF x =- 4080 THEN
            tanh_f := - 1973;
        ELSIF x =- 4079 THEN
            tanh_f := - 1973;
        ELSIF x =- 4078 THEN
            tanh_f := - 1973;
        ELSIF x =- 4077 THEN
            tanh_f := - 1973;
        ELSIF x =- 4076 THEN
            tanh_f := - 1973;
        ELSIF x =- 4075 THEN
            tanh_f := - 1973;
        ELSIF x =- 4074 THEN
            tanh_f := - 1973;
        ELSIF x =- 4073 THEN
            tanh_f := - 1973;
        ELSIF x =- 4072 THEN
            tanh_f := - 1973;
        ELSIF x =- 4071 THEN
            tanh_f := - 1973;
        ELSIF x =- 4070 THEN
            tanh_f := - 1973;
        ELSIF x =- 4069 THEN
            tanh_f := - 1972;
        ELSIF x =- 4068 THEN
            tanh_f := - 1972;
        ELSIF x =- 4067 THEN
            tanh_f := - 1972;
        ELSIF x =- 4066 THEN
            tanh_f := - 1972;
        ELSIF x =- 4065 THEN
            tanh_f := - 1972;
        ELSIF x =- 4064 THEN
            tanh_f := - 1972;
        ELSIF x =- 4063 THEN
            tanh_f := - 1972;
        ELSIF x =- 4062 THEN
            tanh_f := - 1972;
        ELSIF x =- 4061 THEN
            tanh_f := - 1972;
        ELSIF x =- 4060 THEN
            tanh_f := - 1972;
        ELSIF x =- 4059 THEN
            tanh_f := - 1972;
        ELSIF x =- 4058 THEN
            tanh_f := - 1972;
        ELSIF x =- 4057 THEN
            tanh_f := - 1972;
        ELSIF x =- 4056 THEN
            tanh_f := - 1971;
        ELSIF x =- 4055 THEN
            tanh_f := - 1971;
        ELSIF x =- 4054 THEN
            tanh_f := - 1971;
        ELSIF x =- 4053 THEN
            tanh_f := - 1971;
        ELSIF x =- 4052 THEN
            tanh_f := - 1971;
        ELSIF x =- 4051 THEN
            tanh_f := - 1971;
        ELSIF x =- 4050 THEN
            tanh_f := - 1971;
        ELSIF x =- 4049 THEN
            tanh_f := - 1971;
        ELSIF x =- 4048 THEN
            tanh_f := - 1971;
        ELSIF x =- 4047 THEN
            tanh_f := - 1971;
        ELSIF x =- 4046 THEN
            tanh_f := - 1971;
        ELSIF x =- 4045 THEN
            tanh_f := - 1971;
        ELSIF x =- 4044 THEN
            tanh_f := - 1971;
        ELSIF x =- 4043 THEN
            tanh_f := - 1970;
        ELSIF x =- 4042 THEN
            tanh_f := - 1970;
        ELSIF x =- 4041 THEN
            tanh_f := - 1970;
        ELSIF x =- 4040 THEN
            tanh_f := - 1970;
        ELSIF x =- 4039 THEN
            tanh_f := - 1970;
        ELSIF x =- 4038 THEN
            tanh_f := - 1970;
        ELSIF x =- 4037 THEN
            tanh_f := - 1970;
        ELSIF x =- 4036 THEN
            tanh_f := - 1970;
        ELSIF x =- 4035 THEN
            tanh_f := - 1970;
        ELSIF x =- 4034 THEN
            tanh_f := - 1970;
        ELSIF x =- 4033 THEN
            tanh_f := - 1970;
        ELSIF x =- 4032 THEN
            tanh_f := - 1970;
        ELSIF x =- 4031 THEN
            tanh_f := - 1970;
        ELSIF x =- 4030 THEN
            tanh_f := - 1969;
        ELSIF x =- 4029 THEN
            tanh_f := - 1969;
        ELSIF x =- 4028 THEN
            tanh_f := - 1969;
        ELSIF x =- 4027 THEN
            tanh_f := - 1969;
        ELSIF x =- 4026 THEN
            tanh_f := - 1969;
        ELSIF x =- 4025 THEN
            tanh_f := - 1969;
        ELSIF x =- 4024 THEN
            tanh_f := - 1969;
        ELSIF x =- 4023 THEN
            tanh_f := - 1969;
        ELSIF x =- 4022 THEN
            tanh_f := - 1969;
        ELSIF x =- 4021 THEN
            tanh_f := - 1969;
        ELSIF x =- 4020 THEN
            tanh_f := - 1969;
        ELSIF x =- 4019 THEN
            tanh_f := - 1969;
        ELSIF x =- 4018 THEN
            tanh_f := - 1969;
        ELSIF x =- 4017 THEN
            tanh_f := - 1968;
        ELSIF x =- 4016 THEN
            tanh_f := - 1968;
        ELSIF x =- 4015 THEN
            tanh_f := - 1968;
        ELSIF x =- 4014 THEN
            tanh_f := - 1968;
        ELSIF x =- 4013 THEN
            tanh_f := - 1968;
        ELSIF x =- 4012 THEN
            tanh_f := - 1968;
        ELSIF x =- 4011 THEN
            tanh_f := - 1968;
        ELSIF x =- 4010 THEN
            tanh_f := - 1968;
        ELSIF x =- 4009 THEN
            tanh_f := - 1968;
        ELSIF x =- 4008 THEN
            tanh_f := - 1968;
        ELSIF x =- 4007 THEN
            tanh_f := - 1968;
        ELSIF x =- 4006 THEN
            tanh_f := - 1968;
        ELSIF x =- 4005 THEN
            tanh_f := - 1968;
        ELSIF x =- 4004 THEN
            tanh_f := - 1967;
        ELSIF x =- 4003 THEN
            tanh_f := - 1967;
        ELSIF x =- 4002 THEN
            tanh_f := - 1967;
        ELSIF x =- 4001 THEN
            tanh_f := - 1967;
        ELSIF x =- 4000 THEN
            tanh_f := - 1967;
        ELSIF x =- 3999 THEN
            tanh_f := - 1967;
        ELSIF x =- 3998 THEN
            tanh_f := - 1967;
        ELSIF x =- 3997 THEN
            tanh_f := - 1967;
        ELSIF x =- 3996 THEN
            tanh_f := - 1967;
        ELSIF x =- 3995 THEN
            tanh_f := - 1967;
        ELSIF x =- 3994 THEN
            tanh_f := - 1967;
        ELSIF x =- 3993 THEN
            tanh_f := - 1967;
        ELSIF x =- 3992 THEN
            tanh_f := - 1967;
        ELSIF x =- 3991 THEN
            tanh_f := - 1967;
        ELSIF x =- 3990 THEN
            tanh_f := - 1966;
        ELSIF x =- 3989 THEN
            tanh_f := - 1966;
        ELSIF x =- 3988 THEN
            tanh_f := - 1966;
        ELSIF x =- 3987 THEN
            tanh_f := - 1966;
        ELSIF x =- 3986 THEN
            tanh_f := - 1966;
        ELSIF x =- 3985 THEN
            tanh_f := - 1966;
        ELSIF x =- 3984 THEN
            tanh_f := - 1966;
        ELSIF x =- 3983 THEN
            tanh_f := - 1966;
        ELSIF x =- 3982 THEN
            tanh_f := - 1966;
        ELSIF x =- 3981 THEN
            tanh_f := - 1966;
        ELSIF x =- 3980 THEN
            tanh_f := - 1966;
        ELSIF x =- 3979 THEN
            tanh_f := - 1966;
        ELSIF x =- 3978 THEN
            tanh_f := - 1966;
        ELSIF x =- 3977 THEN
            tanh_f := - 1965;
        ELSIF x =- 3976 THEN
            tanh_f := - 1965;
        ELSIF x =- 3975 THEN
            tanh_f := - 1965;
        ELSIF x =- 3974 THEN
            tanh_f := - 1965;
        ELSIF x =- 3973 THEN
            tanh_f := - 1965;
        ELSIF x =- 3972 THEN
            tanh_f := - 1965;
        ELSIF x =- 3971 THEN
            tanh_f := - 1965;
        ELSIF x =- 3970 THEN
            tanh_f := - 1965;
        ELSIF x =- 3969 THEN
            tanh_f := - 1965;
        ELSIF x =- 3968 THEN
            tanh_f := - 1965;
        ELSIF x =- 3967 THEN
            tanh_f := - 1965;
        ELSIF x =- 3966 THEN
            tanh_f := - 1965;
        ELSIF x =- 3965 THEN
            tanh_f := - 1965;
        ELSIF x =- 3964 THEN
            tanh_f := - 1964;
        ELSIF x =- 3963 THEN
            tanh_f := - 1964;
        ELSIF x =- 3962 THEN
            tanh_f := - 1964;
        ELSIF x =- 3961 THEN
            tanh_f := - 1964;
        ELSIF x =- 3960 THEN
            tanh_f := - 1964;
        ELSIF x =- 3959 THEN
            tanh_f := - 1964;
        ELSIF x =- 3958 THEN
            tanh_f := - 1964;
        ELSIF x =- 3957 THEN
            tanh_f := - 1964;
        ELSIF x =- 3956 THEN
            tanh_f := - 1964;
        ELSIF x =- 3955 THEN
            tanh_f := - 1964;
        ELSIF x =- 3954 THEN
            tanh_f := - 1964;
        ELSIF x =- 3953 THEN
            tanh_f := - 1964;
        ELSIF x =- 3952 THEN
            tanh_f := - 1964;
        ELSIF x =- 3951 THEN
            tanh_f := - 1963;
        ELSIF x =- 3950 THEN
            tanh_f := - 1963;
        ELSIF x =- 3949 THEN
            tanh_f := - 1963;
        ELSIF x =- 3948 THEN
            tanh_f := - 1963;
        ELSIF x =- 3947 THEN
            tanh_f := - 1963;
        ELSIF x =- 3946 THEN
            tanh_f := - 1963;
        ELSIF x =- 3945 THEN
            tanh_f := - 1963;
        ELSIF x =- 3944 THEN
            tanh_f := - 1963;
        ELSIF x =- 3943 THEN
            tanh_f := - 1963;
        ELSIF x =- 3942 THEN
            tanh_f := - 1963;
        ELSIF x =- 3941 THEN
            tanh_f := - 1963;
        ELSIF x =- 3940 THEN
            tanh_f := - 1963;
        ELSIF x =- 3939 THEN
            tanh_f := - 1963;
        ELSIF x =- 3938 THEN
            tanh_f := - 1962;
        ELSIF x =- 3937 THEN
            tanh_f := - 1962;
        ELSIF x =- 3936 THEN
            tanh_f := - 1962;
        ELSIF x =- 3935 THEN
            tanh_f := - 1962;
        ELSIF x =- 3934 THEN
            tanh_f := - 1962;
        ELSIF x =- 3933 THEN
            tanh_f := - 1962;
        ELSIF x =- 3932 THEN
            tanh_f := - 1962;
        ELSIF x =- 3931 THEN
            tanh_f := - 1962;
        ELSIF x =- 3930 THEN
            tanh_f := - 1962;
        ELSIF x =- 3929 THEN
            tanh_f := - 1962;
        ELSIF x =- 3928 THEN
            tanh_f := - 1962;
        ELSIF x =- 3927 THEN
            tanh_f := - 1962;
        ELSIF x =- 3926 THEN
            tanh_f := - 1962;
        ELSIF x =- 3925 THEN
            tanh_f := - 1961;
        ELSIF x =- 3924 THEN
            tanh_f := - 1961;
        ELSIF x =- 3923 THEN
            tanh_f := - 1961;
        ELSIF x =- 3922 THEN
            tanh_f := - 1961;
        ELSIF x =- 3921 THEN
            tanh_f := - 1961;
        ELSIF x =- 3920 THEN
            tanh_f := - 1961;
        ELSIF x =- 3919 THEN
            tanh_f := - 1961;
        ELSIF x =- 3918 THEN
            tanh_f := - 1961;
        ELSIF x =- 3917 THEN
            tanh_f := - 1961;
        ELSIF x =- 3916 THEN
            tanh_f := - 1961;
        ELSIF x =- 3915 THEN
            tanh_f := - 1961;
        ELSIF x =- 3914 THEN
            tanh_f := - 1961;
        ELSIF x =- 3913 THEN
            tanh_f := - 1961;
        ELSIF x =- 3912 THEN
            tanh_f := - 1960;
        ELSIF x =- 3911 THEN
            tanh_f := - 1960;
        ELSIF x =- 3910 THEN
            tanh_f := - 1960;
        ELSIF x =- 3909 THEN
            tanh_f := - 1960;
        ELSIF x =- 3908 THEN
            tanh_f := - 1960;
        ELSIF x =- 3907 THEN
            tanh_f := - 1960;
        ELSIF x =- 3906 THEN
            tanh_f := - 1960;
        ELSIF x =- 3905 THEN
            tanh_f := - 1960;
        ELSIF x =- 3904 THEN
            tanh_f := - 1960;
        ELSIF x =- 3903 THEN
            tanh_f := - 1960;
        ELSIF x =- 3902 THEN
            tanh_f := - 1960;
        ELSIF x =- 3901 THEN
            tanh_f := - 1960;
        ELSIF x =- 3900 THEN
            tanh_f := - 1960;
        ELSIF x =- 3899 THEN
            tanh_f := - 1959;
        ELSIF x =- 3898 THEN
            tanh_f := - 1959;
        ELSIF x =- 3897 THEN
            tanh_f := - 1959;
        ELSIF x =- 3896 THEN
            tanh_f := - 1959;
        ELSIF x =- 3895 THEN
            tanh_f := - 1959;
        ELSIF x =- 3894 THEN
            tanh_f := - 1959;
        ELSIF x =- 3893 THEN
            tanh_f := - 1959;
        ELSIF x =- 3892 THEN
            tanh_f := - 1959;
        ELSIF x =- 3891 THEN
            tanh_f := - 1959;
        ELSIF x =- 3890 THEN
            tanh_f := - 1959;
        ELSIF x =- 3889 THEN
            tanh_f := - 1959;
        ELSIF x =- 3888 THEN
            tanh_f := - 1959;
        ELSIF x =- 3887 THEN
            tanh_f := - 1959;
        ELSIF x =- 3886 THEN
            tanh_f := - 1959;
        ELSIF x =- 3885 THEN
            tanh_f := - 1958;
        ELSIF x =- 3884 THEN
            tanh_f := - 1958;
        ELSIF x =- 3883 THEN
            tanh_f := - 1958;
        ELSIF x =- 3882 THEN
            tanh_f := - 1958;
        ELSIF x =- 3881 THEN
            tanh_f := - 1958;
        ELSIF x =- 3880 THEN
            tanh_f := - 1958;
        ELSIF x =- 3879 THEN
            tanh_f := - 1958;
        ELSIF x =- 3878 THEN
            tanh_f := - 1958;
        ELSIF x =- 3877 THEN
            tanh_f := - 1958;
        ELSIF x =- 3876 THEN
            tanh_f := - 1958;
        ELSIF x =- 3875 THEN
            tanh_f := - 1958;
        ELSIF x =- 3874 THEN
            tanh_f := - 1958;
        ELSIF x =- 3873 THEN
            tanh_f := - 1958;
        ELSIF x =- 3872 THEN
            tanh_f := - 1957;
        ELSIF x =- 3871 THEN
            tanh_f := - 1957;
        ELSIF x =- 3870 THEN
            tanh_f := - 1957;
        ELSIF x =- 3869 THEN
            tanh_f := - 1957;
        ELSIF x =- 3868 THEN
            tanh_f := - 1957;
        ELSIF x =- 3867 THEN
            tanh_f := - 1957;
        ELSIF x =- 3866 THEN
            tanh_f := - 1957;
        ELSIF x =- 3865 THEN
            tanh_f := - 1957;
        ELSIF x =- 3864 THEN
            tanh_f := - 1957;
        ELSIF x =- 3863 THEN
            tanh_f := - 1957;
        ELSIF x =- 3862 THEN
            tanh_f := - 1957;
        ELSIF x =- 3861 THEN
            tanh_f := - 1957;
        ELSIF x =- 3860 THEN
            tanh_f := - 1957;
        ELSIF x =- 3859 THEN
            tanh_f := - 1956;
        ELSIF x =- 3858 THEN
            tanh_f := - 1956;
        ELSIF x =- 3857 THEN
            tanh_f := - 1956;
        ELSIF x =- 3856 THEN
            tanh_f := - 1956;
        ELSIF x =- 3855 THEN
            tanh_f := - 1956;
        ELSIF x =- 3854 THEN
            tanh_f := - 1956;
        ELSIF x =- 3853 THEN
            tanh_f := - 1956;
        ELSIF x =- 3852 THEN
            tanh_f := - 1956;
        ELSIF x =- 3851 THEN
            tanh_f := - 1956;
        ELSIF x =- 3850 THEN
            tanh_f := - 1956;
        ELSIF x =- 3849 THEN
            tanh_f := - 1956;
        ELSIF x =- 3848 THEN
            tanh_f := - 1956;
        ELSIF x =- 3847 THEN
            tanh_f := - 1956;
        ELSIF x =- 3846 THEN
            tanh_f := - 1955;
        ELSIF x =- 3845 THEN
            tanh_f := - 1955;
        ELSIF x =- 3844 THEN
            tanh_f := - 1955;
        ELSIF x =- 3843 THEN
            tanh_f := - 1955;
        ELSIF x =- 3842 THEN
            tanh_f := - 1955;
        ELSIF x =- 3841 THEN
            tanh_f := - 1955;
        ELSIF x =- 3840 THEN
            tanh_f := - 1955;
        ELSIF x =- 3839 THEN
            tanh_f := - 1955;
        ELSIF x =- 3838 THEN
            tanh_f := - 1955;
        ELSIF x =- 3837 THEN
            tanh_f := - 1955;
        ELSIF x =- 3836 THEN
            tanh_f := - 1955;
        ELSIF x =- 3835 THEN
            tanh_f := - 1955;
        ELSIF x =- 3834 THEN
            tanh_f := - 1955;
        ELSIF x =- 3833 THEN
            tanh_f := - 1955;
        ELSIF x =- 3832 THEN
            tanh_f := - 1955;
        ELSIF x =- 3831 THEN
            tanh_f := - 1955;
        ELSIF x =- 3830 THEN
            tanh_f := - 1954;
        ELSIF x =- 3829 THEN
            tanh_f := - 1954;
        ELSIF x =- 3828 THEN
            tanh_f := - 1954;
        ELSIF x =- 3827 THEN
            tanh_f := - 1954;
        ELSIF x =- 3826 THEN
            tanh_f := - 1954;
        ELSIF x =- 3825 THEN
            tanh_f := - 1954;
        ELSIF x =- 3824 THEN
            tanh_f := - 1954;
        ELSIF x =- 3823 THEN
            tanh_f := - 1954;
        ELSIF x =- 3822 THEN
            tanh_f := - 1954;
        ELSIF x =- 3821 THEN
            tanh_f := - 1953;
        ELSIF x =- 3820 THEN
            tanh_f := - 1953;
        ELSIF x =- 3819 THEN
            tanh_f := - 1953;
        ELSIF x =- 3818 THEN
            tanh_f := - 1953;
        ELSIF x =- 3817 THEN
            tanh_f := - 1953;
        ELSIF x =- 3816 THEN
            tanh_f := - 1953;
        ELSIF x =- 3815 THEN
            tanh_f := - 1953;
        ELSIF x =- 3814 THEN
            tanh_f := - 1953;
        ELSIF x =- 3813 THEN
            tanh_f := - 1953;
        ELSIF x =- 3812 THEN
            tanh_f := - 1953;
        ELSIF x =- 3811 THEN
            tanh_f := - 1952;
        ELSIF x =- 3810 THEN
            tanh_f := - 1952;
        ELSIF x =- 3809 THEN
            tanh_f := - 1952;
        ELSIF x =- 3808 THEN
            tanh_f := - 1952;
        ELSIF x =- 3807 THEN
            tanh_f := - 1952;
        ELSIF x =- 3806 THEN
            tanh_f := - 1952;
        ELSIF x =- 3805 THEN
            tanh_f := - 1952;
        ELSIF x =- 3804 THEN
            tanh_f := - 1952;
        ELSIF x =- 3803 THEN
            tanh_f := - 1952;
        ELSIF x =- 3802 THEN
            tanh_f := - 1951;
        ELSIF x =- 3801 THEN
            tanh_f := - 1951;
        ELSIF x =- 3800 THEN
            tanh_f := - 1951;
        ELSIF x =- 3799 THEN
            tanh_f := - 1951;
        ELSIF x =- 3798 THEN
            tanh_f := - 1951;
        ELSIF x =- 3797 THEN
            tanh_f := - 1951;
        ELSIF x =- 3796 THEN
            tanh_f := - 1951;
        ELSIF x =- 3795 THEN
            tanh_f := - 1951;
        ELSIF x =- 3794 THEN
            tanh_f := - 1951;
        ELSIF x =- 3793 THEN
            tanh_f := - 1951;
        ELSIF x =- 3792 THEN
            tanh_f := - 1950;
        ELSIF x =- 3791 THEN
            tanh_f := - 1950;
        ELSIF x =- 3790 THEN
            tanh_f := - 1950;
        ELSIF x =- 3789 THEN
            tanh_f := - 1950;
        ELSIF x =- 3788 THEN
            tanh_f := - 1950;
        ELSIF x =- 3787 THEN
            tanh_f := - 1950;
        ELSIF x =- 3786 THEN
            tanh_f := - 1950;
        ELSIF x =- 3785 THEN
            tanh_f := - 1950;
        ELSIF x =- 3784 THEN
            tanh_f := - 1950;
        ELSIF x =- 3783 THEN
            tanh_f := - 1949;
        ELSIF x =- 3782 THEN
            tanh_f := - 1949;
        ELSIF x =- 3781 THEN
            tanh_f := - 1949;
        ELSIF x =- 3780 THEN
            tanh_f := - 1949;
        ELSIF x =- 3779 THEN
            tanh_f := - 1949;
        ELSIF x =- 3778 THEN
            tanh_f := - 1949;
        ELSIF x =- 3777 THEN
            tanh_f := - 1949;
        ELSIF x =- 3776 THEN
            tanh_f := - 1949;
        ELSIF x =- 3775 THEN
            tanh_f := - 1949;
        ELSIF x =- 3774 THEN
            tanh_f := - 1949;
        ELSIF x =- 3773 THEN
            tanh_f := - 1948;
        ELSIF x =- 3772 THEN
            tanh_f := - 1948;
        ELSIF x =- 3771 THEN
            tanh_f := - 1948;
        ELSIF x =- 3770 THEN
            tanh_f := - 1948;
        ELSIF x =- 3769 THEN
            tanh_f := - 1948;
        ELSIF x =- 3768 THEN
            tanh_f := - 1948;
        ELSIF x =- 3767 THEN
            tanh_f := - 1948;
        ELSIF x =- 3766 THEN
            tanh_f := - 1948;
        ELSIF x =- 3765 THEN
            tanh_f := - 1948;
        ELSIF x =- 3764 THEN
            tanh_f := - 1947;
        ELSIF x =- 3763 THEN
            tanh_f := - 1947;
        ELSIF x =- 3762 THEN
            tanh_f := - 1947;
        ELSIF x =- 3761 THEN
            tanh_f := - 1947;
        ELSIF x =- 3760 THEN
            tanh_f := - 1947;
        ELSIF x =- 3759 THEN
            tanh_f := - 1947;
        ELSIF x =- 3758 THEN
            tanh_f := - 1947;
        ELSIF x =- 3757 THEN
            tanh_f := - 1947;
        ELSIF x =- 3756 THEN
            tanh_f := - 1947;
        ELSIF x =- 3755 THEN
            tanh_f := - 1947;
        ELSIF x =- 3754 THEN
            tanh_f := - 1946;
        ELSIF x =- 3753 THEN
            tanh_f := - 1946;
        ELSIF x =- 3752 THEN
            tanh_f := - 1946;
        ELSIF x =- 3751 THEN
            tanh_f := - 1946;
        ELSIF x =- 3750 THEN
            tanh_f := - 1946;
        ELSIF x =- 3749 THEN
            tanh_f := - 1946;
        ELSIF x =- 3748 THEN
            tanh_f := - 1946;
        ELSIF x =- 3747 THEN
            tanh_f := - 1946;
        ELSIF x =- 3746 THEN
            tanh_f := - 1946;
        ELSIF x =- 3745 THEN
            tanh_f := - 1945;
        ELSIF x =- 3744 THEN
            tanh_f := - 1945;
        ELSIF x =- 3743 THEN
            tanh_f := - 1945;
        ELSIF x =- 3742 THEN
            tanh_f := - 1945;
        ELSIF x =- 3741 THEN
            tanh_f := - 1945;
        ELSIF x =- 3740 THEN
            tanh_f := - 1945;
        ELSIF x =- 3739 THEN
            tanh_f := - 1945;
        ELSIF x =- 3738 THEN
            tanh_f := - 1945;
        ELSIF x =- 3737 THEN
            tanh_f := - 1945;
        ELSIF x =- 3736 THEN
            tanh_f := - 1945;
        ELSIF x =- 3735 THEN
            tanh_f := - 1944;
        ELSIF x =- 3734 THEN
            tanh_f := - 1944;
        ELSIF x =- 3733 THEN
            tanh_f := - 1944;
        ELSIF x =- 3732 THEN
            tanh_f := - 1944;
        ELSIF x =- 3731 THEN
            tanh_f := - 1944;
        ELSIF x =- 3730 THEN
            tanh_f := - 1944;
        ELSIF x =- 3729 THEN
            tanh_f := - 1944;
        ELSIF x =- 3728 THEN
            tanh_f := - 1944;
        ELSIF x =- 3727 THEN
            tanh_f := - 1944;
        ELSIF x =- 3726 THEN
            tanh_f := - 1943;
        ELSIF x =- 3725 THEN
            tanh_f := - 1943;
        ELSIF x =- 3724 THEN
            tanh_f := - 1943;
        ELSIF x =- 3723 THEN
            tanh_f := - 1943;
        ELSIF x =- 3722 THEN
            tanh_f := - 1943;
        ELSIF x =- 3721 THEN
            tanh_f := - 1943;
        ELSIF x =- 3720 THEN
            tanh_f := - 1943;
        ELSIF x =- 3719 THEN
            tanh_f := - 1943;
        ELSIF x =- 3718 THEN
            tanh_f := - 1943;
        ELSIF x =- 3717 THEN
            tanh_f := - 1943;
        ELSIF x =- 3716 THEN
            tanh_f := - 1942;
        ELSIF x =- 3715 THEN
            tanh_f := - 1942;
        ELSIF x =- 3714 THEN
            tanh_f := - 1942;
        ELSIF x =- 3713 THEN
            tanh_f := - 1942;
        ELSIF x =- 3712 THEN
            tanh_f := - 1942;
        ELSIF x =- 3711 THEN
            tanh_f := - 1942;
        ELSIF x =- 3710 THEN
            tanh_f := - 1942;
        ELSIF x =- 3709 THEN
            tanh_f := - 1942;
        ELSIF x =- 3708 THEN
            tanh_f := - 1942;
        ELSIF x =- 3707 THEN
            tanh_f := - 1941;
        ELSIF x =- 3706 THEN
            tanh_f := - 1941;
        ELSIF x =- 3705 THEN
            tanh_f := - 1941;
        ELSIF x =- 3704 THEN
            tanh_f := - 1941;
        ELSIF x =- 3703 THEN
            tanh_f := - 1941;
        ELSIF x =- 3702 THEN
            tanh_f := - 1941;
        ELSIF x =- 3701 THEN
            tanh_f := - 1941;
        ELSIF x =- 3700 THEN
            tanh_f := - 1941;
        ELSIF x =- 3699 THEN
            tanh_f := - 1941;
        ELSIF x =- 3698 THEN
            tanh_f := - 1941;
        ELSIF x =- 3697 THEN
            tanh_f := - 1940;
        ELSIF x =- 3696 THEN
            tanh_f := - 1940;
        ELSIF x =- 3695 THEN
            tanh_f := - 1940;
        ELSIF x =- 3694 THEN
            tanh_f := - 1940;
        ELSIF x =- 3693 THEN
            tanh_f := - 1940;
        ELSIF x =- 3692 THEN
            tanh_f := - 1940;
        ELSIF x =- 3691 THEN
            tanh_f := - 1940;
        ELSIF x =- 3690 THEN
            tanh_f := - 1940;
        ELSIF x =- 3689 THEN
            tanh_f := - 1940;
        ELSIF x =- 3688 THEN
            tanh_f := - 1939;
        ELSIF x =- 3687 THEN
            tanh_f := - 1939;
        ELSIF x =- 3686 THEN
            tanh_f := - 1939;
        ELSIF x =- 3685 THEN
            tanh_f := - 1939;
        ELSIF x =- 3684 THEN
            tanh_f := - 1939;
        ELSIF x =- 3683 THEN
            tanh_f := - 1939;
        ELSIF x =- 3682 THEN
            tanh_f := - 1939;
        ELSIF x =- 3681 THEN
            tanh_f := - 1939;
        ELSIF x =- 3680 THEN
            tanh_f := - 1939;
        ELSIF x =- 3679 THEN
            tanh_f := - 1939;
        ELSIF x =- 3678 THEN
            tanh_f := - 1938;
        ELSIF x =- 3677 THEN
            tanh_f := - 1938;
        ELSIF x =- 3676 THEN
            tanh_f := - 1938;
        ELSIF x =- 3675 THEN
            tanh_f := - 1938;
        ELSIF x =- 3674 THEN
            tanh_f := - 1938;
        ELSIF x =- 3673 THEN
            tanh_f := - 1938;
        ELSIF x =- 3672 THEN
            tanh_f := - 1938;
        ELSIF x =- 3671 THEN
            tanh_f := - 1938;
        ELSIF x =- 3670 THEN
            tanh_f := - 1938;
        ELSIF x =- 3669 THEN
            tanh_f := - 1937;
        ELSIF x =- 3668 THEN
            tanh_f := - 1937;
        ELSIF x =- 3667 THEN
            tanh_f := - 1937;
        ELSIF x =- 3666 THEN
            tanh_f := - 1937;
        ELSIF x =- 3665 THEN
            tanh_f := - 1937;
        ELSIF x =- 3664 THEN
            tanh_f := - 1937;
        ELSIF x =- 3663 THEN
            tanh_f := - 1937;
        ELSIF x =- 3662 THEN
            tanh_f := - 1937;
        ELSIF x =- 3661 THEN
            tanh_f := - 1937;
        ELSIF x =- 3660 THEN
            tanh_f := - 1937;
        ELSIF x =- 3659 THEN
            tanh_f := - 1936;
        ELSIF x =- 3658 THEN
            tanh_f := - 1936;
        ELSIF x =- 3657 THEN
            tanh_f := - 1936;
        ELSIF x =- 3656 THEN
            tanh_f := - 1936;
        ELSIF x =- 3655 THEN
            tanh_f := - 1936;
        ELSIF x =- 3654 THEN
            tanh_f := - 1936;
        ELSIF x =- 3653 THEN
            tanh_f := - 1936;
        ELSIF x =- 3652 THEN
            tanh_f := - 1936;
        ELSIF x =- 3651 THEN
            tanh_f := - 1936;
        ELSIF x =- 3650 THEN
            tanh_f := - 1935;
        ELSIF x =- 3649 THEN
            tanh_f := - 1935;
        ELSIF x =- 3648 THEN
            tanh_f := - 1935;
        ELSIF x =- 3647 THEN
            tanh_f := - 1935;
        ELSIF x =- 3646 THEN
            tanh_f := - 1935;
        ELSIF x =- 3645 THEN
            tanh_f := - 1935;
        ELSIF x =- 3644 THEN
            tanh_f := - 1935;
        ELSIF x =- 3643 THEN
            tanh_f := - 1935;
        ELSIF x =- 3642 THEN
            tanh_f := - 1935;
        ELSIF x =- 3641 THEN
            tanh_f := - 1935;
        ELSIF x =- 3640 THEN
            tanh_f := - 1934;
        ELSIF x =- 3639 THEN
            tanh_f := - 1934;
        ELSIF x =- 3638 THEN
            tanh_f := - 1934;
        ELSIF x =- 3637 THEN
            tanh_f := - 1934;
        ELSIF x =- 3636 THEN
            tanh_f := - 1934;
        ELSIF x =- 3635 THEN
            tanh_f := - 1934;
        ELSIF x =- 3634 THEN
            tanh_f := - 1934;
        ELSIF x =- 3633 THEN
            tanh_f := - 1934;
        ELSIF x =- 3632 THEN
            tanh_f := - 1934;
        ELSIF x =- 3631 THEN
            tanh_f := - 1933;
        ELSIF x =- 3630 THEN
            tanh_f := - 1933;
        ELSIF x =- 3629 THEN
            tanh_f := - 1933;
        ELSIF x =- 3628 THEN
            tanh_f := - 1933;
        ELSIF x =- 3627 THEN
            tanh_f := - 1933;
        ELSIF x =- 3626 THEN
            tanh_f := - 1933;
        ELSIF x =- 3625 THEN
            tanh_f := - 1933;
        ELSIF x =- 3624 THEN
            tanh_f := - 1933;
        ELSIF x =- 3623 THEN
            tanh_f := - 1933;
        ELSIF x =- 3622 THEN
            tanh_f := - 1933;
        ELSIF x =- 3621 THEN
            tanh_f := - 1932;
        ELSIF x =- 3620 THEN
            tanh_f := - 1932;
        ELSIF x =- 3619 THEN
            tanh_f := - 1932;
        ELSIF x =- 3618 THEN
            tanh_f := - 1932;
        ELSIF x =- 3617 THEN
            tanh_f := - 1932;
        ELSIF x =- 3616 THEN
            tanh_f := - 1932;
        ELSIF x =- 3615 THEN
            tanh_f := - 1932;
        ELSIF x =- 3614 THEN
            tanh_f := - 1932;
        ELSIF x =- 3613 THEN
            tanh_f := - 1932;
        ELSIF x =- 3612 THEN
            tanh_f := - 1931;
        ELSIF x =- 3611 THEN
            tanh_f := - 1931;
        ELSIF x =- 3610 THEN
            tanh_f := - 1931;
        ELSIF x =- 3609 THEN
            tanh_f := - 1931;
        ELSIF x =- 3608 THEN
            tanh_f := - 1931;
        ELSIF x =- 3607 THEN
            tanh_f := - 1931;
        ELSIF x =- 3606 THEN
            tanh_f := - 1931;
        ELSIF x =- 3605 THEN
            tanh_f := - 1931;
        ELSIF x =- 3604 THEN
            tanh_f := - 1931;
        ELSIF x =- 3603 THEN
            tanh_f := - 1931;
        ELSIF x =- 3602 THEN
            tanh_f := - 1930;
        ELSIF x =- 3601 THEN
            tanh_f := - 1930;
        ELSIF x =- 3600 THEN
            tanh_f := - 1930;
        ELSIF x =- 3599 THEN
            tanh_f := - 1930;
        ELSIF x =- 3598 THEN
            tanh_f := - 1930;
        ELSIF x =- 3597 THEN
            tanh_f := - 1930;
        ELSIF x =- 3596 THEN
            tanh_f := - 1930;
        ELSIF x =- 3595 THEN
            tanh_f := - 1930;
        ELSIF x =- 3594 THEN
            tanh_f := - 1930;
        ELSIF x =- 3593 THEN
            tanh_f := - 1929;
        ELSIF x =- 3592 THEN
            tanh_f := - 1929;
        ELSIF x =- 3591 THEN
            tanh_f := - 1929;
        ELSIF x =- 3590 THEN
            tanh_f := - 1929;
        ELSIF x =- 3589 THEN
            tanh_f := - 1929;
        ELSIF x =- 3588 THEN
            tanh_f := - 1929;
        ELSIF x =- 3587 THEN
            tanh_f := - 1929;
        ELSIF x =- 3586 THEN
            tanh_f := - 1929;
        ELSIF x =- 3585 THEN
            tanh_f := - 1929;
        ELSIF x =- 3584 THEN
            tanh_f := - 1928;
        ELSIF x =- 3583 THEN
            tanh_f := - 1928;
        ELSIF x =- 3582 THEN
            tanh_f := - 1928;
        ELSIF x =- 3581 THEN
            tanh_f := - 1928;
        ELSIF x =- 3580 THEN
            tanh_f := - 1928;
        ELSIF x =- 3579 THEN
            tanh_f := - 1928;
        ELSIF x =- 3578 THEN
            tanh_f := - 1928;
        ELSIF x =- 3577 THEN
            tanh_f := - 1928;
        ELSIF x =- 3576 THEN
            tanh_f := - 1927;
        ELSIF x =- 3575 THEN
            tanh_f := - 1927;
        ELSIF x =- 3574 THEN
            tanh_f := - 1927;
        ELSIF x =- 3573 THEN
            tanh_f := - 1927;
        ELSIF x =- 3572 THEN
            tanh_f := - 1927;
        ELSIF x =- 3571 THEN
            tanh_f := - 1927;
        ELSIF x =- 3570 THEN
            tanh_f := - 1927;
        ELSIF x =- 3569 THEN
            tanh_f := - 1927;
        ELSIF x =- 3568 THEN
            tanh_f := - 1926;
        ELSIF x =- 3567 THEN
            tanh_f := - 1926;
        ELSIF x =- 3566 THEN
            tanh_f := - 1926;
        ELSIF x =- 3565 THEN
            tanh_f := - 1926;
        ELSIF x =- 3564 THEN
            tanh_f := - 1926;
        ELSIF x =- 3563 THEN
            tanh_f := - 1926;
        ELSIF x =- 3562 THEN
            tanh_f := - 1926;
        ELSIF x =- 3561 THEN
            tanh_f := - 1926;
        ELSIF x =- 3560 THEN
            tanh_f := - 1925;
        ELSIF x =- 3559 THEN
            tanh_f := - 1925;
        ELSIF x =- 3558 THEN
            tanh_f := - 1925;
        ELSIF x =- 3557 THEN
            tanh_f := - 1925;
        ELSIF x =- 3556 THEN
            tanh_f := - 1925;
        ELSIF x =- 3555 THEN
            tanh_f := - 1925;
        ELSIF x =- 3554 THEN
            tanh_f := - 1925;
        ELSIF x =- 3553 THEN
            tanh_f := - 1925;
        ELSIF x =- 3552 THEN
            tanh_f := - 1924;
        ELSIF x =- 3551 THEN
            tanh_f := - 1924;
        ELSIF x =- 3550 THEN
            tanh_f := - 1924;
        ELSIF x =- 3549 THEN
            tanh_f := - 1924;
        ELSIF x =- 3548 THEN
            tanh_f := - 1924;
        ELSIF x =- 3547 THEN
            tanh_f := - 1924;
        ELSIF x =- 3546 THEN
            tanh_f := - 1924;
        ELSIF x =- 3545 THEN
            tanh_f := - 1924;
        ELSIF x =- 3544 THEN
            tanh_f := - 1923;
        ELSIF x =- 3543 THEN
            tanh_f := - 1923;
        ELSIF x =- 3542 THEN
            tanh_f := - 1923;
        ELSIF x =- 3541 THEN
            tanh_f := - 1923;
        ELSIF x =- 3540 THEN
            tanh_f := - 1923;
        ELSIF x =- 3539 THEN
            tanh_f := - 1923;
        ELSIF x =- 3538 THEN
            tanh_f := - 1923;
        ELSIF x =- 3537 THEN
            tanh_f := - 1923;
        ELSIF x =- 3536 THEN
            tanh_f := - 1922;
        ELSIF x =- 3535 THEN
            tanh_f := - 1922;
        ELSIF x =- 3534 THEN
            tanh_f := - 1922;
        ELSIF x =- 3533 THEN
            tanh_f := - 1922;
        ELSIF x =- 3532 THEN
            tanh_f := - 1922;
        ELSIF x =- 3531 THEN
            tanh_f := - 1922;
        ELSIF x =- 3530 THEN
            tanh_f := - 1922;
        ELSIF x =- 3529 THEN
            tanh_f := - 1922;
        ELSIF x =- 3528 THEN
            tanh_f := - 1921;
        ELSIF x =- 3527 THEN
            tanh_f := - 1921;
        ELSIF x =- 3526 THEN
            tanh_f := - 1921;
        ELSIF x =- 3525 THEN
            tanh_f := - 1921;
        ELSIF x =- 3524 THEN
            tanh_f := - 1921;
        ELSIF x =- 3523 THEN
            tanh_f := - 1921;
        ELSIF x =- 3522 THEN
            tanh_f := - 1921;
        ELSIF x =- 3521 THEN
            tanh_f := - 1921;
        ELSIF x =- 3520 THEN
            tanh_f := - 1920;
        ELSIF x =- 3519 THEN
            tanh_f := - 1920;
        ELSIF x =- 3518 THEN
            tanh_f := - 1920;
        ELSIF x =- 3517 THEN
            tanh_f := - 1920;
        ELSIF x =- 3516 THEN
            tanh_f := - 1920;
        ELSIF x =- 3515 THEN
            tanh_f := - 1920;
        ELSIF x =- 3514 THEN
            tanh_f := - 1920;
        ELSIF x =- 3513 THEN
            tanh_f := - 1920;
        ELSIF x =- 3512 THEN
            tanh_f := - 1919;
        ELSIF x =- 3511 THEN
            tanh_f := - 1919;
        ELSIF x =- 3510 THEN
            tanh_f := - 1919;
        ELSIF x =- 3509 THEN
            tanh_f := - 1919;
        ELSIF x =- 3508 THEN
            tanh_f := - 1919;
        ELSIF x =- 3507 THEN
            tanh_f := - 1919;
        ELSIF x =- 3506 THEN
            tanh_f := - 1919;
        ELSIF x =- 3505 THEN
            tanh_f := - 1919;
        ELSIF x =- 3504 THEN
            tanh_f := - 1918;
        ELSIF x =- 3503 THEN
            tanh_f := - 1918;
        ELSIF x =- 3502 THEN
            tanh_f := - 1918;
        ELSIF x =- 3501 THEN
            tanh_f := - 1918;
        ELSIF x =- 3500 THEN
            tanh_f := - 1918;
        ELSIF x =- 3499 THEN
            tanh_f := - 1918;
        ELSIF x =- 3498 THEN
            tanh_f := - 1918;
        ELSIF x =- 3497 THEN
            tanh_f := - 1918;
        ELSIF x =- 3496 THEN
            tanh_f := - 1917;
        ELSIF x =- 3495 THEN
            tanh_f := - 1917;
        ELSIF x =- 3494 THEN
            tanh_f := - 1917;
        ELSIF x =- 3493 THEN
            tanh_f := - 1917;
        ELSIF x =- 3492 THEN
            tanh_f := - 1917;
        ELSIF x =- 3491 THEN
            tanh_f := - 1917;
        ELSIF x =- 3490 THEN
            tanh_f := - 1917;
        ELSIF x =- 3489 THEN
            tanh_f := - 1917;
        ELSIF x =- 3488 THEN
            tanh_f := - 1916;
        ELSIF x =- 3487 THEN
            tanh_f := - 1916;
        ELSIF x =- 3486 THEN
            tanh_f := - 1916;
        ELSIF x =- 3485 THEN
            tanh_f := - 1916;
        ELSIF x =- 3484 THEN
            tanh_f := - 1916;
        ELSIF x =- 3483 THEN
            tanh_f := - 1916;
        ELSIF x =- 3482 THEN
            tanh_f := - 1916;
        ELSIF x =- 3481 THEN
            tanh_f := - 1916;
        ELSIF x =- 3480 THEN
            tanh_f := - 1915;
        ELSIF x =- 3479 THEN
            tanh_f := - 1915;
        ELSIF x =- 3478 THEN
            tanh_f := - 1915;
        ELSIF x =- 3477 THEN
            tanh_f := - 1915;
        ELSIF x =- 3476 THEN
            tanh_f := - 1915;
        ELSIF x =- 3475 THEN
            tanh_f := - 1915;
        ELSIF x =- 3474 THEN
            tanh_f := - 1915;
        ELSIF x =- 3473 THEN
            tanh_f := - 1915;
        ELSIF x =- 3472 THEN
            tanh_f := - 1914;
        ELSIF x =- 3471 THEN
            tanh_f := - 1914;
        ELSIF x =- 3470 THEN
            tanh_f := - 1914;
        ELSIF x =- 3469 THEN
            tanh_f := - 1914;
        ELSIF x =- 3468 THEN
            tanh_f := - 1914;
        ELSIF x =- 3467 THEN
            tanh_f := - 1914;
        ELSIF x =- 3466 THEN
            tanh_f := - 1914;
        ELSIF x =- 3465 THEN
            tanh_f := - 1914;
        ELSIF x =- 3464 THEN
            tanh_f := - 1913;
        ELSIF x =- 3463 THEN
            tanh_f := - 1913;
        ELSIF x =- 3462 THEN
            tanh_f := - 1913;
        ELSIF x =- 3461 THEN
            tanh_f := - 1913;
        ELSIF x =- 3460 THEN
            tanh_f := - 1913;
        ELSIF x =- 3459 THEN
            tanh_f := - 1913;
        ELSIF x =- 3458 THEN
            tanh_f := - 1913;
        ELSIF x =- 3457 THEN
            tanh_f := - 1913;
        ELSIF x =- 3456 THEN
            tanh_f := - 1912;
        ELSIF x =- 3455 THEN
            tanh_f := - 1912;
        ELSIF x =- 3454 THEN
            tanh_f := - 1912;
        ELSIF x =- 3453 THEN
            tanh_f := - 1912;
        ELSIF x =- 3452 THEN
            tanh_f := - 1912;
        ELSIF x =- 3451 THEN
            tanh_f := - 1912;
        ELSIF x =- 3450 THEN
            tanh_f := - 1912;
        ELSIF x =- 3449 THEN
            tanh_f := - 1912;
        ELSIF x =- 3448 THEN
            tanh_f := - 1911;
        ELSIF x =- 3447 THEN
            tanh_f := - 1911;
        ELSIF x =- 3446 THEN
            tanh_f := - 1911;
        ELSIF x =- 3445 THEN
            tanh_f := - 1911;
        ELSIF x =- 3444 THEN
            tanh_f := - 1911;
        ELSIF x =- 3443 THEN
            tanh_f := - 1911;
        ELSIF x =- 3442 THEN
            tanh_f := - 1911;
        ELSIF x =- 3441 THEN
            tanh_f := - 1911;
        ELSIF x =- 3440 THEN
            tanh_f := - 1910;
        ELSIF x =- 3439 THEN
            tanh_f := - 1910;
        ELSIF x =- 3438 THEN
            tanh_f := - 1910;
        ELSIF x =- 3437 THEN
            tanh_f := - 1910;
        ELSIF x =- 3436 THEN
            tanh_f := - 1910;
        ELSIF x =- 3435 THEN
            tanh_f := - 1910;
        ELSIF x =- 3434 THEN
            tanh_f := - 1910;
        ELSIF x =- 3433 THEN
            tanh_f := - 1910;
        ELSIF x =- 3432 THEN
            tanh_f := - 1909;
        ELSIF x =- 3431 THEN
            tanh_f := - 1909;
        ELSIF x =- 3430 THEN
            tanh_f := - 1909;
        ELSIF x =- 3429 THEN
            tanh_f := - 1909;
        ELSIF x =- 3428 THEN
            tanh_f := - 1909;
        ELSIF x =- 3427 THEN
            tanh_f := - 1909;
        ELSIF x =- 3426 THEN
            tanh_f := - 1909;
        ELSIF x =- 3425 THEN
            tanh_f := - 1909;
        ELSIF x =- 3424 THEN
            tanh_f := - 1908;
        ELSIF x =- 3423 THEN
            tanh_f := - 1908;
        ELSIF x =- 3422 THEN
            tanh_f := - 1908;
        ELSIF x =- 3421 THEN
            tanh_f := - 1908;
        ELSIF x =- 3420 THEN
            tanh_f := - 1908;
        ELSIF x =- 3419 THEN
            tanh_f := - 1908;
        ELSIF x =- 3418 THEN
            tanh_f := - 1908;
        ELSIF x =- 3417 THEN
            tanh_f := - 1908;
        ELSIF x =- 3416 THEN
            tanh_f := - 1907;
        ELSIF x =- 3415 THEN
            tanh_f := - 1907;
        ELSIF x =- 3414 THEN
            tanh_f := - 1907;
        ELSIF x =- 3413 THEN
            tanh_f := - 1907;
        ELSIF x =- 3412 THEN
            tanh_f := - 1907;
        ELSIF x =- 3411 THEN
            tanh_f := - 1907;
        ELSIF x =- 3410 THEN
            tanh_f := - 1907;
        ELSIF x =- 3409 THEN
            tanh_f := - 1907;
        ELSIF x =- 3408 THEN
            tanh_f := - 1906;
        ELSIF x =- 3407 THEN
            tanh_f := - 1906;
        ELSIF x =- 3406 THEN
            tanh_f := - 1906;
        ELSIF x =- 3405 THEN
            tanh_f := - 1906;
        ELSIF x =- 3404 THEN
            tanh_f := - 1906;
        ELSIF x =- 3403 THEN
            tanh_f := - 1906;
        ELSIF x =- 3402 THEN
            tanh_f := - 1906;
        ELSIF x =- 3401 THEN
            tanh_f := - 1906;
        ELSIF x =- 3400 THEN
            tanh_f := - 1905;
        ELSIF x =- 3399 THEN
            tanh_f := - 1905;
        ELSIF x =- 3398 THEN
            tanh_f := - 1905;
        ELSIF x =- 3397 THEN
            tanh_f := - 1905;
        ELSIF x =- 3396 THEN
            tanh_f := - 1905;
        ELSIF x =- 3395 THEN
            tanh_f := - 1905;
        ELSIF x =- 3394 THEN
            tanh_f := - 1905;
        ELSIF x =- 3393 THEN
            tanh_f := - 1905;
        ELSIF x =- 3392 THEN
            tanh_f := - 1904;
        ELSIF x =- 3391 THEN
            tanh_f := - 1904;
        ELSIF x =- 3390 THEN
            tanh_f := - 1904;
        ELSIF x =- 3389 THEN
            tanh_f := - 1904;
        ELSIF x =- 3388 THEN
            tanh_f := - 1904;
        ELSIF x =- 3387 THEN
            tanh_f := - 1904;
        ELSIF x =- 3386 THEN
            tanh_f := - 1904;
        ELSIF x =- 3385 THEN
            tanh_f := - 1904;
        ELSIF x =- 3384 THEN
            tanh_f := - 1903;
        ELSIF x =- 3383 THEN
            tanh_f := - 1903;
        ELSIF x =- 3382 THEN
            tanh_f := - 1903;
        ELSIF x =- 3381 THEN
            tanh_f := - 1903;
        ELSIF x =- 3380 THEN
            tanh_f := - 1903;
        ELSIF x =- 3379 THEN
            tanh_f := - 1903;
        ELSIF x =- 3378 THEN
            tanh_f := - 1903;
        ELSIF x =- 3377 THEN
            tanh_f := - 1903;
        ELSIF x =- 3376 THEN
            tanh_f := - 1902;
        ELSIF x =- 3375 THEN
            tanh_f := - 1902;
        ELSIF x =- 3374 THEN
            tanh_f := - 1902;
        ELSIF x =- 3373 THEN
            tanh_f := - 1902;
        ELSIF x =- 3372 THEN
            tanh_f := - 1902;
        ELSIF x =- 3371 THEN
            tanh_f := - 1902;
        ELSIF x =- 3370 THEN
            tanh_f := - 1902;
        ELSIF x =- 3369 THEN
            tanh_f := - 1902;
        ELSIF x =- 3368 THEN
            tanh_f := - 1901;
        ELSIF x =- 3367 THEN
            tanh_f := - 1901;
        ELSIF x =- 3366 THEN
            tanh_f := - 1901;
        ELSIF x =- 3365 THEN
            tanh_f := - 1901;
        ELSIF x =- 3364 THEN
            tanh_f := - 1901;
        ELSIF x =- 3363 THEN
            tanh_f := - 1901;
        ELSIF x =- 3362 THEN
            tanh_f := - 1901;
        ELSIF x =- 3361 THEN
            tanh_f := - 1901;
        ELSIF x =- 3360 THEN
            tanh_f := - 1900;
        ELSIF x =- 3359 THEN
            tanh_f := - 1900;
        ELSIF x =- 3358 THEN
            tanh_f := - 1900;
        ELSIF x =- 3357 THEN
            tanh_f := - 1900;
        ELSIF x =- 3356 THEN
            tanh_f := - 1900;
        ELSIF x =- 3355 THEN
            tanh_f := - 1900;
        ELSIF x =- 3354 THEN
            tanh_f := - 1900;
        ELSIF x =- 3353 THEN
            tanh_f := - 1900;
        ELSIF x =- 3352 THEN
            tanh_f := - 1899;
        ELSIF x =- 3351 THEN
            tanh_f := - 1899;
        ELSIF x =- 3350 THEN
            tanh_f := - 1899;
        ELSIF x =- 3349 THEN
            tanh_f := - 1899;
        ELSIF x =- 3348 THEN
            tanh_f := - 1899;
        ELSIF x =- 3347 THEN
            tanh_f := - 1899;
        ELSIF x =- 3346 THEN
            tanh_f := - 1899;
        ELSIF x =- 3345 THEN
            tanh_f := - 1899;
        ELSIF x =- 3344 THEN
            tanh_f := - 1898;
        ELSIF x =- 3343 THEN
            tanh_f := - 1898;
        ELSIF x =- 3342 THEN
            tanh_f := - 1898;
        ELSIF x =- 3341 THEN
            tanh_f := - 1898;
        ELSIF x =- 3340 THEN
            tanh_f := - 1898;
        ELSIF x =- 3339 THEN
            tanh_f := - 1898;
        ELSIF x =- 3338 THEN
            tanh_f := - 1898;
        ELSIF x =- 3337 THEN
            tanh_f := - 1898;
        ELSIF x =- 3336 THEN
            tanh_f := - 1897;
        ELSIF x =- 3335 THEN
            tanh_f := - 1897;
        ELSIF x =- 3334 THEN
            tanh_f := - 1897;
        ELSIF x =- 3333 THEN
            tanh_f := - 1897;
        ELSIF x =- 3332 THEN
            tanh_f := - 1897;
        ELSIF x =- 3331 THEN
            tanh_f := - 1897;
        ELSIF x =- 3330 THEN
            tanh_f := - 1897;
        ELSIF x =- 3329 THEN
            tanh_f := - 1897;
        ELSIF x =- 3328 THEN
            tanh_f := - 1896;
        ELSIF x =- 3327 THEN
            tanh_f := - 1896;
        ELSIF x =- 3326 THEN
            tanh_f := - 1896;
        ELSIF x =- 3325 THEN
            tanh_f := - 1896;
        ELSIF x =- 3324 THEN
            tanh_f := - 1896;
        ELSIF x =- 3323 THEN
            tanh_f := - 1896;
        ELSIF x =- 3322 THEN
            tanh_f := - 1896;
        ELSIF x =- 3321 THEN
            tanh_f := - 1895;
        ELSIF x =- 3320 THEN
            tanh_f := - 1895;
        ELSIF x =- 3319 THEN
            tanh_f := - 1895;
        ELSIF x =- 3318 THEN
            tanh_f := - 1895;
        ELSIF x =- 3317 THEN
            tanh_f := - 1895;
        ELSIF x =- 3316 THEN
            tanh_f := - 1895;
        ELSIF x =- 3315 THEN
            tanh_f := - 1894;
        ELSIF x =- 3314 THEN
            tanh_f := - 1894;
        ELSIF x =- 3313 THEN
            tanh_f := - 1894;
        ELSIF x =- 3312 THEN
            tanh_f := - 1894;
        ELSIF x =- 3311 THEN
            tanh_f := - 1894;
        ELSIF x =- 3310 THEN
            tanh_f := - 1894;
        ELSIF x =- 3309 THEN
            tanh_f := - 1893;
        ELSIF x =- 3308 THEN
            tanh_f := - 1893;
        ELSIF x =- 3307 THEN
            tanh_f := - 1893;
        ELSIF x =- 3306 THEN
            tanh_f := - 1893;
        ELSIF x =- 3305 THEN
            tanh_f := - 1893;
        ELSIF x =- 3304 THEN
            tanh_f := - 1893;
        ELSIF x =- 3303 THEN
            tanh_f := - 1892;
        ELSIF x =- 3302 THEN
            tanh_f := - 1892;
        ELSIF x =- 3301 THEN
            tanh_f := - 1892;
        ELSIF x =- 3300 THEN
            tanh_f := - 1892;
        ELSIF x =- 3299 THEN
            tanh_f := - 1892;
        ELSIF x =- 3298 THEN
            tanh_f := - 1892;
        ELSIF x =- 3297 THEN
            tanh_f := - 1891;
        ELSIF x =- 3296 THEN
            tanh_f := - 1891;
        ELSIF x =- 3295 THEN
            tanh_f := - 1891;
        ELSIF x =- 3294 THEN
            tanh_f := - 1891;
        ELSIF x =- 3293 THEN
            tanh_f := - 1891;
        ELSIF x =- 3292 THEN
            tanh_f := - 1891;
        ELSIF x =- 3291 THEN
            tanh_f := - 1890;
        ELSIF x =- 3290 THEN
            tanh_f := - 1890;
        ELSIF x =- 3289 THEN
            tanh_f := - 1890;
        ELSIF x =- 3288 THEN
            tanh_f := - 1890;
        ELSIF x =- 3287 THEN
            tanh_f := - 1890;
        ELSIF x =- 3286 THEN
            tanh_f := - 1890;
        ELSIF x =- 3285 THEN
            tanh_f := - 1889;
        ELSIF x =- 3284 THEN
            tanh_f := - 1889;
        ELSIF x =- 3283 THEN
            tanh_f := - 1889;
        ELSIF x =- 3282 THEN
            tanh_f := - 1889;
        ELSIF x =- 3281 THEN
            tanh_f := - 1889;
        ELSIF x =- 3280 THEN
            tanh_f := - 1889;
        ELSIF x =- 3279 THEN
            tanh_f := - 1888;
        ELSIF x =- 3278 THEN
            tanh_f := - 1888;
        ELSIF x =- 3277 THEN
            tanh_f := - 1888;
        ELSIF x =- 3276 THEN
            tanh_f := - 1888;
        ELSIF x =- 3275 THEN
            tanh_f := - 1888;
        ELSIF x =- 3274 THEN
            tanh_f := - 1888;
        ELSIF x =- 3273 THEN
            tanh_f := - 1887;
        ELSIF x =- 3272 THEN
            tanh_f := - 1887;
        ELSIF x =- 3271 THEN
            tanh_f := - 1887;
        ELSIF x =- 3270 THEN
            tanh_f := - 1887;
        ELSIF x =- 3269 THEN
            tanh_f := - 1887;
        ELSIF x =- 3268 THEN
            tanh_f := - 1887;
        ELSIF x =- 3267 THEN
            tanh_f := - 1886;
        ELSIF x =- 3266 THEN
            tanh_f := - 1886;
        ELSIF x =- 3265 THEN
            tanh_f := - 1886;
        ELSIF x =- 3264 THEN
            tanh_f := - 1886;
        ELSIF x =- 3263 THEN
            tanh_f := - 1886;
        ELSIF x =- 3262 THEN
            tanh_f := - 1886;
        ELSIF x =- 3261 THEN
            tanh_f := - 1886;
        ELSIF x =- 3260 THEN
            tanh_f := - 1885;
        ELSIF x =- 3259 THEN
            tanh_f := - 1885;
        ELSIF x =- 3258 THEN
            tanh_f := - 1885;
        ELSIF x =- 3257 THEN
            tanh_f := - 1885;
        ELSIF x =- 3256 THEN
            tanh_f := - 1885;
        ELSIF x =- 3255 THEN
            tanh_f := - 1885;
        ELSIF x =- 3254 THEN
            tanh_f := - 1884;
        ELSIF x =- 3253 THEN
            tanh_f := - 1884;
        ELSIF x =- 3252 THEN
            tanh_f := - 1884;
        ELSIF x =- 3251 THEN
            tanh_f := - 1884;
        ELSIF x =- 3250 THEN
            tanh_f := - 1884;
        ELSIF x =- 3249 THEN
            tanh_f := - 1884;
        ELSIF x =- 3248 THEN
            tanh_f := - 1883;
        ELSIF x =- 3247 THEN
            tanh_f := - 1883;
        ELSIF x =- 3246 THEN
            tanh_f := - 1883;
        ELSIF x =- 3245 THEN
            tanh_f := - 1883;
        ELSIF x =- 3244 THEN
            tanh_f := - 1883;
        ELSIF x =- 3243 THEN
            tanh_f := - 1883;
        ELSIF x =- 3242 THEN
            tanh_f := - 1882;
        ELSIF x =- 3241 THEN
            tanh_f := - 1882;
        ELSIF x =- 3240 THEN
            tanh_f := - 1882;
        ELSIF x =- 3239 THEN
            tanh_f := - 1882;
        ELSIF x =- 3238 THEN
            tanh_f := - 1882;
        ELSIF x =- 3237 THEN
            tanh_f := - 1882;
        ELSIF x =- 3236 THEN
            tanh_f := - 1881;
        ELSIF x =- 3235 THEN
            tanh_f := - 1881;
        ELSIF x =- 3234 THEN
            tanh_f := - 1881;
        ELSIF x =- 3233 THEN
            tanh_f := - 1881;
        ELSIF x =- 3232 THEN
            tanh_f := - 1881;
        ELSIF x =- 3231 THEN
            tanh_f := - 1881;
        ELSIF x =- 3230 THEN
            tanh_f := - 1880;
        ELSIF x =- 3229 THEN
            tanh_f := - 1880;
        ELSIF x =- 3228 THEN
            tanh_f := - 1880;
        ELSIF x =- 3227 THEN
            tanh_f := - 1880;
        ELSIF x =- 3226 THEN
            tanh_f := - 1880;
        ELSIF x =- 3225 THEN
            tanh_f := - 1880;
        ELSIF x =- 3224 THEN
            tanh_f := - 1879;
        ELSIF x =- 3223 THEN
            tanh_f := - 1879;
        ELSIF x =- 3222 THEN
            tanh_f := - 1879;
        ELSIF x =- 3221 THEN
            tanh_f := - 1879;
        ELSIF x =- 3220 THEN
            tanh_f := - 1879;
        ELSIF x =- 3219 THEN
            tanh_f := - 1879;
        ELSIF x =- 3218 THEN
            tanh_f := - 1878;
        ELSIF x =- 3217 THEN
            tanh_f := - 1878;
        ELSIF x =- 3216 THEN
            tanh_f := - 1878;
        ELSIF x =- 3215 THEN
            tanh_f := - 1878;
        ELSIF x =- 3214 THEN
            tanh_f := - 1878;
        ELSIF x =- 3213 THEN
            tanh_f := - 1878;
        ELSIF x =- 3212 THEN
            tanh_f := - 1877;
        ELSIF x =- 3211 THEN
            tanh_f := - 1877;
        ELSIF x =- 3210 THEN
            tanh_f := - 1877;
        ELSIF x =- 3209 THEN
            tanh_f := - 1877;
        ELSIF x =- 3208 THEN
            tanh_f := - 1877;
        ELSIF x =- 3207 THEN
            tanh_f := - 1877;
        ELSIF x =- 3206 THEN
            tanh_f := - 1876;
        ELSIF x =- 3205 THEN
            tanh_f := - 1876;
        ELSIF x =- 3204 THEN
            tanh_f := - 1876;
        ELSIF x =- 3203 THEN
            tanh_f := - 1876;
        ELSIF x =- 3202 THEN
            tanh_f := - 1876;
        ELSIF x =- 3201 THEN
            tanh_f := - 1876;
        ELSIF x =- 3200 THEN
            tanh_f := - 1875;
        ELSIF x =- 3199 THEN
            tanh_f := - 1875;
        ELSIF x =- 3198 THEN
            tanh_f := - 1875;
        ELSIF x =- 3197 THEN
            tanh_f := - 1875;
        ELSIF x =- 3196 THEN
            tanh_f := - 1875;
        ELSIF x =- 3195 THEN
            tanh_f := - 1875;
        ELSIF x =- 3194 THEN
            tanh_f := - 1875;
        ELSIF x =- 3193 THEN
            tanh_f := - 1874;
        ELSIF x =- 3192 THEN
            tanh_f := - 1874;
        ELSIF x =- 3191 THEN
            tanh_f := - 1874;
        ELSIF x =- 3190 THEN
            tanh_f := - 1874;
        ELSIF x =- 3189 THEN
            tanh_f := - 1874;
        ELSIF x =- 3188 THEN
            tanh_f := - 1874;
        ELSIF x =- 3187 THEN
            tanh_f := - 1873;
        ELSIF x =- 3186 THEN
            tanh_f := - 1873;
        ELSIF x =- 3185 THEN
            tanh_f := - 1873;
        ELSIF x =- 3184 THEN
            tanh_f := - 1873;
        ELSIF x =- 3183 THEN
            tanh_f := - 1873;
        ELSIF x =- 3182 THEN
            tanh_f := - 1873;
        ELSIF x =- 3181 THEN
            tanh_f := - 1872;
        ELSIF x =- 3180 THEN
            tanh_f := - 1872;
        ELSIF x =- 3179 THEN
            tanh_f := - 1872;
        ELSIF x =- 3178 THEN
            tanh_f := - 1872;
        ELSIF x =- 3177 THEN
            tanh_f := - 1872;
        ELSIF x =- 3176 THEN
            tanh_f := - 1872;
        ELSIF x =- 3175 THEN
            tanh_f := - 1871;
        ELSIF x =- 3174 THEN
            tanh_f := - 1871;
        ELSIF x =- 3173 THEN
            tanh_f := - 1871;
        ELSIF x =- 3172 THEN
            tanh_f := - 1871;
        ELSIF x =- 3171 THEN
            tanh_f := - 1871;
        ELSIF x =- 3170 THEN
            tanh_f := - 1871;
        ELSIF x =- 3169 THEN
            tanh_f := - 1870;
        ELSIF x =- 3168 THEN
            tanh_f := - 1870;
        ELSIF x =- 3167 THEN
            tanh_f := - 1870;
        ELSIF x =- 3166 THEN
            tanh_f := - 1870;
        ELSIF x =- 3165 THEN
            tanh_f := - 1870;
        ELSIF x =- 3164 THEN
            tanh_f := - 1870;
        ELSIF x =- 3163 THEN
            tanh_f := - 1869;
        ELSIF x =- 3162 THEN
            tanh_f := - 1869;
        ELSIF x =- 3161 THEN
            tanh_f := - 1869;
        ELSIF x =- 3160 THEN
            tanh_f := - 1869;
        ELSIF x =- 3159 THEN
            tanh_f := - 1869;
        ELSIF x =- 3158 THEN
            tanh_f := - 1869;
        ELSIF x =- 3157 THEN
            tanh_f := - 1868;
        ELSIF x =- 3156 THEN
            tanh_f := - 1868;
        ELSIF x =- 3155 THEN
            tanh_f := - 1868;
        ELSIF x =- 3154 THEN
            tanh_f := - 1868;
        ELSIF x =- 3153 THEN
            tanh_f := - 1868;
        ELSIF x =- 3152 THEN
            tanh_f := - 1868;
        ELSIF x =- 3151 THEN
            tanh_f := - 1867;
        ELSIF x =- 3150 THEN
            tanh_f := - 1867;
        ELSIF x =- 3149 THEN
            tanh_f := - 1867;
        ELSIF x =- 3148 THEN
            tanh_f := - 1867;
        ELSIF x =- 3147 THEN
            tanh_f := - 1867;
        ELSIF x =- 3146 THEN
            tanh_f := - 1867;
        ELSIF x =- 3145 THEN
            tanh_f := - 1866;
        ELSIF x =- 3144 THEN
            tanh_f := - 1866;
        ELSIF x =- 3143 THEN
            tanh_f := - 1866;
        ELSIF x =- 3142 THEN
            tanh_f := - 1866;
        ELSIF x =- 3141 THEN
            tanh_f := - 1866;
        ELSIF x =- 3140 THEN
            tanh_f := - 1866;
        ELSIF x =- 3139 THEN
            tanh_f := - 1865;
        ELSIF x =- 3138 THEN
            tanh_f := - 1865;
        ELSIF x =- 3137 THEN
            tanh_f := - 1865;
        ELSIF x =- 3136 THEN
            tanh_f := - 1865;
        ELSIF x =- 3135 THEN
            tanh_f := - 1865;
        ELSIF x =- 3134 THEN
            tanh_f := - 1865;
        ELSIF x =- 3133 THEN
            tanh_f := - 1865;
        ELSIF x =- 3132 THEN
            tanh_f := - 1864;
        ELSIF x =- 3131 THEN
            tanh_f := - 1864;
        ELSIF x =- 3130 THEN
            tanh_f := - 1864;
        ELSIF x =- 3129 THEN
            tanh_f := - 1864;
        ELSIF x =- 3128 THEN
            tanh_f := - 1864;
        ELSIF x =- 3127 THEN
            tanh_f := - 1864;
        ELSIF x =- 3126 THEN
            tanh_f := - 1863;
        ELSIF x =- 3125 THEN
            tanh_f := - 1863;
        ELSIF x =- 3124 THEN
            tanh_f := - 1863;
        ELSIF x =- 3123 THEN
            tanh_f := - 1863;
        ELSIF x =- 3122 THEN
            tanh_f := - 1863;
        ELSIF x =- 3121 THEN
            tanh_f := - 1863;
        ELSIF x =- 3120 THEN
            tanh_f := - 1862;
        ELSIF x =- 3119 THEN
            tanh_f := - 1862;
        ELSIF x =- 3118 THEN
            tanh_f := - 1862;
        ELSIF x =- 3117 THEN
            tanh_f := - 1862;
        ELSIF x =- 3116 THEN
            tanh_f := - 1862;
        ELSIF x =- 3115 THEN
            tanh_f := - 1862;
        ELSIF x =- 3114 THEN
            tanh_f := - 1861;
        ELSIF x =- 3113 THEN
            tanh_f := - 1861;
        ELSIF x =- 3112 THEN
            tanh_f := - 1861;
        ELSIF x =- 3111 THEN
            tanh_f := - 1861;
        ELSIF x =- 3110 THEN
            tanh_f := - 1861;
        ELSIF x =- 3109 THEN
            tanh_f := - 1861;
        ELSIF x =- 3108 THEN
            tanh_f := - 1860;
        ELSIF x =- 3107 THEN
            tanh_f := - 1860;
        ELSIF x =- 3106 THEN
            tanh_f := - 1860;
        ELSIF x =- 3105 THEN
            tanh_f := - 1860;
        ELSIF x =- 3104 THEN
            tanh_f := - 1860;
        ELSIF x =- 3103 THEN
            tanh_f := - 1860;
        ELSIF x =- 3102 THEN
            tanh_f := - 1859;
        ELSIF x =- 3101 THEN
            tanh_f := - 1859;
        ELSIF x =- 3100 THEN
            tanh_f := - 1859;
        ELSIF x =- 3099 THEN
            tanh_f := - 1859;
        ELSIF x =- 3098 THEN
            tanh_f := - 1859;
        ELSIF x =- 3097 THEN
            tanh_f := - 1859;
        ELSIF x =- 3096 THEN
            tanh_f := - 1858;
        ELSIF x =- 3095 THEN
            tanh_f := - 1858;
        ELSIF x =- 3094 THEN
            tanh_f := - 1858;
        ELSIF x =- 3093 THEN
            tanh_f := - 1858;
        ELSIF x =- 3092 THEN
            tanh_f := - 1858;
        ELSIF x =- 3091 THEN
            tanh_f := - 1858;
        ELSIF x =- 3090 THEN
            tanh_f := - 1857;
        ELSIF x =- 3089 THEN
            tanh_f := - 1857;
        ELSIF x =- 3088 THEN
            tanh_f := - 1857;
        ELSIF x =- 3087 THEN
            tanh_f := - 1857;
        ELSIF x =- 3086 THEN
            tanh_f := - 1857;
        ELSIF x =- 3085 THEN
            tanh_f := - 1857;
        ELSIF x =- 3084 THEN
            tanh_f := - 1856;
        ELSIF x =- 3083 THEN
            tanh_f := - 1856;
        ELSIF x =- 3082 THEN
            tanh_f := - 1856;
        ELSIF x =- 3081 THEN
            tanh_f := - 1856;
        ELSIF x =- 3080 THEN
            tanh_f := - 1856;
        ELSIF x =- 3079 THEN
            tanh_f := - 1856;
        ELSIF x =- 3078 THEN
            tanh_f := - 1855;
        ELSIF x =- 3077 THEN
            tanh_f := - 1855;
        ELSIF x =- 3076 THEN
            tanh_f := - 1855;
        ELSIF x =- 3075 THEN
            tanh_f := - 1855;
        ELSIF x =- 3074 THEN
            tanh_f := - 1855;
        ELSIF x =- 3073 THEN
            tanh_f := - 1855;
        ELSIF x =- 3072 THEN
            tanh_f := - 1854;
        ELSIF x =- 3071 THEN
            tanh_f := - 1854;
        ELSIF x =- 3070 THEN
            tanh_f := - 1854;
        ELSIF x =- 3069 THEN
            tanh_f := - 1854;
        ELSIF x =- 3068 THEN
            tanh_f := - 1854;
        ELSIF x =- 3067 THEN
            tanh_f := - 1854;
        ELSIF x =- 3066 THEN
            tanh_f := - 1853;
        ELSIF x =- 3065 THEN
            tanh_f := - 1853;
        ELSIF x =- 3064 THEN
            tanh_f := - 1853;
        ELSIF x =- 3063 THEN
            tanh_f := - 1853;
        ELSIF x =- 3062 THEN
            tanh_f := - 1853;
        ELSIF x =- 3061 THEN
            tanh_f := - 1852;
        ELSIF x =- 3060 THEN
            tanh_f := - 1852;
        ELSIF x =- 3059 THEN
            tanh_f := - 1852;
        ELSIF x =- 3058 THEN
            tanh_f := - 1852;
        ELSIF x =- 3057 THEN
            tanh_f := - 1852;
        ELSIF x =- 3056 THEN
            tanh_f := - 1851;
        ELSIF x =- 3055 THEN
            tanh_f := - 1851;
        ELSIF x =- 3054 THEN
            tanh_f := - 1851;
        ELSIF x =- 3053 THEN
            tanh_f := - 1851;
        ELSIF x =- 3052 THEN
            tanh_f := - 1851;
        ELSIF x =- 3051 THEN
            tanh_f := - 1850;
        ELSIF x =- 3050 THEN
            tanh_f := - 1850;
        ELSIF x =- 3049 THEN
            tanh_f := - 1850;
        ELSIF x =- 3048 THEN
            tanh_f := - 1850;
        ELSIF x =- 3047 THEN
            tanh_f := - 1850;
        ELSIF x =- 3046 THEN
            tanh_f := - 1849;
        ELSIF x =- 3045 THEN
            tanh_f := - 1849;
        ELSIF x =- 3044 THEN
            tanh_f := - 1849;
        ELSIF x =- 3043 THEN
            tanh_f := - 1849;
        ELSIF x =- 3042 THEN
            tanh_f := - 1849;
        ELSIF x =- 3041 THEN
            tanh_f := - 1848;
        ELSIF x =- 3040 THEN
            tanh_f := - 1848;
        ELSIF x =- 3039 THEN
            tanh_f := - 1848;
        ELSIF x =- 3038 THEN
            tanh_f := - 1848;
        ELSIF x =- 3037 THEN
            tanh_f := - 1848;
        ELSIF x =- 3036 THEN
            tanh_f := - 1847;
        ELSIF x =- 3035 THEN
            tanh_f := - 1847;
        ELSIF x =- 3034 THEN
            tanh_f := - 1847;
        ELSIF x =- 3033 THEN
            tanh_f := - 1847;
        ELSIF x =- 3032 THEN
            tanh_f := - 1847;
        ELSIF x =- 3031 THEN
            tanh_f := - 1846;
        ELSIF x =- 3030 THEN
            tanh_f := - 1846;
        ELSIF x =- 3029 THEN
            tanh_f := - 1846;
        ELSIF x =- 3028 THEN
            tanh_f := - 1846;
        ELSIF x =- 3027 THEN
            tanh_f := - 1846;
        ELSIF x =- 3026 THEN
            tanh_f := - 1845;
        ELSIF x =- 3025 THEN
            tanh_f := - 1845;
        ELSIF x =- 3024 THEN
            tanh_f := - 1845;
        ELSIF x =- 3023 THEN
            tanh_f := - 1845;
        ELSIF x =- 3022 THEN
            tanh_f := - 1845;
        ELSIF x =- 3021 THEN
            tanh_f := - 1844;
        ELSIF x =- 3020 THEN
            tanh_f := - 1844;
        ELSIF x =- 3019 THEN
            tanh_f := - 1844;
        ELSIF x =- 3018 THEN
            tanh_f := - 1844;
        ELSIF x =- 3017 THEN
            tanh_f := - 1844;
        ELSIF x =- 3016 THEN
            tanh_f := - 1843;
        ELSIF x =- 3015 THEN
            tanh_f := - 1843;
        ELSIF x =- 3014 THEN
            tanh_f := - 1843;
        ELSIF x =- 3013 THEN
            tanh_f := - 1843;
        ELSIF x =- 3012 THEN
            tanh_f := - 1843;
        ELSIF x =- 3011 THEN
            tanh_f := - 1842;
        ELSIF x =- 3010 THEN
            tanh_f := - 1842;
        ELSIF x =- 3009 THEN
            tanh_f := - 1842;
        ELSIF x =- 3008 THEN
            tanh_f := - 1842;
        ELSIF x =- 3007 THEN
            tanh_f := - 1842;
        ELSIF x =- 3006 THEN
            tanh_f := - 1841;
        ELSIF x =- 3005 THEN
            tanh_f := - 1841;
        ELSIF x =- 3004 THEN
            tanh_f := - 1841;
        ELSIF x =- 3003 THEN
            tanh_f := - 1841;
        ELSIF x =- 3002 THEN
            tanh_f := - 1841;
        ELSIF x =- 3001 THEN
            tanh_f := - 1840;
        ELSIF x =- 3000 THEN
            tanh_f := - 1840;
        ELSIF x =- 2999 THEN
            tanh_f := - 1840;
        ELSIF x =- 2998 THEN
            tanh_f := - 1840;
        ELSIF x =- 2997 THEN
            tanh_f := - 1840;
        ELSIF x =- 2996 THEN
            tanh_f := - 1839;
        ELSIF x =- 2995 THEN
            tanh_f := - 1839;
        ELSIF x =- 2994 THEN
            tanh_f := - 1839;
        ELSIF x =- 2993 THEN
            tanh_f := - 1839;
        ELSIF x =- 2992 THEN
            tanh_f := - 1839;
        ELSIF x =- 2991 THEN
            tanh_f := - 1838;
        ELSIF x =- 2990 THEN
            tanh_f := - 1838;
        ELSIF x =- 2989 THEN
            tanh_f := - 1838;
        ELSIF x =- 2988 THEN
            tanh_f := - 1838;
        ELSIF x =- 2987 THEN
            tanh_f := - 1838;
        ELSIF x =- 2986 THEN
            tanh_f := - 1837;
        ELSIF x =- 2985 THEN
            tanh_f := - 1837;
        ELSIF x =- 2984 THEN
            tanh_f := - 1837;
        ELSIF x =- 2983 THEN
            tanh_f := - 1837;
        ELSIF x =- 2982 THEN
            tanh_f := - 1837;
        ELSIF x =- 2981 THEN
            tanh_f := - 1836;
        ELSIF x =- 2980 THEN
            tanh_f := - 1836;
        ELSIF x =- 2979 THEN
            tanh_f := - 1836;
        ELSIF x =- 2978 THEN
            tanh_f := - 1836;
        ELSIF x =- 2977 THEN
            tanh_f := - 1836;
        ELSIF x =- 2976 THEN
            tanh_f := - 1835;
        ELSIF x =- 2975 THEN
            tanh_f := - 1835;
        ELSIF x =- 2974 THEN
            tanh_f := - 1835;
        ELSIF x =- 2973 THEN
            tanh_f := - 1835;
        ELSIF x =- 2972 THEN
            tanh_f := - 1835;
        ELSIF x =- 2971 THEN
            tanh_f := - 1834;
        ELSIF x =- 2970 THEN
            tanh_f := - 1834;
        ELSIF x =- 2969 THEN
            tanh_f := - 1834;
        ELSIF x =- 2968 THEN
            tanh_f := - 1834;
        ELSIF x =- 2967 THEN
            tanh_f := - 1834;
        ELSIF x =- 2966 THEN
            tanh_f := - 1833;
        ELSIF x =- 2965 THEN
            tanh_f := - 1833;
        ELSIF x =- 2964 THEN
            tanh_f := - 1833;
        ELSIF x =- 2963 THEN
            tanh_f := - 1833;
        ELSIF x =- 2962 THEN
            tanh_f := - 1833;
        ELSIF x =- 2961 THEN
            tanh_f := - 1832;
        ELSIF x =- 2960 THEN
            tanh_f := - 1832;
        ELSIF x =- 2959 THEN
            tanh_f := - 1832;
        ELSIF x =- 2958 THEN
            tanh_f := - 1832;
        ELSIF x =- 2957 THEN
            tanh_f := - 1832;
        ELSIF x =- 2956 THEN
            tanh_f := - 1831;
        ELSIF x =- 2955 THEN
            tanh_f := - 1831;
        ELSIF x =- 2954 THEN
            tanh_f := - 1831;
        ELSIF x =- 2953 THEN
            tanh_f := - 1831;
        ELSIF x =- 2952 THEN
            tanh_f := - 1831;
        ELSIF x =- 2951 THEN
            tanh_f := - 1830;
        ELSIF x =- 2950 THEN
            tanh_f := - 1830;
        ELSIF x =- 2949 THEN
            tanh_f := - 1830;
        ELSIF x =- 2948 THEN
            tanh_f := - 1830;
        ELSIF x =- 2947 THEN
            tanh_f := - 1830;
        ELSIF x =- 2946 THEN
            tanh_f := - 1829;
        ELSIF x =- 2945 THEN
            tanh_f := - 1829;
        ELSIF x =- 2944 THEN
            tanh_f := - 1829;
        ELSIF x =- 2943 THEN
            tanh_f := - 1829;
        ELSIF x =- 2942 THEN
            tanh_f := - 1829;
        ELSIF x =- 2941 THEN
            tanh_f := - 1828;
        ELSIF x =- 2940 THEN
            tanh_f := - 1828;
        ELSIF x =- 2939 THEN
            tanh_f := - 1828;
        ELSIF x =- 2938 THEN
            tanh_f := - 1828;
        ELSIF x =- 2937 THEN
            tanh_f := - 1828;
        ELSIF x =- 2936 THEN
            tanh_f := - 1827;
        ELSIF x =- 2935 THEN
            tanh_f := - 1827;
        ELSIF x =- 2934 THEN
            tanh_f := - 1827;
        ELSIF x =- 2933 THEN
            tanh_f := - 1827;
        ELSIF x =- 2932 THEN
            tanh_f := - 1827;
        ELSIF x =- 2931 THEN
            tanh_f := - 1826;
        ELSIF x =- 2930 THEN
            tanh_f := - 1826;
        ELSIF x =- 2929 THEN
            tanh_f := - 1826;
        ELSIF x =- 2928 THEN
            tanh_f := - 1826;
        ELSIF x =- 2927 THEN
            tanh_f := - 1826;
        ELSIF x =- 2926 THEN
            tanh_f := - 1825;
        ELSIF x =- 2925 THEN
            tanh_f := - 1825;
        ELSIF x =- 2924 THEN
            tanh_f := - 1825;
        ELSIF x =- 2923 THEN
            tanh_f := - 1825;
        ELSIF x =- 2922 THEN
            tanh_f := - 1825;
        ELSIF x =- 2921 THEN
            tanh_f := - 1824;
        ELSIF x =- 2920 THEN
            tanh_f := - 1824;
        ELSIF x =- 2919 THEN
            tanh_f := - 1824;
        ELSIF x =- 2918 THEN
            tanh_f := - 1824;
        ELSIF x =- 2917 THEN
            tanh_f := - 1824;
        ELSIF x =- 2916 THEN
            tanh_f := - 1823;
        ELSIF x =- 2915 THEN
            tanh_f := - 1823;
        ELSIF x =- 2914 THEN
            tanh_f := - 1823;
        ELSIF x =- 2913 THEN
            tanh_f := - 1823;
        ELSIF x =- 2912 THEN
            tanh_f := - 1823;
        ELSIF x =- 2911 THEN
            tanh_f := - 1822;
        ELSIF x =- 2910 THEN
            tanh_f := - 1822;
        ELSIF x =- 2909 THEN
            tanh_f := - 1822;
        ELSIF x =- 2908 THEN
            tanh_f := - 1822;
        ELSIF x =- 2907 THEN
            tanh_f := - 1822;
        ELSIF x =- 2906 THEN
            tanh_f := - 1821;
        ELSIF x =- 2905 THEN
            tanh_f := - 1821;
        ELSIF x =- 2904 THEN
            tanh_f := - 1821;
        ELSIF x =- 2903 THEN
            tanh_f := - 1821;
        ELSIF x =- 2902 THEN
            tanh_f := - 1821;
        ELSIF x =- 2901 THEN
            tanh_f := - 1820;
        ELSIF x =- 2900 THEN
            tanh_f := - 1820;
        ELSIF x =- 2899 THEN
            tanh_f := - 1820;
        ELSIF x =- 2898 THEN
            tanh_f := - 1820;
        ELSIF x =- 2897 THEN
            tanh_f := - 1820;
        ELSIF x =- 2896 THEN
            tanh_f := - 1819;
        ELSIF x =- 2895 THEN
            tanh_f := - 1819;
        ELSIF x =- 2894 THEN
            tanh_f := - 1819;
        ELSIF x =- 2893 THEN
            tanh_f := - 1819;
        ELSIF x =- 2892 THEN
            tanh_f := - 1819;
        ELSIF x =- 2891 THEN
            tanh_f := - 1818;
        ELSIF x =- 2890 THEN
            tanh_f := - 1818;
        ELSIF x =- 2889 THEN
            tanh_f := - 1818;
        ELSIF x =- 2888 THEN
            tanh_f := - 1818;
        ELSIF x =- 2887 THEN
            tanh_f := - 1818;
        ELSIF x =- 2886 THEN
            tanh_f := - 1817;
        ELSIF x =- 2885 THEN
            tanh_f := - 1817;
        ELSIF x =- 2884 THEN
            tanh_f := - 1817;
        ELSIF x =- 2883 THEN
            tanh_f := - 1817;
        ELSIF x =- 2882 THEN
            tanh_f := - 1817;
        ELSIF x =- 2881 THEN
            tanh_f := - 1816;
        ELSIF x =- 2880 THEN
            tanh_f := - 1816;
        ELSIF x =- 2879 THEN
            tanh_f := - 1816;
        ELSIF x =- 2878 THEN
            tanh_f := - 1816;
        ELSIF x =- 2877 THEN
            tanh_f := - 1816;
        ELSIF x =- 2876 THEN
            tanh_f := - 1815;
        ELSIF x =- 2875 THEN
            tanh_f := - 1815;
        ELSIF x =- 2874 THEN
            tanh_f := - 1815;
        ELSIF x =- 2873 THEN
            tanh_f := - 1815;
        ELSIF x =- 2872 THEN
            tanh_f := - 1815;
        ELSIF x =- 2871 THEN
            tanh_f := - 1814;
        ELSIF x =- 2870 THEN
            tanh_f := - 1814;
        ELSIF x =- 2869 THEN
            tanh_f := - 1814;
        ELSIF x =- 2868 THEN
            tanh_f := - 1814;
        ELSIF x =- 2867 THEN
            tanh_f := - 1814;
        ELSIF x =- 2866 THEN
            tanh_f := - 1813;
        ELSIF x =- 2865 THEN
            tanh_f := - 1813;
        ELSIF x =- 2864 THEN
            tanh_f := - 1813;
        ELSIF x =- 2863 THEN
            tanh_f := - 1813;
        ELSIF x =- 2862 THEN
            tanh_f := - 1813;
        ELSIF x =- 2861 THEN
            tanh_f := - 1812;
        ELSIF x =- 2860 THEN
            tanh_f := - 1812;
        ELSIF x =- 2859 THEN
            tanh_f := - 1812;
        ELSIF x =- 2858 THEN
            tanh_f := - 1812;
        ELSIF x =- 2857 THEN
            tanh_f := - 1812;
        ELSIF x =- 2856 THEN
            tanh_f := - 1811;
        ELSIF x =- 2855 THEN
            tanh_f := - 1811;
        ELSIF x =- 2854 THEN
            tanh_f := - 1811;
        ELSIF x =- 2853 THEN
            tanh_f := - 1811;
        ELSIF x =- 2852 THEN
            tanh_f := - 1811;
        ELSIF x =- 2851 THEN
            tanh_f := - 1810;
        ELSIF x =- 2850 THEN
            tanh_f := - 1810;
        ELSIF x =- 2849 THEN
            tanh_f := - 1810;
        ELSIF x =- 2848 THEN
            tanh_f := - 1810;
        ELSIF x =- 2847 THEN
            tanh_f := - 1810;
        ELSIF x =- 2846 THEN
            tanh_f := - 1809;
        ELSIF x =- 2845 THEN
            tanh_f := - 1809;
        ELSIF x =- 2844 THEN
            tanh_f := - 1809;
        ELSIF x =- 2843 THEN
            tanh_f := - 1809;
        ELSIF x =- 2842 THEN
            tanh_f := - 1809;
        ELSIF x =- 2841 THEN
            tanh_f := - 1808;
        ELSIF x =- 2840 THEN
            tanh_f := - 1808;
        ELSIF x =- 2839 THEN
            tanh_f := - 1808;
        ELSIF x =- 2838 THEN
            tanh_f := - 1808;
        ELSIF x =- 2837 THEN
            tanh_f := - 1808;
        ELSIF x =- 2836 THEN
            tanh_f := - 1807;
        ELSIF x =- 2835 THEN
            tanh_f := - 1807;
        ELSIF x =- 2834 THEN
            tanh_f := - 1807;
        ELSIF x =- 2833 THEN
            tanh_f := - 1807;
        ELSIF x =- 2832 THEN
            tanh_f := - 1807;
        ELSIF x =- 2831 THEN
            tanh_f := - 1806;
        ELSIF x =- 2830 THEN
            tanh_f := - 1806;
        ELSIF x =- 2829 THEN
            tanh_f := - 1806;
        ELSIF x =- 2828 THEN
            tanh_f := - 1806;
        ELSIF x =- 2827 THEN
            tanh_f := - 1806;
        ELSIF x =- 2826 THEN
            tanh_f := - 1805;
        ELSIF x =- 2825 THEN
            tanh_f := - 1805;
        ELSIF x =- 2824 THEN
            tanh_f := - 1805;
        ELSIF x =- 2823 THEN
            tanh_f := - 1805;
        ELSIF x =- 2822 THEN
            tanh_f := - 1805;
        ELSIF x =- 2821 THEN
            tanh_f := - 1804;
        ELSIF x =- 2820 THEN
            tanh_f := - 1804;
        ELSIF x =- 2819 THEN
            tanh_f := - 1804;
        ELSIF x =- 2818 THEN
            tanh_f := - 1804;
        ELSIF x =- 2817 THEN
            tanh_f := - 1804;
        ELSIF x =- 2816 THEN
            tanh_f := - 1803;
        ELSIF x =- 2815 THEN
            tanh_f := - 1803;
        ELSIF x =- 2814 THEN
            tanh_f := - 1803;
        ELSIF x =- 2813 THEN
            tanh_f := - 1802;
        ELSIF x =- 2812 THEN
            tanh_f := - 1802;
        ELSIF x =- 2811 THEN
            tanh_f := - 1802;
        ELSIF x =- 2810 THEN
            tanh_f := - 1802;
        ELSIF x =- 2809 THEN
            tanh_f := - 1801;
        ELSIF x =- 2808 THEN
            tanh_f := - 1801;
        ELSIF x =- 2807 THEN
            tanh_f := - 1801;
        ELSIF x =- 2806 THEN
            tanh_f := - 1801;
        ELSIF x =- 2805 THEN
            tanh_f := - 1800;
        ELSIF x =- 2804 THEN
            tanh_f := - 1800;
        ELSIF x =- 2803 THEN
            tanh_f := - 1800;
        ELSIF x =- 2802 THEN
            tanh_f := - 1800;
        ELSIF x =- 2801 THEN
            tanh_f := - 1799;
        ELSIF x =- 2800 THEN
            tanh_f := - 1799;
        ELSIF x =- 2799 THEN
            tanh_f := - 1799;
        ELSIF x =- 2798 THEN
            tanh_f := - 1799;
        ELSIF x =- 2797 THEN
            tanh_f := - 1798;
        ELSIF x =- 2796 THEN
            tanh_f := - 1798;
        ELSIF x =- 2795 THEN
            tanh_f := - 1798;
        ELSIF x =- 2794 THEN
            tanh_f := - 1798;
        ELSIF x =- 2793 THEN
            tanh_f := - 1797;
        ELSIF x =- 2792 THEN
            tanh_f := - 1797;
        ELSIF x =- 2791 THEN
            tanh_f := - 1797;
        ELSIF x =- 2790 THEN
            tanh_f := - 1797;
        ELSIF x =- 2789 THEN
            tanh_f := - 1796;
        ELSIF x =- 2788 THEN
            tanh_f := - 1796;
        ELSIF x =- 2787 THEN
            tanh_f := - 1796;
        ELSIF x =- 2786 THEN
            tanh_f := - 1796;
        ELSIF x =- 2785 THEN
            tanh_f := - 1795;
        ELSIF x =- 2784 THEN
            tanh_f := - 1795;
        ELSIF x =- 2783 THEN
            tanh_f := - 1795;
        ELSIF x =- 2782 THEN
            tanh_f := - 1795;
        ELSIF x =- 2781 THEN
            tanh_f := - 1794;
        ELSIF x =- 2780 THEN
            tanh_f := - 1794;
        ELSIF x =- 2779 THEN
            tanh_f := - 1794;
        ELSIF x =- 2778 THEN
            tanh_f := - 1794;
        ELSIF x =- 2777 THEN
            tanh_f := - 1793;
        ELSIF x =- 2776 THEN
            tanh_f := - 1793;
        ELSIF x =- 2775 THEN
            tanh_f := - 1793;
        ELSIF x =- 2774 THEN
            tanh_f := - 1793;
        ELSIF x =- 2773 THEN
            tanh_f := - 1792;
        ELSIF x =- 2772 THEN
            tanh_f := - 1792;
        ELSIF x =- 2771 THEN
            tanh_f := - 1792;
        ELSIF x =- 2770 THEN
            tanh_f := - 1792;
        ELSIF x =- 2769 THEN
            tanh_f := - 1791;
        ELSIF x =- 2768 THEN
            tanh_f := - 1791;
        ELSIF x =- 2767 THEN
            tanh_f := - 1791;
        ELSIF x =- 2766 THEN
            tanh_f := - 1791;
        ELSIF x =- 2765 THEN
            tanh_f := - 1790;
        ELSIF x =- 2764 THEN
            tanh_f := - 1790;
        ELSIF x =- 2763 THEN
            tanh_f := - 1790;
        ELSIF x =- 2762 THEN
            tanh_f := - 1790;
        ELSIF x =- 2761 THEN
            tanh_f := - 1789;
        ELSIF x =- 2760 THEN
            tanh_f := - 1789;
        ELSIF x =- 2759 THEN
            tanh_f := - 1789;
        ELSIF x =- 2758 THEN
            tanh_f := - 1789;
        ELSIF x =- 2757 THEN
            tanh_f := - 1788;
        ELSIF x =- 2756 THEN
            tanh_f := - 1788;
        ELSIF x =- 2755 THEN
            tanh_f := - 1788;
        ELSIF x =- 2754 THEN
            tanh_f := - 1788;
        ELSIF x =- 2753 THEN
            tanh_f := - 1787;
        ELSIF x =- 2752 THEN
            tanh_f := - 1787;
        ELSIF x =- 2751 THEN
            tanh_f := - 1787;
        ELSIF x =- 2750 THEN
            tanh_f := - 1787;
        ELSIF x =- 2749 THEN
            tanh_f := - 1786;
        ELSIF x =- 2748 THEN
            tanh_f := - 1786;
        ELSIF x =- 2747 THEN
            tanh_f := - 1786;
        ELSIF x =- 2746 THEN
            tanh_f := - 1786;
        ELSIF x =- 2745 THEN
            tanh_f := - 1785;
        ELSIF x =- 2744 THEN
            tanh_f := - 1785;
        ELSIF x =- 2743 THEN
            tanh_f := - 1785;
        ELSIF x =- 2742 THEN
            tanh_f := - 1785;
        ELSIF x =- 2741 THEN
            tanh_f := - 1784;
        ELSIF x =- 2740 THEN
            tanh_f := - 1784;
        ELSIF x =- 2739 THEN
            tanh_f := - 1784;
        ELSIF x =- 2738 THEN
            tanh_f := - 1784;
        ELSIF x =- 2737 THEN
            tanh_f := - 1783;
        ELSIF x =- 2736 THEN
            tanh_f := - 1783;
        ELSIF x =- 2735 THEN
            tanh_f := - 1783;
        ELSIF x =- 2734 THEN
            tanh_f := - 1783;
        ELSIF x =- 2733 THEN
            tanh_f := - 1782;
        ELSIF x =- 2732 THEN
            tanh_f := - 1782;
        ELSIF x =- 2731 THEN
            tanh_f := - 1782;
        ELSIF x =- 2730 THEN
            tanh_f := - 1782;
        ELSIF x =- 2729 THEN
            tanh_f := - 1781;
        ELSIF x =- 2728 THEN
            tanh_f := - 1781;
        ELSIF x =- 2727 THEN
            tanh_f := - 1781;
        ELSIF x =- 2726 THEN
            tanh_f := - 1781;
        ELSIF x =- 2725 THEN
            tanh_f := - 1780;
        ELSIF x =- 2724 THEN
            tanh_f := - 1780;
        ELSIF x =- 2723 THEN
            tanh_f := - 1780;
        ELSIF x =- 2722 THEN
            tanh_f := - 1780;
        ELSIF x =- 2721 THEN
            tanh_f := - 1779;
        ELSIF x =- 2720 THEN
            tanh_f := - 1779;
        ELSIF x =- 2719 THEN
            tanh_f := - 1779;
        ELSIF x =- 2718 THEN
            tanh_f := - 1779;
        ELSIF x =- 2717 THEN
            tanh_f := - 1778;
        ELSIF x =- 2716 THEN
            tanh_f := - 1778;
        ELSIF x =- 2715 THEN
            tanh_f := - 1778;
        ELSIF x =- 2714 THEN
            tanh_f := - 1778;
        ELSIF x =- 2713 THEN
            tanh_f := - 1777;
        ELSIF x =- 2712 THEN
            tanh_f := - 1777;
        ELSIF x =- 2711 THEN
            tanh_f := - 1777;
        ELSIF x =- 2710 THEN
            tanh_f := - 1777;
        ELSIF x =- 2709 THEN
            tanh_f := - 1776;
        ELSIF x =- 2708 THEN
            tanh_f := - 1776;
        ELSIF x =- 2707 THEN
            tanh_f := - 1776;
        ELSIF x =- 2706 THEN
            tanh_f := - 1776;
        ELSIF x =- 2705 THEN
            tanh_f := - 1775;
        ELSIF x =- 2704 THEN
            tanh_f := - 1775;
        ELSIF x =- 2703 THEN
            tanh_f := - 1775;
        ELSIF x =- 2702 THEN
            tanh_f := - 1775;
        ELSIF x =- 2701 THEN
            tanh_f := - 1774;
        ELSIF x =- 2700 THEN
            tanh_f := - 1774;
        ELSIF x =- 2699 THEN
            tanh_f := - 1774;
        ELSIF x =- 2698 THEN
            tanh_f := - 1774;
        ELSIF x =- 2697 THEN
            tanh_f := - 1773;
        ELSIF x =- 2696 THEN
            tanh_f := - 1773;
        ELSIF x =- 2695 THEN
            tanh_f := - 1773;
        ELSIF x =- 2694 THEN
            tanh_f := - 1773;
        ELSIF x =- 2693 THEN
            tanh_f := - 1772;
        ELSIF x =- 2692 THEN
            tanh_f := - 1772;
        ELSIF x =- 2691 THEN
            tanh_f := - 1772;
        ELSIF x =- 2690 THEN
            tanh_f := - 1772;
        ELSIF x =- 2689 THEN
            tanh_f := - 1771;
        ELSIF x =- 2688 THEN
            tanh_f := - 1771;
        ELSIF x =- 2687 THEN
            tanh_f := - 1771;
        ELSIF x =- 2686 THEN
            tanh_f := - 1771;
        ELSIF x =- 2685 THEN
            tanh_f := - 1771;
        ELSIF x =- 2684 THEN
            tanh_f := - 1770;
        ELSIF x =- 2683 THEN
            tanh_f := - 1770;
        ELSIF x =- 2682 THEN
            tanh_f := - 1770;
        ELSIF x =- 2681 THEN
            tanh_f := - 1770;
        ELSIF x =- 2680 THEN
            tanh_f := - 1769;
        ELSIF x =- 2679 THEN
            tanh_f := - 1769;
        ELSIF x =- 2678 THEN
            tanh_f := - 1769;
        ELSIF x =- 2677 THEN
            tanh_f := - 1769;
        ELSIF x =- 2676 THEN
            tanh_f := - 1768;
        ELSIF x =- 2675 THEN
            tanh_f := - 1768;
        ELSIF x =- 2674 THEN
            tanh_f := - 1768;
        ELSIF x =- 2673 THEN
            tanh_f := - 1768;
        ELSIF x =- 2672 THEN
            tanh_f := - 1767;
        ELSIF x =- 2671 THEN
            tanh_f := - 1767;
        ELSIF x =- 2670 THEN
            tanh_f := - 1767;
        ELSIF x =- 2669 THEN
            tanh_f := - 1767;
        ELSIF x =- 2668 THEN
            tanh_f := - 1766;
        ELSIF x =- 2667 THEN
            tanh_f := - 1766;
        ELSIF x =- 2666 THEN
            tanh_f := - 1766;
        ELSIF x =- 2665 THEN
            tanh_f := - 1766;
        ELSIF x =- 2664 THEN
            tanh_f := - 1765;
        ELSIF x =- 2663 THEN
            tanh_f := - 1765;
        ELSIF x =- 2662 THEN
            tanh_f := - 1765;
        ELSIF x =- 2661 THEN
            tanh_f := - 1765;
        ELSIF x =- 2660 THEN
            tanh_f := - 1764;
        ELSIF x =- 2659 THEN
            tanh_f := - 1764;
        ELSIF x =- 2658 THEN
            tanh_f := - 1764;
        ELSIF x =- 2657 THEN
            tanh_f := - 1764;
        ELSIF x =- 2656 THEN
            tanh_f := - 1763;
        ELSIF x =- 2655 THEN
            tanh_f := - 1763;
        ELSIF x =- 2654 THEN
            tanh_f := - 1763;
        ELSIF x =- 2653 THEN
            tanh_f := - 1763;
        ELSIF x =- 2652 THEN
            tanh_f := - 1762;
        ELSIF x =- 2651 THEN
            tanh_f := - 1762;
        ELSIF x =- 2650 THEN
            tanh_f := - 1762;
        ELSIF x =- 2649 THEN
            tanh_f := - 1762;
        ELSIF x =- 2648 THEN
            tanh_f := - 1761;
        ELSIF x =- 2647 THEN
            tanh_f := - 1761;
        ELSIF x =- 2646 THEN
            tanh_f := - 1761;
        ELSIF x =- 2645 THEN
            tanh_f := - 1761;
        ELSIF x =- 2644 THEN
            tanh_f := - 1760;
        ELSIF x =- 2643 THEN
            tanh_f := - 1760;
        ELSIF x =- 2642 THEN
            tanh_f := - 1760;
        ELSIF x =- 2641 THEN
            tanh_f := - 1760;
        ELSIF x =- 2640 THEN
            tanh_f := - 1759;
        ELSIF x =- 2639 THEN
            tanh_f := - 1759;
        ELSIF x =- 2638 THEN
            tanh_f := - 1759;
        ELSIF x =- 2637 THEN
            tanh_f := - 1759;
        ELSIF x =- 2636 THEN
            tanh_f := - 1758;
        ELSIF x =- 2635 THEN
            tanh_f := - 1758;
        ELSIF x =- 2634 THEN
            tanh_f := - 1758;
        ELSIF x =- 2633 THEN
            tanh_f := - 1758;
        ELSIF x =- 2632 THEN
            tanh_f := - 1757;
        ELSIF x =- 2631 THEN
            tanh_f := - 1757;
        ELSIF x =- 2630 THEN
            tanh_f := - 1757;
        ELSIF x =- 2629 THEN
            tanh_f := - 1757;
        ELSIF x =- 2628 THEN
            tanh_f := - 1756;
        ELSIF x =- 2627 THEN
            tanh_f := - 1756;
        ELSIF x =- 2626 THEN
            tanh_f := - 1756;
        ELSIF x =- 2625 THEN
            tanh_f := - 1756;
        ELSIF x =- 2624 THEN
            tanh_f := - 1755;
        ELSIF x =- 2623 THEN
            tanh_f := - 1755;
        ELSIF x =- 2622 THEN
            tanh_f := - 1755;
        ELSIF x =- 2621 THEN
            tanh_f := - 1755;
        ELSIF x =- 2620 THEN
            tanh_f := - 1754;
        ELSIF x =- 2619 THEN
            tanh_f := - 1754;
        ELSIF x =- 2618 THEN
            tanh_f := - 1754;
        ELSIF x =- 2617 THEN
            tanh_f := - 1754;
        ELSIF x =- 2616 THEN
            tanh_f := - 1753;
        ELSIF x =- 2615 THEN
            tanh_f := - 1753;
        ELSIF x =- 2614 THEN
            tanh_f := - 1753;
        ELSIF x =- 2613 THEN
            tanh_f := - 1753;
        ELSIF x =- 2612 THEN
            tanh_f := - 1752;
        ELSIF x =- 2611 THEN
            tanh_f := - 1752;
        ELSIF x =- 2610 THEN
            tanh_f := - 1752;
        ELSIF x =- 2609 THEN
            tanh_f := - 1752;
        ELSIF x =- 2608 THEN
            tanh_f := - 1751;
        ELSIF x =- 2607 THEN
            tanh_f := - 1751;
        ELSIF x =- 2606 THEN
            tanh_f := - 1751;
        ELSIF x =- 2605 THEN
            tanh_f := - 1751;
        ELSIF x =- 2604 THEN
            tanh_f := - 1750;
        ELSIF x =- 2603 THEN
            tanh_f := - 1750;
        ELSIF x =- 2602 THEN
            tanh_f := - 1750;
        ELSIF x =- 2601 THEN
            tanh_f := - 1750;
        ELSIF x =- 2600 THEN
            tanh_f := - 1749;
        ELSIF x =- 2599 THEN
            tanh_f := - 1749;
        ELSIF x =- 2598 THEN
            tanh_f := - 1749;
        ELSIF x =- 2597 THEN
            tanh_f := - 1749;
        ELSIF x =- 2596 THEN
            tanh_f := - 1748;
        ELSIF x =- 2595 THEN
            tanh_f := - 1748;
        ELSIF x =- 2594 THEN
            tanh_f := - 1748;
        ELSIF x =- 2593 THEN
            tanh_f := - 1748;
        ELSIF x =- 2592 THEN
            tanh_f := - 1747;
        ELSIF x =- 2591 THEN
            tanh_f := - 1747;
        ELSIF x =- 2590 THEN
            tanh_f := - 1747;
        ELSIF x =- 2589 THEN
            tanh_f := - 1747;
        ELSIF x =- 2588 THEN
            tanh_f := - 1746;
        ELSIF x =- 2587 THEN
            tanh_f := - 1746;
        ELSIF x =- 2586 THEN
            tanh_f := - 1746;
        ELSIF x =- 2585 THEN
            tanh_f := - 1746;
        ELSIF x =- 2584 THEN
            tanh_f := - 1745;
        ELSIF x =- 2583 THEN
            tanh_f := - 1745;
        ELSIF x =- 2582 THEN
            tanh_f := - 1745;
        ELSIF x =- 2581 THEN
            tanh_f := - 1745;
        ELSIF x =- 2580 THEN
            tanh_f := - 1744;
        ELSIF x =- 2579 THEN
            tanh_f := - 1744;
        ELSIF x =- 2578 THEN
            tanh_f := - 1744;
        ELSIF x =- 2577 THEN
            tanh_f := - 1744;
        ELSIF x =- 2576 THEN
            tanh_f := - 1743;
        ELSIF x =- 2575 THEN
            tanh_f := - 1743;
        ELSIF x =- 2574 THEN
            tanh_f := - 1743;
        ELSIF x =- 2573 THEN
            tanh_f := - 1743;
        ELSIF x =- 2572 THEN
            tanh_f := - 1742;
        ELSIF x =- 2571 THEN
            tanh_f := - 1742;
        ELSIF x =- 2570 THEN
            tanh_f := - 1742;
        ELSIF x =- 2569 THEN
            tanh_f := - 1742;
        ELSIF x =- 2568 THEN
            tanh_f := - 1741;
        ELSIF x =- 2567 THEN
            tanh_f := - 1741;
        ELSIF x =- 2566 THEN
            tanh_f := - 1741;
        ELSIF x =- 2565 THEN
            tanh_f := - 1741;
        ELSIF x =- 2564 THEN
            tanh_f := - 1740;
        ELSIF x =- 2563 THEN
            tanh_f := - 1740;
        ELSIF x =- 2562 THEN
            tanh_f := - 1740;
        ELSIF x =- 2561 THEN
            tanh_f := - 1740;
        ELSIF x =- 2560 THEN
            tanh_f := - 1739;
        ELSIF x =- 2559 THEN
            tanh_f := - 1739;
        ELSIF x =- 2558 THEN
            tanh_f := - 1739;
        ELSIF x =- 2557 THEN
            tanh_f := - 1739;
        ELSIF x =- 2556 THEN
            tanh_f := - 1738;
        ELSIF x =- 2555 THEN
            tanh_f := - 1738;
        ELSIF x =- 2554 THEN
            tanh_f := - 1738;
        ELSIF x =- 2553 THEN
            tanh_f := - 1737;
        ELSIF x =- 2552 THEN
            tanh_f := - 1737;
        ELSIF x =- 2551 THEN
            tanh_f := - 1737;
        ELSIF x =- 2550 THEN
            tanh_f := - 1736;
        ELSIF x =- 2549 THEN
            tanh_f := - 1736;
        ELSIF x =- 2548 THEN
            tanh_f := - 1736;
        ELSIF x =- 2547 THEN
            tanh_f := - 1735;
        ELSIF x =- 2546 THEN
            tanh_f := - 1735;
        ELSIF x =- 2545 THEN
            tanh_f := - 1735;
        ELSIF x =- 2544 THEN
            tanh_f := - 1734;
        ELSIF x =- 2543 THEN
            tanh_f := - 1734;
        ELSIF x =- 2542 THEN
            tanh_f := - 1734;
        ELSIF x =- 2541 THEN
            tanh_f := - 1734;
        ELSIF x =- 2540 THEN
            tanh_f := - 1733;
        ELSIF x =- 2539 THEN
            tanh_f := - 1733;
        ELSIF x =- 2538 THEN
            tanh_f := - 1733;
        ELSIF x =- 2537 THEN
            tanh_f := - 1732;
        ELSIF x =- 2536 THEN
            tanh_f := - 1732;
        ELSIF x =- 2535 THEN
            tanh_f := - 1732;
        ELSIF x =- 2534 THEN
            tanh_f := - 1731;
        ELSIF x =- 2533 THEN
            tanh_f := - 1731;
        ELSIF x =- 2532 THEN
            tanh_f := - 1731;
        ELSIF x =- 2531 THEN
            tanh_f := - 1730;
        ELSIF x =- 2530 THEN
            tanh_f := - 1730;
        ELSIF x =- 2529 THEN
            tanh_f := - 1730;
        ELSIF x =- 2528 THEN
            tanh_f := - 1729;
        ELSIF x =- 2527 THEN
            tanh_f := - 1729;
        ELSIF x =- 2526 THEN
            tanh_f := - 1729;
        ELSIF x =- 2525 THEN
            tanh_f := - 1728;
        ELSIF x =- 2524 THEN
            tanh_f := - 1728;
        ELSIF x =- 2523 THEN
            tanh_f := - 1728;
        ELSIF x =- 2522 THEN
            tanh_f := - 1728;
        ELSIF x =- 2521 THEN
            tanh_f := - 1727;
        ELSIF x =- 2520 THEN
            tanh_f := - 1727;
        ELSIF x =- 2519 THEN
            tanh_f := - 1727;
        ELSIF x =- 2518 THEN
            tanh_f := - 1726;
        ELSIF x =- 2517 THEN
            tanh_f := - 1726;
        ELSIF x =- 2516 THEN
            tanh_f := - 1726;
        ELSIF x =- 2515 THEN
            tanh_f := - 1725;
        ELSIF x =- 2514 THEN
            tanh_f := - 1725;
        ELSIF x =- 2513 THEN
            tanh_f := - 1725;
        ELSIF x =- 2512 THEN
            tanh_f := - 1724;
        ELSIF x =- 2511 THEN
            tanh_f := - 1724;
        ELSIF x =- 2510 THEN
            tanh_f := - 1724;
        ELSIF x =- 2509 THEN
            tanh_f := - 1723;
        ELSIF x =- 2508 THEN
            tanh_f := - 1723;
        ELSIF x =- 2507 THEN
            tanh_f := - 1723;
        ELSIF x =- 2506 THEN
            tanh_f := - 1723;
        ELSIF x =- 2505 THEN
            tanh_f := - 1722;
        ELSIF x =- 2504 THEN
            tanh_f := - 1722;
        ELSIF x =- 2503 THEN
            tanh_f := - 1722;
        ELSIF x =- 2502 THEN
            tanh_f := - 1721;
        ELSIF x =- 2501 THEN
            tanh_f := - 1721;
        ELSIF x =- 2500 THEN
            tanh_f := - 1721;
        ELSIF x =- 2499 THEN
            tanh_f := - 1720;
        ELSIF x =- 2498 THEN
            tanh_f := - 1720;
        ELSIF x =- 2497 THEN
            tanh_f := - 1720;
        ELSIF x =- 2496 THEN
            tanh_f := - 1719;
        ELSIF x =- 2495 THEN
            tanh_f := - 1719;
        ELSIF x =- 2494 THEN
            tanh_f := - 1719;
        ELSIF x =- 2493 THEN
            tanh_f := - 1718;
        ELSIF x =- 2492 THEN
            tanh_f := - 1718;
        ELSIF x =- 2491 THEN
            tanh_f := - 1718;
        ELSIF x =- 2490 THEN
            tanh_f := - 1717;
        ELSIF x =- 2489 THEN
            tanh_f := - 1717;
        ELSIF x =- 2488 THEN
            tanh_f := - 1717;
        ELSIF x =- 2487 THEN
            tanh_f := - 1717;
        ELSIF x =- 2486 THEN
            tanh_f := - 1716;
        ELSIF x =- 2485 THEN
            tanh_f := - 1716;
        ELSIF x =- 2484 THEN
            tanh_f := - 1716;
        ELSIF x =- 2483 THEN
            tanh_f := - 1715;
        ELSIF x =- 2482 THEN
            tanh_f := - 1715;
        ELSIF x =- 2481 THEN
            tanh_f := - 1715;
        ELSIF x =- 2480 THEN
            tanh_f := - 1714;
        ELSIF x =- 2479 THEN
            tanh_f := - 1714;
        ELSIF x =- 2478 THEN
            tanh_f := - 1714;
        ELSIF x =- 2477 THEN
            tanh_f := - 1713;
        ELSIF x =- 2476 THEN
            tanh_f := - 1713;
        ELSIF x =- 2475 THEN
            tanh_f := - 1713;
        ELSIF x =- 2474 THEN
            tanh_f := - 1712;
        ELSIF x =- 2473 THEN
            tanh_f := - 1712;
        ELSIF x =- 2472 THEN
            tanh_f := - 1712;
        ELSIF x =- 2471 THEN
            tanh_f := - 1712;
        ELSIF x =- 2470 THEN
            tanh_f := - 1711;
        ELSIF x =- 2469 THEN
            tanh_f := - 1711;
        ELSIF x =- 2468 THEN
            tanh_f := - 1711;
        ELSIF x =- 2467 THEN
            tanh_f := - 1710;
        ELSIF x =- 2466 THEN
            tanh_f := - 1710;
        ELSIF x =- 2465 THEN
            tanh_f := - 1710;
        ELSIF x =- 2464 THEN
            tanh_f := - 1709;
        ELSIF x =- 2463 THEN
            tanh_f := - 1709;
        ELSIF x =- 2462 THEN
            tanh_f := - 1709;
        ELSIF x =- 2461 THEN
            tanh_f := - 1708;
        ELSIF x =- 2460 THEN
            tanh_f := - 1708;
        ELSIF x =- 2459 THEN
            tanh_f := - 1708;
        ELSIF x =- 2458 THEN
            tanh_f := - 1707;
        ELSIF x =- 2457 THEN
            tanh_f := - 1707;
        ELSIF x =- 2456 THEN
            tanh_f := - 1707;
        ELSIF x =- 2455 THEN
            tanh_f := - 1706;
        ELSIF x =- 2454 THEN
            tanh_f := - 1706;
        ELSIF x =- 2453 THEN
            tanh_f := - 1706;
        ELSIF x =- 2452 THEN
            tanh_f := - 1706;
        ELSIF x =- 2451 THEN
            tanh_f := - 1705;
        ELSIF x =- 2450 THEN
            tanh_f := - 1705;
        ELSIF x =- 2449 THEN
            tanh_f := - 1705;
        ELSIF x =- 2448 THEN
            tanh_f := - 1704;
        ELSIF x =- 2447 THEN
            tanh_f := - 1704;
        ELSIF x =- 2446 THEN
            tanh_f := - 1704;
        ELSIF x =- 2445 THEN
            tanh_f := - 1703;
        ELSIF x =- 2444 THEN
            tanh_f := - 1703;
        ELSIF x =- 2443 THEN
            tanh_f := - 1703;
        ELSIF x =- 2442 THEN
            tanh_f := - 1702;
        ELSIF x =- 2441 THEN
            tanh_f := - 1702;
        ELSIF x =- 2440 THEN
            tanh_f := - 1702;
        ELSIF x =- 2439 THEN
            tanh_f := - 1701;
        ELSIF x =- 2438 THEN
            tanh_f := - 1701;
        ELSIF x =- 2437 THEN
            tanh_f := - 1701;
        ELSIF x =- 2436 THEN
            tanh_f := - 1701;
        ELSIF x =- 2435 THEN
            tanh_f := - 1700;
        ELSIF x =- 2434 THEN
            tanh_f := - 1700;
        ELSIF x =- 2433 THEN
            tanh_f := - 1700;
        ELSIF x =- 2432 THEN
            tanh_f := - 1699;
        ELSIF x =- 2431 THEN
            tanh_f := - 1699;
        ELSIF x =- 2430 THEN
            tanh_f := - 1699;
        ELSIF x =- 2429 THEN
            tanh_f := - 1698;
        ELSIF x =- 2428 THEN
            tanh_f := - 1698;
        ELSIF x =- 2427 THEN
            tanh_f := - 1698;
        ELSIF x =- 2426 THEN
            tanh_f := - 1697;
        ELSIF x =- 2425 THEN
            tanh_f := - 1697;
        ELSIF x =- 2424 THEN
            tanh_f := - 1697;
        ELSIF x =- 2423 THEN
            tanh_f := - 1696;
        ELSIF x =- 2422 THEN
            tanh_f := - 1696;
        ELSIF x =- 2421 THEN
            tanh_f := - 1696;
        ELSIF x =- 2420 THEN
            tanh_f := - 1695;
        ELSIF x =- 2419 THEN
            tanh_f := - 1695;
        ELSIF x =- 2418 THEN
            tanh_f := - 1695;
        ELSIF x =- 2417 THEN
            tanh_f := - 1695;
        ELSIF x =- 2416 THEN
            tanh_f := - 1694;
        ELSIF x =- 2415 THEN
            tanh_f := - 1694;
        ELSIF x =- 2414 THEN
            tanh_f := - 1694;
        ELSIF x =- 2413 THEN
            tanh_f := - 1693;
        ELSIF x =- 2412 THEN
            tanh_f := - 1693;
        ELSIF x =- 2411 THEN
            tanh_f := - 1693;
        ELSIF x =- 2410 THEN
            tanh_f := - 1692;
        ELSIF x =- 2409 THEN
            tanh_f := - 1692;
        ELSIF x =- 2408 THEN
            tanh_f := - 1692;
        ELSIF x =- 2407 THEN
            tanh_f := - 1691;
        ELSIF x =- 2406 THEN
            tanh_f := - 1691;
        ELSIF x =- 2405 THEN
            tanh_f := - 1691;
        ELSIF x =- 2404 THEN
            tanh_f := - 1690;
        ELSIF x =- 2403 THEN
            tanh_f := - 1690;
        ELSIF x =- 2402 THEN
            tanh_f := - 1690;
        ELSIF x =- 2401 THEN
            tanh_f := - 1690;
        ELSIF x =- 2400 THEN
            tanh_f := - 1689;
        ELSIF x =- 2399 THEN
            tanh_f := - 1689;
        ELSIF x =- 2398 THEN
            tanh_f := - 1689;
        ELSIF x =- 2397 THEN
            tanh_f := - 1688;
        ELSIF x =- 2396 THEN
            tanh_f := - 1688;
        ELSIF x =- 2395 THEN
            tanh_f := - 1688;
        ELSIF x =- 2394 THEN
            tanh_f := - 1687;
        ELSIF x =- 2393 THEN
            tanh_f := - 1687;
        ELSIF x =- 2392 THEN
            tanh_f := - 1687;
        ELSIF x =- 2391 THEN
            tanh_f := - 1686;
        ELSIF x =- 2390 THEN
            tanh_f := - 1686;
        ELSIF x =- 2389 THEN
            tanh_f := - 1686;
        ELSIF x =- 2388 THEN
            tanh_f := - 1685;
        ELSIF x =- 2387 THEN
            tanh_f := - 1685;
        ELSIF x =- 2386 THEN
            tanh_f := - 1685;
        ELSIF x =- 2385 THEN
            tanh_f := - 1684;
        ELSIF x =- 2384 THEN
            tanh_f := - 1684;
        ELSIF x =- 2383 THEN
            tanh_f := - 1684;
        ELSIF x =- 2382 THEN
            tanh_f := - 1684;
        ELSIF x =- 2381 THEN
            tanh_f := - 1683;
        ELSIF x =- 2380 THEN
            tanh_f := - 1683;
        ELSIF x =- 2379 THEN
            tanh_f := - 1683;
        ELSIF x =- 2378 THEN
            tanh_f := - 1682;
        ELSIF x =- 2377 THEN
            tanh_f := - 1682;
        ELSIF x =- 2376 THEN
            tanh_f := - 1682;
        ELSIF x =- 2375 THEN
            tanh_f := - 1681;
        ELSIF x =- 2374 THEN
            tanh_f := - 1681;
        ELSIF x =- 2373 THEN
            tanh_f := - 1681;
        ELSIF x =- 2372 THEN
            tanh_f := - 1680;
        ELSIF x =- 2371 THEN
            tanh_f := - 1680;
        ELSIF x =- 2370 THEN
            tanh_f := - 1680;
        ELSIF x =- 2369 THEN
            tanh_f := - 1679;
        ELSIF x =- 2368 THEN
            tanh_f := - 1679;
        ELSIF x =- 2367 THEN
            tanh_f := - 1679;
        ELSIF x =- 2366 THEN
            tanh_f := - 1678;
        ELSIF x =- 2365 THEN
            tanh_f := - 1678;
        ELSIF x =- 2364 THEN
            tanh_f := - 1678;
        ELSIF x =- 2363 THEN
            tanh_f := - 1678;
        ELSIF x =- 2362 THEN
            tanh_f := - 1677;
        ELSIF x =- 2361 THEN
            tanh_f := - 1677;
        ELSIF x =- 2360 THEN
            tanh_f := - 1677;
        ELSIF x =- 2359 THEN
            tanh_f := - 1676;
        ELSIF x =- 2358 THEN
            tanh_f := - 1676;
        ELSIF x =- 2357 THEN
            tanh_f := - 1676;
        ELSIF x =- 2356 THEN
            tanh_f := - 1675;
        ELSIF x =- 2355 THEN
            tanh_f := - 1675;
        ELSIF x =- 2354 THEN
            tanh_f := - 1675;
        ELSIF x =- 2353 THEN
            tanh_f := - 1674;
        ELSIF x =- 2352 THEN
            tanh_f := - 1674;
        ELSIF x =- 2351 THEN
            tanh_f := - 1674;
        ELSIF x =- 2350 THEN
            tanh_f := - 1673;
        ELSIF x =- 2349 THEN
            tanh_f := - 1673;
        ELSIF x =- 2348 THEN
            tanh_f := - 1673;
        ELSIF x =- 2347 THEN
            tanh_f := - 1673;
        ELSIF x =- 2346 THEN
            tanh_f := - 1672;
        ELSIF x =- 2345 THEN
            tanh_f := - 1672;
        ELSIF x =- 2344 THEN
            tanh_f := - 1672;
        ELSIF x =- 2343 THEN
            tanh_f := - 1671;
        ELSIF x =- 2342 THEN
            tanh_f := - 1671;
        ELSIF x =- 2341 THEN
            tanh_f := - 1671;
        ELSIF x =- 2340 THEN
            tanh_f := - 1670;
        ELSIF x =- 2339 THEN
            tanh_f := - 1670;
        ELSIF x =- 2338 THEN
            tanh_f := - 1670;
        ELSIF x =- 2337 THEN
            tanh_f := - 1669;
        ELSIF x =- 2336 THEN
            tanh_f := - 1669;
        ELSIF x =- 2335 THEN
            tanh_f := - 1669;
        ELSIF x =- 2334 THEN
            tanh_f := - 1668;
        ELSIF x =- 2333 THEN
            tanh_f := - 1668;
        ELSIF x =- 2332 THEN
            tanh_f := - 1668;
        ELSIF x =- 2331 THEN
            tanh_f := - 1667;
        ELSIF x =- 2330 THEN
            tanh_f := - 1667;
        ELSIF x =- 2329 THEN
            tanh_f := - 1667;
        ELSIF x =- 2328 THEN
            tanh_f := - 1667;
        ELSIF x =- 2327 THEN
            tanh_f := - 1666;
        ELSIF x =- 2326 THEN
            tanh_f := - 1666;
        ELSIF x =- 2325 THEN
            tanh_f := - 1666;
        ELSIF x =- 2324 THEN
            tanh_f := - 1665;
        ELSIF x =- 2323 THEN
            tanh_f := - 1665;
        ELSIF x =- 2322 THEN
            tanh_f := - 1665;
        ELSIF x =- 2321 THEN
            tanh_f := - 1664;
        ELSIF x =- 2320 THEN
            tanh_f := - 1664;
        ELSIF x =- 2319 THEN
            tanh_f := - 1664;
        ELSIF x =- 2318 THEN
            tanh_f := - 1663;
        ELSIF x =- 2317 THEN
            tanh_f := - 1663;
        ELSIF x =- 2316 THEN
            tanh_f := - 1663;
        ELSIF x =- 2315 THEN
            tanh_f := - 1662;
        ELSIF x =- 2314 THEN
            tanh_f := - 1662;
        ELSIF x =- 2313 THEN
            tanh_f := - 1662;
        ELSIF x =- 2312 THEN
            tanh_f := - 1662;
        ELSIF x =- 2311 THEN
            tanh_f := - 1661;
        ELSIF x =- 2310 THEN
            tanh_f := - 1661;
        ELSIF x =- 2309 THEN
            tanh_f := - 1661;
        ELSIF x =- 2308 THEN
            tanh_f := - 1660;
        ELSIF x =- 2307 THEN
            tanh_f := - 1660;
        ELSIF x =- 2306 THEN
            tanh_f := - 1660;
        ELSIF x =- 2305 THEN
            tanh_f := - 1659;
        ELSIF x =- 2304 THEN
            tanh_f := - 1659;
        ELSIF x =- 2303 THEN
            tanh_f := - 1659;
        ELSIF x =- 2302 THEN
            tanh_f := - 1658;
        ELSIF x =- 2301 THEN
            tanh_f := - 1658;
        ELSIF x =- 2300 THEN
            tanh_f := - 1657;
        ELSIF x =- 2299 THEN
            tanh_f := - 1657;
        ELSIF x =- 2298 THEN
            tanh_f := - 1657;
        ELSIF x =- 2297 THEN
            tanh_f := - 1656;
        ELSIF x =- 2296 THEN
            tanh_f := - 1656;
        ELSIF x =- 2295 THEN
            tanh_f := - 1656;
        ELSIF x =- 2294 THEN
            tanh_f := - 1655;
        ELSIF x =- 2293 THEN
            tanh_f := - 1655;
        ELSIF x =- 2292 THEN
            tanh_f := - 1654;
        ELSIF x =- 2291 THEN
            tanh_f := - 1654;
        ELSIF x =- 2290 THEN
            tanh_f := - 1654;
        ELSIF x =- 2289 THEN
            tanh_f := - 1653;
        ELSIF x =- 2288 THEN
            tanh_f := - 1653;
        ELSIF x =- 2287 THEN
            tanh_f := - 1653;
        ELSIF x =- 2286 THEN
            tanh_f := - 1652;
        ELSIF x =- 2285 THEN
            tanh_f := - 1652;
        ELSIF x =- 2284 THEN
            tanh_f := - 1651;
        ELSIF x =- 2283 THEN
            tanh_f := - 1651;
        ELSIF x =- 2282 THEN
            tanh_f := - 1651;
        ELSIF x =- 2281 THEN
            tanh_f := - 1650;
        ELSIF x =- 2280 THEN
            tanh_f := - 1650;
        ELSIF x =- 2279 THEN
            tanh_f := - 1650;
        ELSIF x =- 2278 THEN
            tanh_f := - 1649;
        ELSIF x =- 2277 THEN
            tanh_f := - 1649;
        ELSIF x =- 2276 THEN
            tanh_f := - 1648;
        ELSIF x =- 2275 THEN
            tanh_f := - 1648;
        ELSIF x =- 2274 THEN
            tanh_f := - 1648;
        ELSIF x =- 2273 THEN
            tanh_f := - 1647;
        ELSIF x =- 2272 THEN
            tanh_f := - 1647;
        ELSIF x =- 2271 THEN
            tanh_f := - 1647;
        ELSIF x =- 2270 THEN
            tanh_f := - 1646;
        ELSIF x =- 2269 THEN
            tanh_f := - 1646;
        ELSIF x =- 2268 THEN
            tanh_f := - 1645;
        ELSIF x =- 2267 THEN
            tanh_f := - 1645;
        ELSIF x =- 2266 THEN
            tanh_f := - 1645;
        ELSIF x =- 2265 THEN
            tanh_f := - 1644;
        ELSIF x =- 2264 THEN
            tanh_f := - 1644;
        ELSIF x =- 2263 THEN
            tanh_f := - 1644;
        ELSIF x =- 2262 THEN
            tanh_f := - 1643;
        ELSIF x =- 2261 THEN
            tanh_f := - 1643;
        ELSIF x =- 2260 THEN
            tanh_f := - 1642;
        ELSIF x =- 2259 THEN
            tanh_f := - 1642;
        ELSIF x =- 2258 THEN
            tanh_f := - 1642;
        ELSIF x =- 2257 THEN
            tanh_f := - 1641;
        ELSIF x =- 2256 THEN
            tanh_f := - 1641;
        ELSIF x =- 2255 THEN
            tanh_f := - 1641;
        ELSIF x =- 2254 THEN
            tanh_f := - 1640;
        ELSIF x =- 2253 THEN
            tanh_f := - 1640;
        ELSIF x =- 2252 THEN
            tanh_f := - 1639;
        ELSIF x =- 2251 THEN
            tanh_f := - 1639;
        ELSIF x =- 2250 THEN
            tanh_f := - 1639;
        ELSIF x =- 2249 THEN
            tanh_f := - 1638;
        ELSIF x =- 2248 THEN
            tanh_f := - 1638;
        ELSIF x =- 2247 THEN
            tanh_f := - 1638;
        ELSIF x =- 2246 THEN
            tanh_f := - 1637;
        ELSIF x =- 2245 THEN
            tanh_f := - 1637;
        ELSIF x =- 2244 THEN
            tanh_f := - 1636;
        ELSIF x =- 2243 THEN
            tanh_f := - 1636;
        ELSIF x =- 2242 THEN
            tanh_f := - 1636;
        ELSIF x =- 2241 THEN
            tanh_f := - 1635;
        ELSIF x =- 2240 THEN
            tanh_f := - 1635;
        ELSIF x =- 2239 THEN
            tanh_f := - 1634;
        ELSIF x =- 2238 THEN
            tanh_f := - 1634;
        ELSIF x =- 2237 THEN
            tanh_f := - 1634;
        ELSIF x =- 2236 THEN
            tanh_f := - 1633;
        ELSIF x =- 2235 THEN
            tanh_f := - 1633;
        ELSIF x =- 2234 THEN
            tanh_f := - 1633;
        ELSIF x =- 2233 THEN
            tanh_f := - 1632;
        ELSIF x =- 2232 THEN
            tanh_f := - 1632;
        ELSIF x =- 2231 THEN
            tanh_f := - 1631;
        ELSIF x =- 2230 THEN
            tanh_f := - 1631;
        ELSIF x =- 2229 THEN
            tanh_f := - 1631;
        ELSIF x =- 2228 THEN
            tanh_f := - 1630;
        ELSIF x =- 2227 THEN
            tanh_f := - 1630;
        ELSIF x =- 2226 THEN
            tanh_f := - 1630;
        ELSIF x =- 2225 THEN
            tanh_f := - 1629;
        ELSIF x =- 2224 THEN
            tanh_f := - 1629;
        ELSIF x =- 2223 THEN
            tanh_f := - 1628;
        ELSIF x =- 2222 THEN
            tanh_f := - 1628;
        ELSIF x =- 2221 THEN
            tanh_f := - 1628;
        ELSIF x =- 2220 THEN
            tanh_f := - 1627;
        ELSIF x =- 2219 THEN
            tanh_f := - 1627;
        ELSIF x =- 2218 THEN
            tanh_f := - 1627;
        ELSIF x =- 2217 THEN
            tanh_f := - 1626;
        ELSIF x =- 2216 THEN
            tanh_f := - 1626;
        ELSIF x =- 2215 THEN
            tanh_f := - 1625;
        ELSIF x =- 2214 THEN
            tanh_f := - 1625;
        ELSIF x =- 2213 THEN
            tanh_f := - 1625;
        ELSIF x =- 2212 THEN
            tanh_f := - 1624;
        ELSIF x =- 2211 THEN
            tanh_f := - 1624;
        ELSIF x =- 2210 THEN
            tanh_f := - 1624;
        ELSIF x =- 2209 THEN
            tanh_f := - 1623;
        ELSIF x =- 2208 THEN
            tanh_f := - 1623;
        ELSIF x =- 2207 THEN
            tanh_f := - 1622;
        ELSIF x =- 2206 THEN
            tanh_f := - 1622;
        ELSIF x =- 2205 THEN
            tanh_f := - 1622;
        ELSIF x =- 2204 THEN
            tanh_f := - 1621;
        ELSIF x =- 2203 THEN
            tanh_f := - 1621;
        ELSIF x =- 2202 THEN
            tanh_f := - 1621;
        ELSIF x =- 2201 THEN
            tanh_f := - 1620;
        ELSIF x =- 2200 THEN
            tanh_f := - 1620;
        ELSIF x =- 2199 THEN
            tanh_f := - 1619;
        ELSIF x =- 2198 THEN
            tanh_f := - 1619;
        ELSIF x =- 2197 THEN
            tanh_f := - 1619;
        ELSIF x =- 2196 THEN
            tanh_f := - 1618;
        ELSIF x =- 2195 THEN
            tanh_f := - 1618;
        ELSIF x =- 2194 THEN
            tanh_f := - 1618;
        ELSIF x =- 2193 THEN
            tanh_f := - 1617;
        ELSIF x =- 2192 THEN
            tanh_f := - 1617;
        ELSIF x =- 2191 THEN
            tanh_f := - 1616;
        ELSIF x =- 2190 THEN
            tanh_f := - 1616;
        ELSIF x =- 2189 THEN
            tanh_f := - 1616;
        ELSIF x =- 2188 THEN
            tanh_f := - 1615;
        ELSIF x =- 2187 THEN
            tanh_f := - 1615;
        ELSIF x =- 2186 THEN
            tanh_f := - 1615;
        ELSIF x =- 2185 THEN
            tanh_f := - 1614;
        ELSIF x =- 2184 THEN
            tanh_f := - 1614;
        ELSIF x =- 2183 THEN
            tanh_f := - 1613;
        ELSIF x =- 2182 THEN
            tanh_f := - 1613;
        ELSIF x =- 2181 THEN
            tanh_f := - 1613;
        ELSIF x =- 2180 THEN
            tanh_f := - 1612;
        ELSIF x =- 2179 THEN
            tanh_f := - 1612;
        ELSIF x =- 2178 THEN
            tanh_f := - 1612;
        ELSIF x =- 2177 THEN
            tanh_f := - 1611;
        ELSIF x =- 2176 THEN
            tanh_f := - 1611;
        ELSIF x =- 2175 THEN
            tanh_f := - 1610;
        ELSIF x =- 2174 THEN
            tanh_f := - 1610;
        ELSIF x =- 2173 THEN
            tanh_f := - 1610;
        ELSIF x =- 2172 THEN
            tanh_f := - 1609;
        ELSIF x =- 2171 THEN
            tanh_f := - 1609;
        ELSIF x =- 2170 THEN
            tanh_f := - 1608;
        ELSIF x =- 2169 THEN
            tanh_f := - 1608;
        ELSIF x =- 2168 THEN
            tanh_f := - 1608;
        ELSIF x =- 2167 THEN
            tanh_f := - 1607;
        ELSIF x =- 2166 THEN
            tanh_f := - 1607;
        ELSIF x =- 2165 THEN
            tanh_f := - 1607;
        ELSIF x =- 2164 THEN
            tanh_f := - 1606;
        ELSIF x =- 2163 THEN
            tanh_f := - 1606;
        ELSIF x =- 2162 THEN
            tanh_f := - 1605;
        ELSIF x =- 2161 THEN
            tanh_f := - 1605;
        ELSIF x =- 2160 THEN
            tanh_f := - 1605;
        ELSIF x =- 2159 THEN
            tanh_f := - 1604;
        ELSIF x =- 2158 THEN
            tanh_f := - 1604;
        ELSIF x =- 2157 THEN
            tanh_f := - 1604;
        ELSIF x =- 2156 THEN
            tanh_f := - 1603;
        ELSIF x =- 2155 THEN
            tanh_f := - 1603;
        ELSIF x =- 2154 THEN
            tanh_f := - 1602;
        ELSIF x =- 2153 THEN
            tanh_f := - 1602;
        ELSIF x =- 2152 THEN
            tanh_f := - 1602;
        ELSIF x =- 2151 THEN
            tanh_f := - 1601;
        ELSIF x =- 2150 THEN
            tanh_f := - 1601;
        ELSIF x =- 2149 THEN
            tanh_f := - 1601;
        ELSIF x =- 2148 THEN
            tanh_f := - 1600;
        ELSIF x =- 2147 THEN
            tanh_f := - 1600;
        ELSIF x =- 2146 THEN
            tanh_f := - 1599;
        ELSIF x =- 2145 THEN
            tanh_f := - 1599;
        ELSIF x =- 2144 THEN
            tanh_f := - 1599;
        ELSIF x =- 2143 THEN
            tanh_f := - 1598;
        ELSIF x =- 2142 THEN
            tanh_f := - 1598;
        ELSIF x =- 2141 THEN
            tanh_f := - 1598;
        ELSIF x =- 2140 THEN
            tanh_f := - 1597;
        ELSIF x =- 2139 THEN
            tanh_f := - 1597;
        ELSIF x =- 2138 THEN
            tanh_f := - 1596;
        ELSIF x =- 2137 THEN
            tanh_f := - 1596;
        ELSIF x =- 2136 THEN
            tanh_f := - 1596;
        ELSIF x =- 2135 THEN
            tanh_f := - 1595;
        ELSIF x =- 2134 THEN
            tanh_f := - 1595;
        ELSIF x =- 2133 THEN
            tanh_f := - 1595;
        ELSIF x =- 2132 THEN
            tanh_f := - 1594;
        ELSIF x =- 2131 THEN
            tanh_f := - 1594;
        ELSIF x =- 2130 THEN
            tanh_f := - 1593;
        ELSIF x =- 2129 THEN
            tanh_f := - 1593;
        ELSIF x =- 2128 THEN
            tanh_f := - 1593;
        ELSIF x =- 2127 THEN
            tanh_f := - 1592;
        ELSIF x =- 2126 THEN
            tanh_f := - 1592;
        ELSIF x =- 2125 THEN
            tanh_f := - 1592;
        ELSIF x =- 2124 THEN
            tanh_f := - 1591;
        ELSIF x =- 2123 THEN
            tanh_f := - 1591;
        ELSIF x =- 2122 THEN
            tanh_f := - 1590;
        ELSIF x =- 2121 THEN
            tanh_f := - 1590;
        ELSIF x =- 2120 THEN
            tanh_f := - 1590;
        ELSIF x =- 2119 THEN
            tanh_f := - 1589;
        ELSIF x =- 2118 THEN
            tanh_f := - 1589;
        ELSIF x =- 2117 THEN
            tanh_f := - 1589;
        ELSIF x =- 2116 THEN
            tanh_f := - 1588;
        ELSIF x =- 2115 THEN
            tanh_f := - 1588;
        ELSIF x =- 2114 THEN
            tanh_f := - 1587;
        ELSIF x =- 2113 THEN
            tanh_f := - 1587;
        ELSIF x =- 2112 THEN
            tanh_f := - 1587;
        ELSIF x =- 2111 THEN
            tanh_f := - 1586;
        ELSIF x =- 2110 THEN
            tanh_f := - 1586;
        ELSIF x =- 2109 THEN
            tanh_f := - 1585;
        ELSIF x =- 2108 THEN
            tanh_f := - 1585;
        ELSIF x =- 2107 THEN
            tanh_f := - 1585;
        ELSIF x =- 2106 THEN
            tanh_f := - 1584;
        ELSIF x =- 2105 THEN
            tanh_f := - 1584;
        ELSIF x =- 2104 THEN
            tanh_f := - 1584;
        ELSIF x =- 2103 THEN
            tanh_f := - 1583;
        ELSIF x =- 2102 THEN
            tanh_f := - 1583;
        ELSIF x =- 2101 THEN
            tanh_f := - 1582;
        ELSIF x =- 2100 THEN
            tanh_f := - 1582;
        ELSIF x =- 2099 THEN
            tanh_f := - 1582;
        ELSIF x =- 2098 THEN
            tanh_f := - 1581;
        ELSIF x =- 2097 THEN
            tanh_f := - 1581;
        ELSIF x =- 2096 THEN
            tanh_f := - 1581;
        ELSIF x =- 2095 THEN
            tanh_f := - 1580;
        ELSIF x =- 2094 THEN
            tanh_f := - 1580;
        ELSIF x =- 2093 THEN
            tanh_f := - 1579;
        ELSIF x =- 2092 THEN
            tanh_f := - 1579;
        ELSIF x =- 2091 THEN
            tanh_f := - 1579;
        ELSIF x =- 2090 THEN
            tanh_f := - 1578;
        ELSIF x =- 2089 THEN
            tanh_f := - 1578;
        ELSIF x =- 2088 THEN
            tanh_f := - 1578;
        ELSIF x =- 2087 THEN
            tanh_f := - 1577;
        ELSIF x =- 2086 THEN
            tanh_f := - 1577;
        ELSIF x =- 2085 THEN
            tanh_f := - 1576;
        ELSIF x =- 2084 THEN
            tanh_f := - 1576;
        ELSIF x =- 2083 THEN
            tanh_f := - 1576;
        ELSIF x =- 2082 THEN
            tanh_f := - 1575;
        ELSIF x =- 2081 THEN
            tanh_f := - 1575;
        ELSIF x =- 2080 THEN
            tanh_f := - 1575;
        ELSIF x =- 2079 THEN
            tanh_f := - 1574;
        ELSIF x =- 2078 THEN
            tanh_f := - 1574;
        ELSIF x =- 2077 THEN
            tanh_f := - 1573;
        ELSIF x =- 2076 THEN
            tanh_f := - 1573;
        ELSIF x =- 2075 THEN
            tanh_f := - 1573;
        ELSIF x =- 2074 THEN
            tanh_f := - 1572;
        ELSIF x =- 2073 THEN
            tanh_f := - 1572;
        ELSIF x =- 2072 THEN
            tanh_f := - 1572;
        ELSIF x =- 2071 THEN
            tanh_f := - 1571;
        ELSIF x =- 2070 THEN
            tanh_f := - 1571;
        ELSIF x =- 2069 THEN
            tanh_f := - 1570;
        ELSIF x =- 2068 THEN
            tanh_f := - 1570;
        ELSIF x =- 2067 THEN
            tanh_f := - 1570;
        ELSIF x =- 2066 THEN
            tanh_f := - 1569;
        ELSIF x =- 2065 THEN
            tanh_f := - 1569;
        ELSIF x =- 2064 THEN
            tanh_f := - 1569;
        ELSIF x =- 2063 THEN
            tanh_f := - 1568;
        ELSIF x =- 2062 THEN
            tanh_f := - 1568;
        ELSIF x =- 2061 THEN
            tanh_f := - 1567;
        ELSIF x =- 2060 THEN
            tanh_f := - 1567;
        ELSIF x =- 2059 THEN
            tanh_f := - 1567;
        ELSIF x =- 2058 THEN
            tanh_f := - 1566;
        ELSIF x =- 2057 THEN
            tanh_f := - 1566;
        ELSIF x =- 2056 THEN
            tanh_f := - 1566;
        ELSIF x =- 2055 THEN
            tanh_f := - 1565;
        ELSIF x =- 2054 THEN
            tanh_f := - 1565;
        ELSIF x =- 2053 THEN
            tanh_f := - 1564;
        ELSIF x =- 2052 THEN
            tanh_f := - 1564;
        ELSIF x =- 2051 THEN
            tanh_f := - 1564;
        ELSIF x =- 2050 THEN
            tanh_f := - 1563;
        ELSIF x =- 2049 THEN
            tanh_f := - 1563;
        ELSIF x =- 2048 THEN
            tanh_f := - 1562;
        ELSIF x =- 2047 THEN
            tanh_f := - 1562;
        ELSIF x =- 2046 THEN
            tanh_f := - 1562;
        ELSIF x =- 2045 THEN
            tanh_f := - 1561;
        ELSIF x =- 2044 THEN
            tanh_f := - 1561;
        ELSIF x =- 2043 THEN
            tanh_f := - 1560;
        ELSIF x =- 2042 THEN
            tanh_f := - 1560;
        ELSIF x =- 2041 THEN
            tanh_f := - 1559;
        ELSIF x =- 2040 THEN
            tanh_f := - 1559;
        ELSIF x =- 2039 THEN
            tanh_f := - 1558;
        ELSIF x =- 2038 THEN
            tanh_f := - 1558;
        ELSIF x =- 2037 THEN
            tanh_f := - 1557;
        ELSIF x =- 2036 THEN
            tanh_f := - 1557;
        ELSIF x =- 2035 THEN
            tanh_f := - 1556;
        ELSIF x =- 2034 THEN
            tanh_f := - 1556;
        ELSIF x =- 2033 THEN
            tanh_f := - 1556;
        ELSIF x =- 2032 THEN
            tanh_f := - 1555;
        ELSIF x =- 2031 THEN
            tanh_f := - 1555;
        ELSIF x =- 2030 THEN
            tanh_f := - 1554;
        ELSIF x =- 2029 THEN
            tanh_f := - 1554;
        ELSIF x =- 2028 THEN
            tanh_f := - 1553;
        ELSIF x =- 2027 THEN
            tanh_f := - 1553;
        ELSIF x =- 2026 THEN
            tanh_f := - 1552;
        ELSIF x =- 2025 THEN
            tanh_f := - 1552;
        ELSIF x =- 2024 THEN
            tanh_f := - 1551;
        ELSIF x =- 2023 THEN
            tanh_f := - 1551;
        ELSIF x =- 2022 THEN
            tanh_f := - 1550;
        ELSIF x =- 2021 THEN
            tanh_f := - 1550;
        ELSIF x =- 2020 THEN
            tanh_f := - 1549;
        ELSIF x =- 2019 THEN
            tanh_f := - 1549;
        ELSIF x =- 2018 THEN
            tanh_f := - 1549;
        ELSIF x =- 2017 THEN
            tanh_f := - 1548;
        ELSIF x =- 2016 THEN
            tanh_f := - 1548;
        ELSIF x =- 2015 THEN
            tanh_f := - 1547;
        ELSIF x =- 2014 THEN
            tanh_f := - 1547;
        ELSIF x =- 2013 THEN
            tanh_f := - 1546;
        ELSIF x =- 2012 THEN
            tanh_f := - 1546;
        ELSIF x =- 2011 THEN
            tanh_f := - 1545;
        ELSIF x =- 2010 THEN
            tanh_f := - 1545;
        ELSIF x =- 2009 THEN
            tanh_f := - 1544;
        ELSIF x =- 2008 THEN
            tanh_f := - 1544;
        ELSIF x =- 2007 THEN
            tanh_f := - 1543;
        ELSIF x =- 2006 THEN
            tanh_f := - 1543;
        ELSIF x =- 2005 THEN
            tanh_f := - 1543;
        ELSIF x =- 2004 THEN
            tanh_f := - 1542;
        ELSIF x =- 2003 THEN
            tanh_f := - 1542;
        ELSIF x =- 2002 THEN
            tanh_f := - 1541;
        ELSIF x =- 2001 THEN
            tanh_f := - 1541;
        ELSIF x =- 2000 THEN
            tanh_f := - 1540;
        ELSIF x =- 1999 THEN
            tanh_f := - 1540;
        ELSIF x =- 1998 THEN
            tanh_f := - 1539;
        ELSIF x =- 1997 THEN
            tanh_f := - 1539;
        ELSIF x =- 1996 THEN
            tanh_f := - 1538;
        ELSIF x =- 1995 THEN
            tanh_f := - 1538;
        ELSIF x =- 1994 THEN
            tanh_f := - 1537;
        ELSIF x =- 1993 THEN
            tanh_f := - 1537;
        ELSIF x =- 1992 THEN
            tanh_f := - 1536;
        ELSIF x =- 1991 THEN
            tanh_f := - 1536;
        ELSIF x =- 1990 THEN
            tanh_f := - 1536;
        ELSIF x =- 1989 THEN
            tanh_f := - 1535;
        ELSIF x =- 1988 THEN
            tanh_f := - 1535;
        ELSIF x =- 1987 THEN
            tanh_f := - 1534;
        ELSIF x =- 1986 THEN
            tanh_f := - 1534;
        ELSIF x =- 1985 THEN
            tanh_f := - 1533;
        ELSIF x =- 1984 THEN
            tanh_f := - 1533;
        ELSIF x =- 1983 THEN
            tanh_f := - 1532;
        ELSIF x =- 1982 THEN
            tanh_f := - 1532;
        ELSIF x =- 1981 THEN
            tanh_f := - 1531;
        ELSIF x =- 1980 THEN
            tanh_f := - 1531;
        ELSIF x =- 1979 THEN
            tanh_f := - 1530;
        ELSIF x =- 1978 THEN
            tanh_f := - 1530;
        ELSIF x =- 1977 THEN
            tanh_f := - 1529;
        ELSIF x =- 1976 THEN
            tanh_f := - 1529;
        ELSIF x =- 1975 THEN
            tanh_f := - 1529;
        ELSIF x =- 1974 THEN
            tanh_f := - 1528;
        ELSIF x =- 1973 THEN
            tanh_f := - 1528;
        ELSIF x =- 1972 THEN
            tanh_f := - 1527;
        ELSIF x =- 1971 THEN
            tanh_f := - 1527;
        ELSIF x =- 1970 THEN
            tanh_f := - 1526;
        ELSIF x =- 1969 THEN
            tanh_f := - 1526;
        ELSIF x =- 1968 THEN
            tanh_f := - 1525;
        ELSIF x =- 1967 THEN
            tanh_f := - 1525;
        ELSIF x =- 1966 THEN
            tanh_f := - 1524;
        ELSIF x =- 1965 THEN
            tanh_f := - 1524;
        ELSIF x =- 1964 THEN
            tanh_f := - 1523;
        ELSIF x =- 1963 THEN
            tanh_f := - 1523;
        ELSIF x =- 1962 THEN
            tanh_f := - 1523;
        ELSIF x =- 1961 THEN
            tanh_f := - 1522;
        ELSIF x =- 1960 THEN
            tanh_f := - 1522;
        ELSIF x =- 1959 THEN
            tanh_f := - 1521;
        ELSIF x =- 1958 THEN
            tanh_f := - 1521;
        ELSIF x =- 1957 THEN
            tanh_f := - 1520;
        ELSIF x =- 1956 THEN
            tanh_f := - 1520;
        ELSIF x =- 1955 THEN
            tanh_f := - 1519;
        ELSIF x =- 1954 THEN
            tanh_f := - 1519;
        ELSIF x =- 1953 THEN
            tanh_f := - 1518;
        ELSIF x =- 1952 THEN
            tanh_f := - 1518;
        ELSIF x =- 1951 THEN
            tanh_f := - 1517;
        ELSIF x =- 1950 THEN
            tanh_f := - 1517;
        ELSIF x =- 1949 THEN
            tanh_f := - 1516;
        ELSIF x =- 1948 THEN
            tanh_f := - 1516;
        ELSIF x =- 1947 THEN
            tanh_f := - 1516;
        ELSIF x =- 1946 THEN
            tanh_f := - 1515;
        ELSIF x =- 1945 THEN
            tanh_f := - 1515;
        ELSIF x =- 1944 THEN
            tanh_f := - 1514;
        ELSIF x =- 1943 THEN
            tanh_f := - 1514;
        ELSIF x =- 1942 THEN
            tanh_f := - 1513;
        ELSIF x =- 1941 THEN
            tanh_f := - 1513;
        ELSIF x =- 1940 THEN
            tanh_f := - 1512;
        ELSIF x =- 1939 THEN
            tanh_f := - 1512;
        ELSIF x =- 1938 THEN
            tanh_f := - 1511;
        ELSIF x =- 1937 THEN
            tanh_f := - 1511;
        ELSIF x =- 1936 THEN
            tanh_f := - 1510;
        ELSIF x =- 1935 THEN
            tanh_f := - 1510;
        ELSIF x =- 1934 THEN
            tanh_f := - 1510;
        ELSIF x =- 1933 THEN
            tanh_f := - 1509;
        ELSIF x =- 1932 THEN
            tanh_f := - 1509;
        ELSIF x =- 1931 THEN
            tanh_f := - 1508;
        ELSIF x =- 1930 THEN
            tanh_f := - 1508;
        ELSIF x =- 1929 THEN
            tanh_f := - 1507;
        ELSIF x =- 1928 THEN
            tanh_f := - 1507;
        ELSIF x =- 1927 THEN
            tanh_f := - 1506;
        ELSIF x =- 1926 THEN
            tanh_f := - 1506;
        ELSIF x =- 1925 THEN
            tanh_f := - 1505;
        ELSIF x =- 1924 THEN
            tanh_f := - 1505;
        ELSIF x =- 1923 THEN
            tanh_f := - 1504;
        ELSIF x =- 1922 THEN
            tanh_f := - 1504;
        ELSIF x =- 1921 THEN
            tanh_f := - 1503;
        ELSIF x =- 1920 THEN
            tanh_f := - 1503;
        ELSIF x =- 1919 THEN
            tanh_f := - 1503;
        ELSIF x =- 1918 THEN
            tanh_f := - 1502;
        ELSIF x =- 1917 THEN
            tanh_f := - 1502;
        ELSIF x =- 1916 THEN
            tanh_f := - 1501;
        ELSIF x =- 1915 THEN
            tanh_f := - 1501;
        ELSIF x =- 1914 THEN
            tanh_f := - 1500;
        ELSIF x =- 1913 THEN
            tanh_f := - 1500;
        ELSIF x =- 1912 THEN
            tanh_f := - 1499;
        ELSIF x =- 1911 THEN
            tanh_f := - 1499;
        ELSIF x =- 1910 THEN
            tanh_f := - 1498;
        ELSIF x =- 1909 THEN
            tanh_f := - 1498;
        ELSIF x =- 1908 THEN
            tanh_f := - 1497;
        ELSIF x =- 1907 THEN
            tanh_f := - 1497;
        ELSIF x =- 1906 THEN
            tanh_f := - 1496;
        ELSIF x =- 1905 THEN
            tanh_f := - 1496;
        ELSIF x =- 1904 THEN
            tanh_f := - 1496;
        ELSIF x =- 1903 THEN
            tanh_f := - 1495;
        ELSIF x =- 1902 THEN
            tanh_f := - 1495;
        ELSIF x =- 1901 THEN
            tanh_f := - 1494;
        ELSIF x =- 1900 THEN
            tanh_f := - 1494;
        ELSIF x =- 1899 THEN
            tanh_f := - 1493;
        ELSIF x =- 1898 THEN
            tanh_f := - 1493;
        ELSIF x =- 1897 THEN
            tanh_f := - 1492;
        ELSIF x =- 1896 THEN
            tanh_f := - 1492;
        ELSIF x =- 1895 THEN
            tanh_f := - 1491;
        ELSIF x =- 1894 THEN
            tanh_f := - 1491;
        ELSIF x =- 1893 THEN
            tanh_f := - 1490;
        ELSIF x =- 1892 THEN
            tanh_f := - 1490;
        ELSIF x =- 1891 THEN
            tanh_f := - 1490;
        ELSIF x =- 1890 THEN
            tanh_f := - 1489;
        ELSIF x =- 1889 THEN
            tanh_f := - 1489;
        ELSIF x =- 1888 THEN
            tanh_f := - 1488;
        ELSIF x =- 1887 THEN
            tanh_f := - 1488;
        ELSIF x =- 1886 THEN
            tanh_f := - 1487;
        ELSIF x =- 1885 THEN
            tanh_f := - 1487;
        ELSIF x =- 1884 THEN
            tanh_f := - 1486;
        ELSIF x =- 1883 THEN
            tanh_f := - 1486;
        ELSIF x =- 1882 THEN
            tanh_f := - 1485;
        ELSIF x =- 1881 THEN
            tanh_f := - 1485;
        ELSIF x =- 1880 THEN
            tanh_f := - 1484;
        ELSIF x =- 1879 THEN
            tanh_f := - 1484;
        ELSIF x =- 1878 THEN
            tanh_f := - 1483;
        ELSIF x =- 1877 THEN
            tanh_f := - 1483;
        ELSIF x =- 1876 THEN
            tanh_f := - 1483;
        ELSIF x =- 1875 THEN
            tanh_f := - 1482;
        ELSIF x =- 1874 THEN
            tanh_f := - 1482;
        ELSIF x =- 1873 THEN
            tanh_f := - 1481;
        ELSIF x =- 1872 THEN
            tanh_f := - 1481;
        ELSIF x =- 1871 THEN
            tanh_f := - 1480;
        ELSIF x =- 1870 THEN
            tanh_f := - 1480;
        ELSIF x =- 1869 THEN
            tanh_f := - 1479;
        ELSIF x =- 1868 THEN
            tanh_f := - 1479;
        ELSIF x =- 1867 THEN
            tanh_f := - 1478;
        ELSIF x =- 1866 THEN
            tanh_f := - 1478;
        ELSIF x =- 1865 THEN
            tanh_f := - 1477;
        ELSIF x =- 1864 THEN
            tanh_f := - 1477;
        ELSIF x =- 1863 THEN
            tanh_f := - 1477;
        ELSIF x =- 1862 THEN
            tanh_f := - 1476;
        ELSIF x =- 1861 THEN
            tanh_f := - 1476;
        ELSIF x =- 1860 THEN
            tanh_f := - 1475;
        ELSIF x =- 1859 THEN
            tanh_f := - 1475;
        ELSIF x =- 1858 THEN
            tanh_f := - 1474;
        ELSIF x =- 1857 THEN
            tanh_f := - 1474;
        ELSIF x =- 1856 THEN
            tanh_f := - 1473;
        ELSIF x =- 1855 THEN
            tanh_f := - 1473;
        ELSIF x =- 1854 THEN
            tanh_f := - 1472;
        ELSIF x =- 1853 THEN
            tanh_f := - 1472;
        ELSIF x =- 1852 THEN
            tanh_f := - 1471;
        ELSIF x =- 1851 THEN
            tanh_f := - 1471;
        ELSIF x =- 1850 THEN
            tanh_f := - 1470;
        ELSIF x =- 1849 THEN
            tanh_f := - 1470;
        ELSIF x =- 1848 THEN
            tanh_f := - 1470;
        ELSIF x =- 1847 THEN
            tanh_f := - 1469;
        ELSIF x =- 1846 THEN
            tanh_f := - 1469;
        ELSIF x =- 1845 THEN
            tanh_f := - 1468;
        ELSIF x =- 1844 THEN
            tanh_f := - 1468;
        ELSIF x =- 1843 THEN
            tanh_f := - 1467;
        ELSIF x =- 1842 THEN
            tanh_f := - 1467;
        ELSIF x =- 1841 THEN
            tanh_f := - 1466;
        ELSIF x =- 1840 THEN
            tanh_f := - 1466;
        ELSIF x =- 1839 THEN
            tanh_f := - 1465;
        ELSIF x =- 1838 THEN
            tanh_f := - 1465;
        ELSIF x =- 1837 THEN
            tanh_f := - 1464;
        ELSIF x =- 1836 THEN
            tanh_f := - 1464;
        ELSIF x =- 1835 THEN
            tanh_f := - 1463;
        ELSIF x =- 1834 THEN
            tanh_f := - 1463;
        ELSIF x =- 1833 THEN
            tanh_f := - 1463;
        ELSIF x =- 1832 THEN
            tanh_f := - 1462;
        ELSIF x =- 1831 THEN
            tanh_f := - 1462;
        ELSIF x =- 1830 THEN
            tanh_f := - 1461;
        ELSIF x =- 1829 THEN
            tanh_f := - 1461;
        ELSIF x =- 1828 THEN
            tanh_f := - 1460;
        ELSIF x =- 1827 THEN
            tanh_f := - 1460;
        ELSIF x =- 1826 THEN
            tanh_f := - 1459;
        ELSIF x =- 1825 THEN
            tanh_f := - 1459;
        ELSIF x =- 1824 THEN
            tanh_f := - 1458;
        ELSIF x =- 1823 THEN
            tanh_f := - 1458;
        ELSIF x =- 1822 THEN
            tanh_f := - 1457;
        ELSIF x =- 1821 THEN
            tanh_f := - 1457;
        ELSIF x =- 1820 THEN
            tanh_f := - 1457;
        ELSIF x =- 1819 THEN
            tanh_f := - 1456;
        ELSIF x =- 1818 THEN
            tanh_f := - 1456;
        ELSIF x =- 1817 THEN
            tanh_f := - 1455;
        ELSIF x =- 1816 THEN
            tanh_f := - 1455;
        ELSIF x =- 1815 THEN
            tanh_f := - 1454;
        ELSIF x =- 1814 THEN
            tanh_f := - 1454;
        ELSIF x =- 1813 THEN
            tanh_f := - 1453;
        ELSIF x =- 1812 THEN
            tanh_f := - 1453;
        ELSIF x =- 1811 THEN
            tanh_f := - 1452;
        ELSIF x =- 1810 THEN
            tanh_f := - 1452;
        ELSIF x =- 1809 THEN
            tanh_f := - 1451;
        ELSIF x =- 1808 THEN
            tanh_f := - 1451;
        ELSIF x =- 1807 THEN
            tanh_f := - 1450;
        ELSIF x =- 1806 THEN
            tanh_f := - 1450;
        ELSIF x =- 1805 THEN
            tanh_f := - 1450;
        ELSIF x =- 1804 THEN
            tanh_f := - 1449;
        ELSIF x =- 1803 THEN
            tanh_f := - 1449;
        ELSIF x =- 1802 THEN
            tanh_f := - 1448;
        ELSIF x =- 1801 THEN
            tanh_f := - 1448;
        ELSIF x =- 1800 THEN
            tanh_f := - 1447;
        ELSIF x =- 1799 THEN
            tanh_f := - 1447;
        ELSIF x =- 1798 THEN
            tanh_f := - 1446;
        ELSIF x =- 1797 THEN
            tanh_f := - 1446;
        ELSIF x =- 1796 THEN
            tanh_f := - 1445;
        ELSIF x =- 1795 THEN
            tanh_f := - 1445;
        ELSIF x =- 1794 THEN
            tanh_f := - 1444;
        ELSIF x =- 1793 THEN
            tanh_f := - 1444;
        ELSIF x =- 1792 THEN
            tanh_f := - 1443;
        ELSIF x =- 1791 THEN
            tanh_f := - 1443;
        ELSIF x =- 1790 THEN
            tanh_f := - 1443;
        ELSIF x =- 1789 THEN
            tanh_f := - 1442;
        ELSIF x =- 1788 THEN
            tanh_f := - 1442;
        ELSIF x =- 1787 THEN
            tanh_f := - 1441;
        ELSIF x =- 1786 THEN
            tanh_f := - 1441;
        ELSIF x =- 1785 THEN
            tanh_f := - 1440;
        ELSIF x =- 1784 THEN
            tanh_f := - 1440;
        ELSIF x =- 1783 THEN
            tanh_f := - 1439;
        ELSIF x =- 1782 THEN
            tanh_f := - 1439;
        ELSIF x =- 1781 THEN
            tanh_f := - 1438;
        ELSIF x =- 1780 THEN
            tanh_f := - 1437;
        ELSIF x =- 1779 THEN
            tanh_f := - 1437;
        ELSIF x =- 1778 THEN
            tanh_f := - 1436;
        ELSIF x =- 1777 THEN
            tanh_f := - 1436;
        ELSIF x =- 1776 THEN
            tanh_f := - 1435;
        ELSIF x =- 1775 THEN
            tanh_f := - 1435;
        ELSIF x =- 1774 THEN
            tanh_f := - 1434;
        ELSIF x =- 1773 THEN
            tanh_f := - 1434;
        ELSIF x =- 1772 THEN
            tanh_f := - 1433;
        ELSIF x =- 1771 THEN
            tanh_f := - 1432;
        ELSIF x =- 1770 THEN
            tanh_f := - 1432;
        ELSIF x =- 1769 THEN
            tanh_f := - 1431;
        ELSIF x =- 1768 THEN
            tanh_f := - 1431;
        ELSIF x =- 1767 THEN
            tanh_f := - 1430;
        ELSIF x =- 1766 THEN
            tanh_f := - 1430;
        ELSIF x =- 1765 THEN
            tanh_f := - 1429;
        ELSIF x =- 1764 THEN
            tanh_f := - 1429;
        ELSIF x =- 1763 THEN
            tanh_f := - 1428;
        ELSIF x =- 1762 THEN
            tanh_f := - 1428;
        ELSIF x =- 1761 THEN
            tanh_f := - 1427;
        ELSIF x =- 1760 THEN
            tanh_f := - 1426;
        ELSIF x =- 1759 THEN
            tanh_f := - 1426;
        ELSIF x =- 1758 THEN
            tanh_f := - 1425;
        ELSIF x =- 1757 THEN
            tanh_f := - 1425;
        ELSIF x =- 1756 THEN
            tanh_f := - 1424;
        ELSIF x =- 1755 THEN
            tanh_f := - 1424;
        ELSIF x =- 1754 THEN
            tanh_f := - 1423;
        ELSIF x =- 1753 THEN
            tanh_f := - 1423;
        ELSIF x =- 1752 THEN
            tanh_f := - 1422;
        ELSIF x =- 1751 THEN
            tanh_f := - 1421;
        ELSIF x =- 1750 THEN
            tanh_f := - 1421;
        ELSIF x =- 1749 THEN
            tanh_f := - 1420;
        ELSIF x =- 1748 THEN
            tanh_f := - 1420;
        ELSIF x =- 1747 THEN
            tanh_f := - 1419;
        ELSIF x =- 1746 THEN
            tanh_f := - 1419;
        ELSIF x =- 1745 THEN
            tanh_f := - 1418;
        ELSIF x =- 1744 THEN
            tanh_f := - 1418;
        ELSIF x =- 1743 THEN
            tanh_f := - 1417;
        ELSIF x =- 1742 THEN
            tanh_f := - 1417;
        ELSIF x =- 1741 THEN
            tanh_f := - 1416;
        ELSIF x =- 1740 THEN
            tanh_f := - 1415;
        ELSIF x =- 1739 THEN
            tanh_f := - 1415;
        ELSIF x =- 1738 THEN
            tanh_f := - 1414;
        ELSIF x =- 1737 THEN
            tanh_f := - 1414;
        ELSIF x =- 1736 THEN
            tanh_f := - 1413;
        ELSIF x =- 1735 THEN
            tanh_f := - 1413;
        ELSIF x =- 1734 THEN
            tanh_f := - 1412;
        ELSIF x =- 1733 THEN
            tanh_f := - 1412;
        ELSIF x =- 1732 THEN
            tanh_f := - 1411;
        ELSIF x =- 1731 THEN
            tanh_f := - 1411;
        ELSIF x =- 1730 THEN
            tanh_f := - 1410;
        ELSIF x =- 1729 THEN
            tanh_f := - 1409;
        ELSIF x =- 1728 THEN
            tanh_f := - 1409;
        ELSIF x =- 1727 THEN
            tanh_f := - 1408;
        ELSIF x =- 1726 THEN
            tanh_f := - 1408;
        ELSIF x =- 1725 THEN
            tanh_f := - 1407;
        ELSIF x =- 1724 THEN
            tanh_f := - 1407;
        ELSIF x =- 1723 THEN
            tanh_f := - 1406;
        ELSIF x =- 1722 THEN
            tanh_f := - 1406;
        ELSIF x =- 1721 THEN
            tanh_f := - 1405;
        ELSIF x =- 1720 THEN
            tanh_f := - 1404;
        ELSIF x =- 1719 THEN
            tanh_f := - 1404;
        ELSIF x =- 1718 THEN
            tanh_f := - 1403;
        ELSIF x =- 1717 THEN
            tanh_f := - 1403;
        ELSIF x =- 1716 THEN
            tanh_f := - 1402;
        ELSIF x =- 1715 THEN
            tanh_f := - 1402;
        ELSIF x =- 1714 THEN
            tanh_f := - 1401;
        ELSIF x =- 1713 THEN
            tanh_f := - 1401;
        ELSIF x =- 1712 THEN
            tanh_f := - 1400;
        ELSIF x =- 1711 THEN
            tanh_f := - 1400;
        ELSIF x =- 1710 THEN
            tanh_f := - 1399;
        ELSIF x =- 1709 THEN
            tanh_f := - 1398;
        ELSIF x =- 1708 THEN
            tanh_f := - 1398;
        ELSIF x =- 1707 THEN
            tanh_f := - 1397;
        ELSIF x =- 1706 THEN
            tanh_f := - 1397;
        ELSIF x =- 1705 THEN
            tanh_f := - 1396;
        ELSIF x =- 1704 THEN
            tanh_f := - 1396;
        ELSIF x =- 1703 THEN
            tanh_f := - 1395;
        ELSIF x =- 1702 THEN
            tanh_f := - 1395;
        ELSIF x =- 1701 THEN
            tanh_f := - 1394;
        ELSIF x =- 1700 THEN
            tanh_f := - 1394;
        ELSIF x =- 1699 THEN
            tanh_f := - 1393;
        ELSIF x =- 1698 THEN
            tanh_f := - 1392;
        ELSIF x =- 1697 THEN
            tanh_f := - 1392;
        ELSIF x =- 1696 THEN
            tanh_f := - 1391;
        ELSIF x =- 1695 THEN
            tanh_f := - 1391;
        ELSIF x =- 1694 THEN
            tanh_f := - 1390;
        ELSIF x =- 1693 THEN
            tanh_f := - 1390;
        ELSIF x =- 1692 THEN
            tanh_f := - 1389;
        ELSIF x =- 1691 THEN
            tanh_f := - 1389;
        ELSIF x =- 1690 THEN
            tanh_f := - 1388;
        ELSIF x =- 1689 THEN
            tanh_f := - 1387;
        ELSIF x =- 1688 THEN
            tanh_f := - 1387;
        ELSIF x =- 1687 THEN
            tanh_f := - 1386;
        ELSIF x =- 1686 THEN
            tanh_f := - 1386;
        ELSIF x =- 1685 THEN
            tanh_f := - 1385;
        ELSIF x =- 1684 THEN
            tanh_f := - 1385;
        ELSIF x =- 1683 THEN
            tanh_f := - 1384;
        ELSIF x =- 1682 THEN
            tanh_f := - 1384;
        ELSIF x =- 1681 THEN
            tanh_f := - 1383;
        ELSIF x =- 1680 THEN
            tanh_f := - 1383;
        ELSIF x =- 1679 THEN
            tanh_f := - 1382;
        ELSIF x =- 1678 THEN
            tanh_f := - 1381;
        ELSIF x =- 1677 THEN
            tanh_f := - 1381;
        ELSIF x =- 1676 THEN
            tanh_f := - 1380;
        ELSIF x =- 1675 THEN
            tanh_f := - 1380;
        ELSIF x =- 1674 THEN
            tanh_f := - 1379;
        ELSIF x =- 1673 THEN
            tanh_f := - 1379;
        ELSIF x =- 1672 THEN
            tanh_f := - 1378;
        ELSIF x =- 1671 THEN
            tanh_f := - 1378;
        ELSIF x =- 1670 THEN
            tanh_f := - 1377;
        ELSIF x =- 1669 THEN
            tanh_f := - 1376;
        ELSIF x =- 1668 THEN
            tanh_f := - 1376;
        ELSIF x =- 1667 THEN
            tanh_f := - 1375;
        ELSIF x =- 1666 THEN
            tanh_f := - 1375;
        ELSIF x =- 1665 THEN
            tanh_f := - 1374;
        ELSIF x =- 1664 THEN
            tanh_f := - 1374;
        ELSIF x =- 1663 THEN
            tanh_f := - 1373;
        ELSIF x =- 1662 THEN
            tanh_f := - 1373;
        ELSIF x =- 1661 THEN
            tanh_f := - 1372;
        ELSIF x =- 1660 THEN
            tanh_f := - 1372;
        ELSIF x =- 1659 THEN
            tanh_f := - 1371;
        ELSIF x =- 1658 THEN
            tanh_f := - 1370;
        ELSIF x =- 1657 THEN
            tanh_f := - 1370;
        ELSIF x =- 1656 THEN
            tanh_f := - 1369;
        ELSIF x =- 1655 THEN
            tanh_f := - 1369;
        ELSIF x =- 1654 THEN
            tanh_f := - 1368;
        ELSIF x =- 1653 THEN
            tanh_f := - 1368;
        ELSIF x =- 1652 THEN
            tanh_f := - 1367;
        ELSIF x =- 1651 THEN
            tanh_f := - 1367;
        ELSIF x =- 1650 THEN
            tanh_f := - 1366;
        ELSIF x =- 1649 THEN
            tanh_f := - 1366;
        ELSIF x =- 1648 THEN
            tanh_f := - 1365;
        ELSIF x =- 1647 THEN
            tanh_f := - 1364;
        ELSIF x =- 1646 THEN
            tanh_f := - 1364;
        ELSIF x =- 1645 THEN
            tanh_f := - 1363;
        ELSIF x =- 1644 THEN
            tanh_f := - 1363;
        ELSIF x =- 1643 THEN
            tanh_f := - 1362;
        ELSIF x =- 1642 THEN
            tanh_f := - 1362;
        ELSIF x =- 1641 THEN
            tanh_f := - 1361;
        ELSIF x =- 1640 THEN
            tanh_f := - 1361;
        ELSIF x =- 1639 THEN
            tanh_f := - 1360;
        ELSIF x =- 1638 THEN
            tanh_f := - 1359;
        ELSIF x =- 1637 THEN
            tanh_f := - 1359;
        ELSIF x =- 1636 THEN
            tanh_f := - 1358;
        ELSIF x =- 1635 THEN
            tanh_f := - 1358;
        ELSIF x =- 1634 THEN
            tanh_f := - 1357;
        ELSIF x =- 1633 THEN
            tanh_f := - 1357;
        ELSIF x =- 1632 THEN
            tanh_f := - 1356;
        ELSIF x =- 1631 THEN
            tanh_f := - 1356;
        ELSIF x =- 1630 THEN
            tanh_f := - 1355;
        ELSIF x =- 1629 THEN
            tanh_f := - 1355;
        ELSIF x =- 1628 THEN
            tanh_f := - 1354;
        ELSIF x =- 1627 THEN
            tanh_f := - 1353;
        ELSIF x =- 1626 THEN
            tanh_f := - 1353;
        ELSIF x =- 1625 THEN
            tanh_f := - 1352;
        ELSIF x =- 1624 THEN
            tanh_f := - 1352;
        ELSIF x =- 1623 THEN
            tanh_f := - 1351;
        ELSIF x =- 1622 THEN
            tanh_f := - 1351;
        ELSIF x =- 1621 THEN
            tanh_f := - 1350;
        ELSIF x =- 1620 THEN
            tanh_f := - 1350;
        ELSIF x =- 1619 THEN
            tanh_f := - 1349;
        ELSIF x =- 1618 THEN
            tanh_f := - 1349;
        ELSIF x =- 1617 THEN
            tanh_f := - 1348;
        ELSIF x =- 1616 THEN
            tanh_f := - 1347;
        ELSIF x =- 1615 THEN
            tanh_f := - 1347;
        ELSIF x =- 1614 THEN
            tanh_f := - 1346;
        ELSIF x =- 1613 THEN
            tanh_f := - 1346;
        ELSIF x =- 1612 THEN
            tanh_f := - 1345;
        ELSIF x =- 1611 THEN
            tanh_f := - 1345;
        ELSIF x =- 1610 THEN
            tanh_f := - 1344;
        ELSIF x =- 1609 THEN
            tanh_f := - 1344;
        ELSIF x =- 1608 THEN
            tanh_f := - 1343;
        ELSIF x =- 1607 THEN
            tanh_f := - 1342;
        ELSIF x =- 1606 THEN
            tanh_f := - 1342;
        ELSIF x =- 1605 THEN
            tanh_f := - 1341;
        ELSIF x =- 1604 THEN
            tanh_f := - 1341;
        ELSIF x =- 1603 THEN
            tanh_f := - 1340;
        ELSIF x =- 1602 THEN
            tanh_f := - 1340;
        ELSIF x =- 1601 THEN
            tanh_f := - 1339;
        ELSIF x =- 1600 THEN
            tanh_f := - 1339;
        ELSIF x =- 1599 THEN
            tanh_f := - 1338;
        ELSIF x =- 1598 THEN
            tanh_f := - 1338;
        ELSIF x =- 1597 THEN
            tanh_f := - 1337;
        ELSIF x =- 1596 THEN
            tanh_f := - 1336;
        ELSIF x =- 1595 THEN
            tanh_f := - 1336;
        ELSIF x =- 1594 THEN
            tanh_f := - 1335;
        ELSIF x =- 1593 THEN
            tanh_f := - 1335;
        ELSIF x =- 1592 THEN
            tanh_f := - 1334;
        ELSIF x =- 1591 THEN
            tanh_f := - 1334;
        ELSIF x =- 1590 THEN
            tanh_f := - 1333;
        ELSIF x =- 1589 THEN
            tanh_f := - 1333;
        ELSIF x =- 1588 THEN
            tanh_f := - 1332;
        ELSIF x =- 1587 THEN
            tanh_f := - 1331;
        ELSIF x =- 1586 THEN
            tanh_f := - 1331;
        ELSIF x =- 1585 THEN
            tanh_f := - 1330;
        ELSIF x =- 1584 THEN
            tanh_f := - 1330;
        ELSIF x =- 1583 THEN
            tanh_f := - 1329;
        ELSIF x =- 1582 THEN
            tanh_f := - 1329;
        ELSIF x =- 1581 THEN
            tanh_f := - 1328;
        ELSIF x =- 1580 THEN
            tanh_f := - 1328;
        ELSIF x =- 1579 THEN
            tanh_f := - 1327;
        ELSIF x =- 1578 THEN
            tanh_f := - 1327;
        ELSIF x =- 1577 THEN
            tanh_f := - 1326;
        ELSIF x =- 1576 THEN
            tanh_f := - 1325;
        ELSIF x =- 1575 THEN
            tanh_f := - 1325;
        ELSIF x =- 1574 THEN
            tanh_f := - 1324;
        ELSIF x =- 1573 THEN
            tanh_f := - 1324;
        ELSIF x =- 1572 THEN
            tanh_f := - 1323;
        ELSIF x =- 1571 THEN
            tanh_f := - 1323;
        ELSIF x =- 1570 THEN
            tanh_f := - 1322;
        ELSIF x =- 1569 THEN
            tanh_f := - 1322;
        ELSIF x =- 1568 THEN
            tanh_f := - 1321;
        ELSIF x =- 1567 THEN
            tanh_f := - 1321;
        ELSIF x =- 1566 THEN
            tanh_f := - 1320;
        ELSIF x =- 1565 THEN
            tanh_f := - 1319;
        ELSIF x =- 1564 THEN
            tanh_f := - 1319;
        ELSIF x =- 1563 THEN
            tanh_f := - 1318;
        ELSIF x =- 1562 THEN
            tanh_f := - 1318;
        ELSIF x =- 1561 THEN
            tanh_f := - 1317;
        ELSIF x =- 1560 THEN
            tanh_f := - 1317;
        ELSIF x =- 1559 THEN
            tanh_f := - 1316;
        ELSIF x =- 1558 THEN
            tanh_f := - 1316;
        ELSIF x =- 1557 THEN
            tanh_f := - 1315;
        ELSIF x =- 1556 THEN
            tanh_f := - 1314;
        ELSIF x =- 1555 THEN
            tanh_f := - 1314;
        ELSIF x =- 1554 THEN
            tanh_f := - 1313;
        ELSIF x =- 1553 THEN
            tanh_f := - 1313;
        ELSIF x =- 1552 THEN
            tanh_f := - 1312;
        ELSIF x =- 1551 THEN
            tanh_f := - 1312;
        ELSIF x =- 1550 THEN
            tanh_f := - 1311;
        ELSIF x =- 1549 THEN
            tanh_f := - 1311;
        ELSIF x =- 1548 THEN
            tanh_f := - 1310;
        ELSIF x =- 1547 THEN
            tanh_f := - 1310;
        ELSIF x =- 1546 THEN
            tanh_f := - 1309;
        ELSIF x =- 1545 THEN
            tanh_f := - 1308;
        ELSIF x =- 1544 THEN
            tanh_f := - 1308;
        ELSIF x =- 1543 THEN
            tanh_f := - 1307;
        ELSIF x =- 1542 THEN
            tanh_f := - 1307;
        ELSIF x =- 1541 THEN
            tanh_f := - 1306;
        ELSIF x =- 1540 THEN
            tanh_f := - 1306;
        ELSIF x =- 1539 THEN
            tanh_f := - 1305;
        ELSIF x =- 1538 THEN
            tanh_f := - 1305;
        ELSIF x =- 1537 THEN
            tanh_f := - 1304;
        ELSIF x =- 1536 THEN
            tanh_f := - 1303;
        ELSIF x =- 1535 THEN
            tanh_f := - 1303;
        ELSIF x =- 1534 THEN
            tanh_f := - 1302;
        ELSIF x =- 1533 THEN
            tanh_f := - 1302;
        ELSIF x =- 1532 THEN
            tanh_f := - 1301;
        ELSIF x =- 1531 THEN
            tanh_f := - 1300;
        ELSIF x =- 1530 THEN
            tanh_f := - 1300;
        ELSIF x =- 1529 THEN
            tanh_f := - 1299;
        ELSIF x =- 1528 THEN
            tanh_f := - 1298;
        ELSIF x =- 1527 THEN
            tanh_f := - 1298;
        ELSIF x =- 1526 THEN
            tanh_f := - 1297;
        ELSIF x =- 1525 THEN
            tanh_f := - 1296;
        ELSIF x =- 1524 THEN
            tanh_f := - 1296;
        ELSIF x =- 1523 THEN
            tanh_f := - 1295;
        ELSIF x =- 1522 THEN
            tanh_f := - 1295;
        ELSIF x =- 1521 THEN
            tanh_f := - 1294;
        ELSIF x =- 1520 THEN
            tanh_f := - 1293;
        ELSIF x =- 1519 THEN
            tanh_f := - 1293;
        ELSIF x =- 1518 THEN
            tanh_f := - 1292;
        ELSIF x =- 1517 THEN
            tanh_f := - 1291;
        ELSIF x =- 1516 THEN
            tanh_f := - 1291;
        ELSIF x =- 1515 THEN
            tanh_f := - 1290;
        ELSIF x =- 1514 THEN
            tanh_f := - 1289;
        ELSIF x =- 1513 THEN
            tanh_f := - 1289;
        ELSIF x =- 1512 THEN
            tanh_f := - 1288;
        ELSIF x =- 1511 THEN
            tanh_f := - 1287;
        ELSIF x =- 1510 THEN
            tanh_f := - 1287;
        ELSIF x =- 1509 THEN
            tanh_f := - 1286;
        ELSIF x =- 1508 THEN
            tanh_f := - 1286;
        ELSIF x =- 1507 THEN
            tanh_f := - 1285;
        ELSIF x =- 1506 THEN
            tanh_f := - 1284;
        ELSIF x =- 1505 THEN
            tanh_f := - 1284;
        ELSIF x =- 1504 THEN
            tanh_f := - 1283;
        ELSIF x =- 1503 THEN
            tanh_f := - 1282;
        ELSIF x =- 1502 THEN
            tanh_f := - 1282;
        ELSIF x =- 1501 THEN
            tanh_f := - 1281;
        ELSIF x =- 1500 THEN
            tanh_f := - 1280;
        ELSIF x =- 1499 THEN
            tanh_f := - 1280;
        ELSIF x =- 1498 THEN
            tanh_f := - 1279;
        ELSIF x =- 1497 THEN
            tanh_f := - 1278;
        ELSIF x =- 1496 THEN
            tanh_f := - 1278;
        ELSIF x =- 1495 THEN
            tanh_f := - 1277;
        ELSIF x =- 1494 THEN
            tanh_f := - 1277;
        ELSIF x =- 1493 THEN
            tanh_f := - 1276;
        ELSIF x =- 1492 THEN
            tanh_f := - 1275;
        ELSIF x =- 1491 THEN
            tanh_f := - 1275;
        ELSIF x =- 1490 THEN
            tanh_f := - 1274;
        ELSIF x =- 1489 THEN
            tanh_f := - 1273;
        ELSIF x =- 1488 THEN
            tanh_f := - 1273;
        ELSIF x =- 1487 THEN
            tanh_f := - 1272;
        ELSIF x =- 1486 THEN
            tanh_f := - 1271;
        ELSIF x =- 1485 THEN
            tanh_f := - 1271;
        ELSIF x =- 1484 THEN
            tanh_f := - 1270;
        ELSIF x =- 1483 THEN
            tanh_f := - 1269;
        ELSIF x =- 1482 THEN
            tanh_f := - 1269;
        ELSIF x =- 1481 THEN
            tanh_f := - 1268;
        ELSIF x =- 1480 THEN
            tanh_f := - 1268;
        ELSIF x =- 1479 THEN
            tanh_f := - 1267;
        ELSIF x =- 1478 THEN
            tanh_f := - 1266;
        ELSIF x =- 1477 THEN
            tanh_f := - 1266;
        ELSIF x =- 1476 THEN
            tanh_f := - 1265;
        ELSIF x =- 1475 THEN
            tanh_f := - 1264;
        ELSIF x =- 1474 THEN
            tanh_f := - 1264;
        ELSIF x =- 1473 THEN
            tanh_f := - 1263;
        ELSIF x =- 1472 THEN
            tanh_f := - 1262;
        ELSIF x =- 1471 THEN
            tanh_f := - 1262;
        ELSIF x =- 1470 THEN
            tanh_f := - 1261;
        ELSIF x =- 1469 THEN
            tanh_f := - 1260;
        ELSIF x =- 1468 THEN
            tanh_f := - 1260;
        ELSIF x =- 1467 THEN
            tanh_f := - 1259;
        ELSIF x =- 1466 THEN
            tanh_f := - 1259;
        ELSIF x =- 1465 THEN
            tanh_f := - 1258;
        ELSIF x =- 1464 THEN
            tanh_f := - 1257;
        ELSIF x =- 1463 THEN
            tanh_f := - 1257;
        ELSIF x =- 1462 THEN
            tanh_f := - 1256;
        ELSIF x =- 1461 THEN
            tanh_f := - 1255;
        ELSIF x =- 1460 THEN
            tanh_f := - 1255;
        ELSIF x =- 1459 THEN
            tanh_f := - 1254;
        ELSIF x =- 1458 THEN
            tanh_f := - 1253;
        ELSIF x =- 1457 THEN
            tanh_f := - 1253;
        ELSIF x =- 1456 THEN
            tanh_f := - 1252;
        ELSIF x =- 1455 THEN
            tanh_f := - 1251;
        ELSIF x =- 1454 THEN
            tanh_f := - 1251;
        ELSIF x =- 1453 THEN
            tanh_f := - 1250;
        ELSIF x =- 1452 THEN
            tanh_f := - 1250;
        ELSIF x =- 1451 THEN
            tanh_f := - 1249;
        ELSIF x =- 1450 THEN
            tanh_f := - 1248;
        ELSIF x =- 1449 THEN
            tanh_f := - 1248;
        ELSIF x =- 1448 THEN
            tanh_f := - 1247;
        ELSIF x =- 1447 THEN
            tanh_f := - 1246;
        ELSIF x =- 1446 THEN
            tanh_f := - 1246;
        ELSIF x =- 1445 THEN
            tanh_f := - 1245;
        ELSIF x =- 1444 THEN
            tanh_f := - 1244;
        ELSIF x =- 1443 THEN
            tanh_f := - 1244;
        ELSIF x =- 1442 THEN
            tanh_f := - 1243;
        ELSIF x =- 1441 THEN
            tanh_f := - 1242;
        ELSIF x =- 1440 THEN
            tanh_f := - 1242;
        ELSIF x =- 1439 THEN
            tanh_f := - 1241;
        ELSIF x =- 1438 THEN
            tanh_f := - 1241;
        ELSIF x =- 1437 THEN
            tanh_f := - 1240;
        ELSIF x =- 1436 THEN
            tanh_f := - 1239;
        ELSIF x =- 1435 THEN
            tanh_f := - 1239;
        ELSIF x =- 1434 THEN
            tanh_f := - 1238;
        ELSIF x =- 1433 THEN
            tanh_f := - 1237;
        ELSIF x =- 1432 THEN
            tanh_f := - 1237;
        ELSIF x =- 1431 THEN
            tanh_f := - 1236;
        ELSIF x =- 1430 THEN
            tanh_f := - 1235;
        ELSIF x =- 1429 THEN
            tanh_f := - 1235;
        ELSIF x =- 1428 THEN
            tanh_f := - 1234;
        ELSIF x =- 1427 THEN
            tanh_f := - 1233;
        ELSIF x =- 1426 THEN
            tanh_f := - 1233;
        ELSIF x =- 1425 THEN
            tanh_f := - 1232;
        ELSIF x =- 1424 THEN
            tanh_f := - 1232;
        ELSIF x =- 1423 THEN
            tanh_f := - 1231;
        ELSIF x =- 1422 THEN
            tanh_f := - 1230;
        ELSIF x =- 1421 THEN
            tanh_f := - 1230;
        ELSIF x =- 1420 THEN
            tanh_f := - 1229;
        ELSIF x =- 1419 THEN
            tanh_f := - 1228;
        ELSIF x =- 1418 THEN
            tanh_f := - 1228;
        ELSIF x =- 1417 THEN
            tanh_f := - 1227;
        ELSIF x =- 1416 THEN
            tanh_f := - 1226;
        ELSIF x =- 1415 THEN
            tanh_f := - 1226;
        ELSIF x =- 1414 THEN
            tanh_f := - 1225;
        ELSIF x =- 1413 THEN
            tanh_f := - 1224;
        ELSIF x =- 1412 THEN
            tanh_f := - 1224;
        ELSIF x =- 1411 THEN
            tanh_f := - 1223;
        ELSIF x =- 1410 THEN
            tanh_f := - 1223;
        ELSIF x =- 1409 THEN
            tanh_f := - 1222;
        ELSIF x =- 1408 THEN
            tanh_f := - 1221;
        ELSIF x =- 1407 THEN
            tanh_f := - 1221;
        ELSIF x =- 1406 THEN
            tanh_f := - 1220;
        ELSIF x =- 1405 THEN
            tanh_f := - 1219;
        ELSIF x =- 1404 THEN
            tanh_f := - 1219;
        ELSIF x =- 1403 THEN
            tanh_f := - 1218;
        ELSIF x =- 1402 THEN
            tanh_f := - 1217;
        ELSIF x =- 1401 THEN
            tanh_f := - 1217;
        ELSIF x =- 1400 THEN
            tanh_f := - 1216;
        ELSIF x =- 1399 THEN
            tanh_f := - 1215;
        ELSIF x =- 1398 THEN
            tanh_f := - 1215;
        ELSIF x =- 1397 THEN
            tanh_f := - 1214;
        ELSIF x =- 1396 THEN
            tanh_f := - 1214;
        ELSIF x =- 1395 THEN
            tanh_f := - 1213;
        ELSIF x =- 1394 THEN
            tanh_f := - 1212;
        ELSIF x =- 1393 THEN
            tanh_f := - 1212;
        ELSIF x =- 1392 THEN
            tanh_f := - 1211;
        ELSIF x =- 1391 THEN
            tanh_f := - 1210;
        ELSIF x =- 1390 THEN
            tanh_f := - 1210;
        ELSIF x =- 1389 THEN
            tanh_f := - 1209;
        ELSIF x =- 1388 THEN
            tanh_f := - 1208;
        ELSIF x =- 1387 THEN
            tanh_f := - 1208;
        ELSIF x =- 1386 THEN
            tanh_f := - 1207;
        ELSIF x =- 1385 THEN
            tanh_f := - 1206;
        ELSIF x =- 1384 THEN
            tanh_f := - 1206;
        ELSIF x =- 1383 THEN
            tanh_f := - 1205;
        ELSIF x =- 1382 THEN
            tanh_f := - 1205;
        ELSIF x =- 1381 THEN
            tanh_f := - 1204;
        ELSIF x =- 1380 THEN
            tanh_f := - 1203;
        ELSIF x =- 1379 THEN
            tanh_f := - 1203;
        ELSIF x =- 1378 THEN
            tanh_f := - 1202;
        ELSIF x =- 1377 THEN
            tanh_f := - 1201;
        ELSIF x =- 1376 THEN
            tanh_f := - 1201;
        ELSIF x =- 1375 THEN
            tanh_f := - 1200;
        ELSIF x =- 1374 THEN
            tanh_f := - 1199;
        ELSIF x =- 1373 THEN
            tanh_f := - 1199;
        ELSIF x =- 1372 THEN
            tanh_f := - 1198;
        ELSIF x =- 1371 THEN
            tanh_f := - 1197;
        ELSIF x =- 1370 THEN
            tanh_f := - 1197;
        ELSIF x =- 1369 THEN
            tanh_f := - 1196;
        ELSIF x =- 1368 THEN
            tanh_f := - 1196;
        ELSIF x =- 1367 THEN
            tanh_f := - 1195;
        ELSIF x =- 1366 THEN
            tanh_f := - 1194;
        ELSIF x =- 1365 THEN
            tanh_f := - 1194;
        ELSIF x =- 1364 THEN
            tanh_f := - 1193;
        ELSIF x =- 1363 THEN
            tanh_f := - 1192;
        ELSIF x =- 1362 THEN
            tanh_f := - 1192;
        ELSIF x =- 1361 THEN
            tanh_f := - 1191;
        ELSIF x =- 1360 THEN
            tanh_f := - 1190;
        ELSIF x =- 1359 THEN
            tanh_f := - 1190;
        ELSIF x =- 1358 THEN
            tanh_f := - 1189;
        ELSIF x =- 1357 THEN
            tanh_f := - 1188;
        ELSIF x =- 1356 THEN
            tanh_f := - 1188;
        ELSIF x =- 1355 THEN
            tanh_f := - 1187;
        ELSIF x =- 1354 THEN
            tanh_f := - 1187;
        ELSIF x =- 1353 THEN
            tanh_f := - 1186;
        ELSIF x =- 1352 THEN
            tanh_f := - 1185;
        ELSIF x =- 1351 THEN
            tanh_f := - 1185;
        ELSIF x =- 1350 THEN
            tanh_f := - 1184;
        ELSIF x =- 1349 THEN
            tanh_f := - 1183;
        ELSIF x =- 1348 THEN
            tanh_f := - 1183;
        ELSIF x =- 1347 THEN
            tanh_f := - 1182;
        ELSIF x =- 1346 THEN
            tanh_f := - 1181;
        ELSIF x =- 1345 THEN
            tanh_f := - 1181;
        ELSIF x =- 1344 THEN
            tanh_f := - 1180;
        ELSIF x =- 1343 THEN
            tanh_f := - 1179;
        ELSIF x =- 1342 THEN
            tanh_f := - 1179;
        ELSIF x =- 1341 THEN
            tanh_f := - 1178;
        ELSIF x =- 1340 THEN
            tanh_f := - 1178;
        ELSIF x =- 1339 THEN
            tanh_f := - 1177;
        ELSIF x =- 1338 THEN
            tanh_f := - 1176;
        ELSIF x =- 1337 THEN
            tanh_f := - 1176;
        ELSIF x =- 1336 THEN
            tanh_f := - 1175;
        ELSIF x =- 1335 THEN
            tanh_f := - 1174;
        ELSIF x =- 1334 THEN
            tanh_f := - 1174;
        ELSIF x =- 1333 THEN
            tanh_f := - 1173;
        ELSIF x =- 1332 THEN
            tanh_f := - 1172;
        ELSIF x =- 1331 THEN
            tanh_f := - 1172;
        ELSIF x =- 1330 THEN
            tanh_f := - 1171;
        ELSIF x =- 1329 THEN
            tanh_f := - 1170;
        ELSIF x =- 1328 THEN
            tanh_f := - 1170;
        ELSIF x =- 1327 THEN
            tanh_f := - 1169;
        ELSIF x =- 1326 THEN
            tanh_f := - 1169;
        ELSIF x =- 1325 THEN
            tanh_f := - 1168;
        ELSIF x =- 1324 THEN
            tanh_f := - 1167;
        ELSIF x =- 1323 THEN
            tanh_f := - 1167;
        ELSIF x =- 1322 THEN
            tanh_f := - 1166;
        ELSIF x =- 1321 THEN
            tanh_f := - 1165;
        ELSIF x =- 1320 THEN
            tanh_f := - 1165;
        ELSIF x =- 1319 THEN
            tanh_f := - 1164;
        ELSIF x =- 1318 THEN
            tanh_f := - 1163;
        ELSIF x =- 1317 THEN
            tanh_f := - 1163;
        ELSIF x =- 1316 THEN
            tanh_f := - 1162;
        ELSIF x =- 1315 THEN
            tanh_f := - 1161;
        ELSIF x =- 1314 THEN
            tanh_f := - 1161;
        ELSIF x =- 1313 THEN
            tanh_f := - 1160;
        ELSIF x =- 1312 THEN
            tanh_f := - 1160;
        ELSIF x =- 1311 THEN
            tanh_f := - 1159;
        ELSIF x =- 1310 THEN
            tanh_f := - 1158;
        ELSIF x =- 1309 THEN
            tanh_f := - 1158;
        ELSIF x =- 1308 THEN
            tanh_f := - 1157;
        ELSIF x =- 1307 THEN
            tanh_f := - 1156;
        ELSIF x =- 1306 THEN
            tanh_f := - 1156;
        ELSIF x =- 1305 THEN
            tanh_f := - 1155;
        ELSIF x =- 1304 THEN
            tanh_f := - 1154;
        ELSIF x =- 1303 THEN
            tanh_f := - 1154;
        ELSIF x =- 1302 THEN
            tanh_f := - 1153;
        ELSIF x =- 1301 THEN
            tanh_f := - 1152;
        ELSIF x =- 1300 THEN
            tanh_f := - 1152;
        ELSIF x =- 1299 THEN
            tanh_f := - 1151;
        ELSIF x =- 1298 THEN
            tanh_f := - 1151;
        ELSIF x =- 1297 THEN
            tanh_f := - 1150;
        ELSIF x =- 1296 THEN
            tanh_f := - 1149;
        ELSIF x =- 1295 THEN
            tanh_f := - 1149;
        ELSIF x =- 1294 THEN
            tanh_f := - 1148;
        ELSIF x =- 1293 THEN
            tanh_f := - 1147;
        ELSIF x =- 1292 THEN
            tanh_f := - 1147;
        ELSIF x =- 1291 THEN
            tanh_f := - 1146;
        ELSIF x =- 1290 THEN
            tanh_f := - 1145;
        ELSIF x =- 1289 THEN
            tanh_f := - 1145;
        ELSIF x =- 1288 THEN
            tanh_f := - 1144;
        ELSIF x =- 1287 THEN
            tanh_f := - 1143;
        ELSIF x =- 1286 THEN
            tanh_f := - 1143;
        ELSIF x =- 1285 THEN
            tanh_f := - 1142;
        ELSIF x =- 1284 THEN
            tanh_f := - 1142;
        ELSIF x =- 1283 THEN
            tanh_f := - 1141;
        ELSIF x =- 1282 THEN
            tanh_f := - 1140;
        ELSIF x =- 1281 THEN
            tanh_f := - 1140;
        ELSIF x =- 1280 THEN
            tanh_f := - 1139;
        ELSIF x =- 1279 THEN
            tanh_f := - 1138;
        ELSIF x =- 1278 THEN
            tanh_f := - 1138;
        ELSIF x =- 1277 THEN
            tanh_f := - 1137;
        ELSIF x =- 1276 THEN
            tanh_f := - 1136;
        ELSIF x =- 1275 THEN
            tanh_f := - 1135;
        ELSIF x =- 1274 THEN
            tanh_f := - 1135;
        ELSIF x =- 1273 THEN
            tanh_f := - 1134;
        ELSIF x =- 1272 THEN
            tanh_f := - 1133;
        ELSIF x =- 1271 THEN
            tanh_f := - 1132;
        ELSIF x =- 1270 THEN
            tanh_f := - 1132;
        ELSIF x =- 1269 THEN
            tanh_f := - 1131;
        ELSIF x =- 1268 THEN
            tanh_f := - 1130;
        ELSIF x =- 1267 THEN
            tanh_f := - 1129;
        ELSIF x =- 1266 THEN
            tanh_f := - 1129;
        ELSIF x =- 1265 THEN
            tanh_f := - 1128;
        ELSIF x =- 1264 THEN
            tanh_f := - 1127;
        ELSIF x =- 1263 THEN
            tanh_f := - 1126;
        ELSIF x =- 1262 THEN
            tanh_f := - 1126;
        ELSIF x =- 1261 THEN
            tanh_f := - 1125;
        ELSIF x =- 1260 THEN
            tanh_f := - 1124;
        ELSIF x =- 1259 THEN
            tanh_f := - 1123;
        ELSIF x =- 1258 THEN
            tanh_f := - 1123;
        ELSIF x =- 1257 THEN
            tanh_f := - 1122;
        ELSIF x =- 1256 THEN
            tanh_f := - 1121;
        ELSIF x =- 1255 THEN
            tanh_f := - 1120;
        ELSIF x =- 1254 THEN
            tanh_f := - 1120;
        ELSIF x =- 1253 THEN
            tanh_f := - 1119;
        ELSIF x =- 1252 THEN
            tanh_f := - 1118;
        ELSIF x =- 1251 THEN
            tanh_f := - 1117;
        ELSIF x =- 1250 THEN
            tanh_f := - 1117;
        ELSIF x =- 1249 THEN
            tanh_f := - 1116;
        ELSIF x =- 1248 THEN
            tanh_f := - 1115;
        ELSIF x =- 1247 THEN
            tanh_f := - 1114;
        ELSIF x =- 1246 THEN
            tanh_f := - 1114;
        ELSIF x =- 1245 THEN
            tanh_f := - 1113;
        ELSIF x =- 1244 THEN
            tanh_f := - 1112;
        ELSIF x =- 1243 THEN
            tanh_f := - 1111;
        ELSIF x =- 1242 THEN
            tanh_f := - 1111;
        ELSIF x =- 1241 THEN
            tanh_f := - 1110;
        ELSIF x =- 1240 THEN
            tanh_f := - 1109;
        ELSIF x =- 1239 THEN
            tanh_f := - 1108;
        ELSIF x =- 1238 THEN
            tanh_f := - 1108;
        ELSIF x =- 1237 THEN
            tanh_f := - 1107;
        ELSIF x =- 1236 THEN
            tanh_f := - 1106;
        ELSIF x =- 1235 THEN
            tanh_f := - 1106;
        ELSIF x =- 1234 THEN
            tanh_f := - 1105;
        ELSIF x =- 1233 THEN
            tanh_f := - 1104;
        ELSIF x =- 1232 THEN
            tanh_f := - 1103;
        ELSIF x =- 1231 THEN
            tanh_f := - 1103;
        ELSIF x =- 1230 THEN
            tanh_f := - 1102;
        ELSIF x =- 1229 THEN
            tanh_f := - 1101;
        ELSIF x =- 1228 THEN
            tanh_f := - 1100;
        ELSIF x =- 1227 THEN
            tanh_f := - 1100;
        ELSIF x =- 1226 THEN
            tanh_f := - 1099;
        ELSIF x =- 1225 THEN
            tanh_f := - 1098;
        ELSIF x =- 1224 THEN
            tanh_f := - 1097;
        ELSIF x =- 1223 THEN
            tanh_f := - 1097;
        ELSIF x =- 1222 THEN
            tanh_f := - 1096;
        ELSIF x =- 1221 THEN
            tanh_f := - 1095;
        ELSIF x =- 1220 THEN
            tanh_f := - 1094;
        ELSIF x =- 1219 THEN
            tanh_f := - 1094;
        ELSIF x =- 1218 THEN
            tanh_f := - 1093;
        ELSIF x =- 1217 THEN
            tanh_f := - 1092;
        ELSIF x =- 1216 THEN
            tanh_f := - 1091;
        ELSIF x =- 1215 THEN
            tanh_f := - 1091;
        ELSIF x =- 1214 THEN
            tanh_f := - 1090;
        ELSIF x =- 1213 THEN
            tanh_f := - 1089;
        ELSIF x =- 1212 THEN
            tanh_f := - 1088;
        ELSIF x =- 1211 THEN
            tanh_f := - 1088;
        ELSIF x =- 1210 THEN
            tanh_f := - 1087;
        ELSIF x =- 1209 THEN
            tanh_f := - 1086;
        ELSIF x =- 1208 THEN
            tanh_f := - 1085;
        ELSIF x =- 1207 THEN
            tanh_f := - 1085;
        ELSIF x =- 1206 THEN
            tanh_f := - 1084;
        ELSIF x =- 1205 THEN
            tanh_f := - 1083;
        ELSIF x =- 1204 THEN
            tanh_f := - 1082;
        ELSIF x =- 1203 THEN
            tanh_f := - 1082;
        ELSIF x =- 1202 THEN
            tanh_f := - 1081;
        ELSIF x =- 1201 THEN
            tanh_f := - 1080;
        ELSIF x =- 1200 THEN
            tanh_f := - 1079;
        ELSIF x =- 1199 THEN
            tanh_f := - 1079;
        ELSIF x =- 1198 THEN
            tanh_f := - 1078;
        ELSIF x =- 1197 THEN
            tanh_f := - 1077;
        ELSIF x =- 1196 THEN
            tanh_f := - 1076;
        ELSIF x =- 1195 THEN
            tanh_f := - 1076;
        ELSIF x =- 1194 THEN
            tanh_f := - 1075;
        ELSIF x =- 1193 THEN
            tanh_f := - 1074;
        ELSIF x =- 1192 THEN
            tanh_f := - 1074;
        ELSIF x =- 1191 THEN
            tanh_f := - 1073;
        ELSIF x =- 1190 THEN
            tanh_f := - 1072;
        ELSIF x =- 1189 THEN
            tanh_f := - 1071;
        ELSIF x =- 1188 THEN
            tanh_f := - 1071;
        ELSIF x =- 1187 THEN
            tanh_f := - 1070;
        ELSIF x =- 1186 THEN
            tanh_f := - 1069;
        ELSIF x =- 1185 THEN
            tanh_f := - 1068;
        ELSIF x =- 1184 THEN
            tanh_f := - 1068;
        ELSIF x =- 1183 THEN
            tanh_f := - 1067;
        ELSIF x =- 1182 THEN
            tanh_f := - 1066;
        ELSIF x =- 1181 THEN
            tanh_f := - 1065;
        ELSIF x =- 1180 THEN
            tanh_f := - 1065;
        ELSIF x =- 1179 THEN
            tanh_f := - 1064;
        ELSIF x =- 1178 THEN
            tanh_f := - 1063;
        ELSIF x =- 1177 THEN
            tanh_f := - 1062;
        ELSIF x =- 1176 THEN
            tanh_f := - 1062;
        ELSIF x =- 1175 THEN
            tanh_f := - 1061;
        ELSIF x =- 1174 THEN
            tanh_f := - 1060;
        ELSIF x =- 1173 THEN
            tanh_f := - 1059;
        ELSIF x =- 1172 THEN
            tanh_f := - 1059;
        ELSIF x =- 1171 THEN
            tanh_f := - 1058;
        ELSIF x =- 1170 THEN
            tanh_f := - 1057;
        ELSIF x =- 1169 THEN
            tanh_f := - 1056;
        ELSIF x =- 1168 THEN
            tanh_f := - 1056;
        ELSIF x =- 1167 THEN
            tanh_f := - 1055;
        ELSIF x =- 1166 THEN
            tanh_f := - 1054;
        ELSIF x =- 1165 THEN
            tanh_f := - 1053;
        ELSIF x =- 1164 THEN
            tanh_f := - 1053;
        ELSIF x =- 1163 THEN
            tanh_f := - 1052;
        ELSIF x =- 1162 THEN
            tanh_f := - 1051;
        ELSIF x =- 1161 THEN
            tanh_f := - 1050;
        ELSIF x =- 1160 THEN
            tanh_f := - 1050;
        ELSIF x =- 1159 THEN
            tanh_f := - 1049;
        ELSIF x =- 1158 THEN
            tanh_f := - 1048;
        ELSIF x =- 1157 THEN
            tanh_f := - 1047;
        ELSIF x =- 1156 THEN
            tanh_f := - 1047;
        ELSIF x =- 1155 THEN
            tanh_f := - 1046;
        ELSIF x =- 1154 THEN
            tanh_f := - 1045;
        ELSIF x =- 1153 THEN
            tanh_f := - 1044;
        ELSIF x =- 1152 THEN
            tanh_f := - 1044;
        ELSIF x =- 1151 THEN
            tanh_f := - 1043;
        ELSIF x =- 1150 THEN
            tanh_f := - 1042;
        ELSIF x =- 1149 THEN
            tanh_f := - 1042;
        ELSIF x =- 1148 THEN
            tanh_f := - 1041;
        ELSIF x =- 1147 THEN
            tanh_f := - 1040;
        ELSIF x =- 1146 THEN
            tanh_f := - 1039;
        ELSIF x =- 1145 THEN
            tanh_f := - 1039;
        ELSIF x =- 1144 THEN
            tanh_f := - 1038;
        ELSIF x =- 1143 THEN
            tanh_f := - 1037;
        ELSIF x =- 1142 THEN
            tanh_f := - 1036;
        ELSIF x =- 1141 THEN
            tanh_f := - 1036;
        ELSIF x =- 1140 THEN
            tanh_f := - 1035;
        ELSIF x =- 1139 THEN
            tanh_f := - 1034;
        ELSIF x =- 1138 THEN
            tanh_f := - 1033;
        ELSIF x =- 1137 THEN
            tanh_f := - 1033;
        ELSIF x =- 1136 THEN
            tanh_f := - 1032;
        ELSIF x =- 1135 THEN
            tanh_f := - 1031;
        ELSIF x =- 1134 THEN
            tanh_f := - 1030;
        ELSIF x =- 1133 THEN
            tanh_f := - 1030;
        ELSIF x =- 1132 THEN
            tanh_f := - 1029;
        ELSIF x =- 1131 THEN
            tanh_f := - 1028;
        ELSIF x =- 1130 THEN
            tanh_f := - 1027;
        ELSIF x =- 1129 THEN
            tanh_f := - 1027;
        ELSIF x =- 1128 THEN
            tanh_f := - 1026;
        ELSIF x =- 1127 THEN
            tanh_f := - 1025;
        ELSIF x =- 1126 THEN
            tanh_f := - 1024;
        ELSIF x =- 1125 THEN
            tanh_f := - 1024;
        ELSIF x =- 1124 THEN
            tanh_f := - 1023;
        ELSIF x =- 1123 THEN
            tanh_f := - 1022;
        ELSIF x =- 1122 THEN
            tanh_f := - 1021;
        ELSIF x =- 1121 THEN
            tanh_f := - 1021;
        ELSIF x =- 1120 THEN
            tanh_f := - 1020;
        ELSIF x =- 1119 THEN
            tanh_f := - 1019;
        ELSIF x =- 1118 THEN
            tanh_f := - 1018;
        ELSIF x =- 1117 THEN
            tanh_f := - 1018;
        ELSIF x =- 1116 THEN
            tanh_f := - 1017;
        ELSIF x =- 1115 THEN
            tanh_f := - 1016;
        ELSIF x =- 1114 THEN
            tanh_f := - 1015;
        ELSIF x =- 1113 THEN
            tanh_f := - 1015;
        ELSIF x =- 1112 THEN
            tanh_f := - 1014;
        ELSIF x =- 1111 THEN
            tanh_f := - 1013;
        ELSIF x =- 1110 THEN
            tanh_f := - 1012;
        ELSIF x =- 1109 THEN
            tanh_f := - 1012;
        ELSIF x =- 1108 THEN
            tanh_f := - 1011;
        ELSIF x =- 1107 THEN
            tanh_f := - 1010;
        ELSIF x =- 1106 THEN
            tanh_f := - 1010;
        ELSIF x =- 1105 THEN
            tanh_f := - 1009;
        ELSIF x =- 1104 THEN
            tanh_f := - 1008;
        ELSIF x =- 1103 THEN
            tanh_f := - 1007;
        ELSIF x =- 1102 THEN
            tanh_f := - 1007;
        ELSIF x =- 1101 THEN
            tanh_f := - 1006;
        ELSIF x =- 1100 THEN
            tanh_f := - 1005;
        ELSIF x =- 1099 THEN
            tanh_f := - 1004;
        ELSIF x =- 1098 THEN
            tanh_f := - 1004;
        ELSIF x =- 1097 THEN
            tanh_f := - 1003;
        ELSIF x =- 1096 THEN
            tanh_f := - 1002;
        ELSIF x =- 1095 THEN
            tanh_f := - 1001;
        ELSIF x =- 1094 THEN
            tanh_f := - 1001;
        ELSIF x =- 1093 THEN
            tanh_f := - 1000;
        ELSIF x =- 1092 THEN
            tanh_f := - 999;
        ELSIF x =- 1091 THEN
            tanh_f := - 998;
        ELSIF x =- 1090 THEN
            tanh_f := - 998;
        ELSIF x =- 1089 THEN
            tanh_f := - 997;
        ELSIF x =- 1088 THEN
            tanh_f := - 996;
        ELSIF x =- 1087 THEN
            tanh_f := - 995;
        ELSIF x =- 1086 THEN
            tanh_f := - 995;
        ELSIF x =- 1085 THEN
            tanh_f := - 994;
        ELSIF x =- 1084 THEN
            tanh_f := - 993;
        ELSIF x =- 1083 THEN
            tanh_f := - 992;
        ELSIF x =- 1082 THEN
            tanh_f := - 992;
        ELSIF x =- 1081 THEN
            tanh_f := - 991;
        ELSIF x =- 1080 THEN
            tanh_f := - 990;
        ELSIF x =- 1079 THEN
            tanh_f := - 989;
        ELSIF x =- 1078 THEN
            tanh_f := - 989;
        ELSIF x =- 1077 THEN
            tanh_f := - 988;
        ELSIF x =- 1076 THEN
            tanh_f := - 987;
        ELSIF x =- 1075 THEN
            tanh_f := - 986;
        ELSIF x =- 1074 THEN
            tanh_f := - 986;
        ELSIF x =- 1073 THEN
            tanh_f := - 985;
        ELSIF x =- 1072 THEN
            tanh_f := - 984;
        ELSIF x =- 1071 THEN
            tanh_f := - 983;
        ELSIF x =- 1070 THEN
            tanh_f := - 983;
        ELSIF x =- 1069 THEN
            tanh_f := - 982;
        ELSIF x =- 1068 THEN
            tanh_f := - 981;
        ELSIF x =- 1067 THEN
            tanh_f := - 980;
        ELSIF x =- 1066 THEN
            tanh_f := - 980;
        ELSIF x =- 1065 THEN
            tanh_f := - 979;
        ELSIF x =- 1064 THEN
            tanh_f := - 978;
        ELSIF x =- 1063 THEN
            tanh_f := - 978;
        ELSIF x =- 1062 THEN
            tanh_f := - 977;
        ELSIF x =- 1061 THEN
            tanh_f := - 976;
        ELSIF x =- 1060 THEN
            tanh_f := - 975;
        ELSIF x =- 1059 THEN
            tanh_f := - 975;
        ELSIF x =- 1058 THEN
            tanh_f := - 974;
        ELSIF x =- 1057 THEN
            tanh_f := - 973;
        ELSIF x =- 1056 THEN
            tanh_f := - 972;
        ELSIF x =- 1055 THEN
            tanh_f := - 972;
        ELSIF x =- 1054 THEN
            tanh_f := - 971;
        ELSIF x =- 1053 THEN
            tanh_f := - 970;
        ELSIF x =- 1052 THEN
            tanh_f := - 969;
        ELSIF x =- 1051 THEN
            tanh_f := - 969;
        ELSIF x =- 1050 THEN
            tanh_f := - 968;
        ELSIF x =- 1049 THEN
            tanh_f := - 967;
        ELSIF x =- 1048 THEN
            tanh_f := - 966;
        ELSIF x =- 1047 THEN
            tanh_f := - 966;
        ELSIF x =- 1046 THEN
            tanh_f := - 965;
        ELSIF x =- 1045 THEN
            tanh_f := - 964;
        ELSIF x =- 1044 THEN
            tanh_f := - 963;
        ELSIF x =- 1043 THEN
            tanh_f := - 963;
        ELSIF x =- 1042 THEN
            tanh_f := - 962;
        ELSIF x =- 1041 THEN
            tanh_f := - 961;
        ELSIF x =- 1040 THEN
            tanh_f := - 960;
        ELSIF x =- 1039 THEN
            tanh_f := - 960;
        ELSIF x =- 1038 THEN
            tanh_f := - 959;
        ELSIF x =- 1037 THEN
            tanh_f := - 958;
        ELSIF x =- 1036 THEN
            tanh_f := - 957;
        ELSIF x =- 1035 THEN
            tanh_f := - 957;
        ELSIF x =- 1034 THEN
            tanh_f := - 956;
        ELSIF x =- 1033 THEN
            tanh_f := - 955;
        ELSIF x =- 1032 THEN
            tanh_f := - 954;
        ELSIF x =- 1031 THEN
            tanh_f := - 954;
        ELSIF x =- 1030 THEN
            tanh_f := - 953;
        ELSIF x =- 1029 THEN
            tanh_f := - 952;
        ELSIF x =- 1028 THEN
            tanh_f := - 951;
        ELSIF x =- 1027 THEN
            tanh_f := - 951;
        ELSIF x =- 1026 THEN
            tanh_f := - 950;
        ELSIF x =- 1025 THEN
            tanh_f := - 949;
        ELSIF x =- 1024 THEN
            tanh_f := - 948;
        ELSIF x =- 1023 THEN
            tanh_f := - 948;
        ELSIF x =- 1022 THEN
            tanh_f := - 947;
        ELSIF x =- 1021 THEN
            tanh_f := - 946;
        ELSIF x =- 1020 THEN
            tanh_f := - 945;
        ELSIF x =- 1019 THEN
            tanh_f := - 944;
        ELSIF x =- 1018 THEN
            tanh_f := - 944;
        ELSIF x =- 1017 THEN
            tanh_f := - 943;
        ELSIF x =- 1016 THEN
            tanh_f := - 942;
        ELSIF x =- 1015 THEN
            tanh_f := - 941;
        ELSIF x =- 1014 THEN
            tanh_f := - 940;
        ELSIF x =- 1013 THEN
            tanh_f := - 939;
        ELSIF x =- 1012 THEN
            tanh_f := - 939;
        ELSIF x =- 1011 THEN
            tanh_f := - 938;
        ELSIF x =- 1010 THEN
            tanh_f := - 937;
        ELSIF x =- 1009 THEN
            tanh_f := - 936;
        ELSIF x =- 1008 THEN
            tanh_f := - 935;
        ELSIF x =- 1007 THEN
            tanh_f := - 934;
        ELSIF x =- 1006 THEN
            tanh_f := - 934;
        ELSIF x =- 1005 THEN
            tanh_f := - 933;
        ELSIF x =- 1004 THEN
            tanh_f := - 932;
        ELSIF x =- 1003 THEN
            tanh_f := - 931;
        ELSIF x =- 1002 THEN
            tanh_f := - 930;
        ELSIF x =- 1001 THEN
            tanh_f := - 929;
        ELSIF x =- 1000 THEN
            tanh_f := - 929;
        ELSIF x =- 999 THEN
            tanh_f := - 928;
        ELSIF x =- 998 THEN
            tanh_f := - 927;
        ELSIF x =- 997 THEN
            tanh_f := - 926;
        ELSIF x =- 996 THEN
            tanh_f := - 925;
        ELSIF x =- 995 THEN
            tanh_f := - 924;
        ELSIF x =- 994 THEN
            tanh_f := - 924;
        ELSIF x =- 993 THEN
            tanh_f := - 923;
        ELSIF x =- 992 THEN
            tanh_f := - 922;
        ELSIF x =- 991 THEN
            tanh_f := - 921;
        ELSIF x =- 990 THEN
            tanh_f := - 920;
        ELSIF x =- 989 THEN
            tanh_f := - 920;
        ELSIF x =- 988 THEN
            tanh_f := - 919;
        ELSIF x =- 987 THEN
            tanh_f := - 918;
        ELSIF x =- 986 THEN
            tanh_f := - 917;
        ELSIF x =- 985 THEN
            tanh_f := - 916;
        ELSIF x =- 984 THEN
            tanh_f := - 915;
        ELSIF x =- 983 THEN
            tanh_f := - 915;
        ELSIF x =- 982 THEN
            tanh_f := - 914;
        ELSIF x =- 981 THEN
            tanh_f := - 913;
        ELSIF x =- 980 THEN
            tanh_f := - 912;
        ELSIF x =- 979 THEN
            tanh_f := - 911;
        ELSIF x =- 978 THEN
            tanh_f := - 910;
        ELSIF x =- 977 THEN
            tanh_f := - 910;
        ELSIF x =- 976 THEN
            tanh_f := - 909;
        ELSIF x =- 975 THEN
            tanh_f := - 908;
        ELSIF x =- 974 THEN
            tanh_f := - 907;
        ELSIF x =- 973 THEN
            tanh_f := - 906;
        ELSIF x =- 972 THEN
            tanh_f := - 905;
        ELSIF x =- 971 THEN
            tanh_f := - 905;
        ELSIF x =- 970 THEN
            tanh_f := - 904;
        ELSIF x =- 969 THEN
            tanh_f := - 903;
        ELSIF x =- 968 THEN
            tanh_f := - 902;
        ELSIF x =- 967 THEN
            tanh_f := - 901;
        ELSIF x =- 966 THEN
            tanh_f := - 900;
        ELSIF x =- 965 THEN
            tanh_f := - 900;
        ELSIF x =- 964 THEN
            tanh_f := - 899;
        ELSIF x =- 963 THEN
            tanh_f := - 898;
        ELSIF x =- 962 THEN
            tanh_f := - 897;
        ELSIF x =- 961 THEN
            tanh_f := - 896;
        ELSIF x =- 960 THEN
            tanh_f := - 895;
        ELSIF x =- 959 THEN
            tanh_f := - 895;
        ELSIF x =- 958 THEN
            tanh_f := - 894;
        ELSIF x =- 957 THEN
            tanh_f := - 893;
        ELSIF x =- 956 THEN
            tanh_f := - 892;
        ELSIF x =- 955 THEN
            tanh_f := - 891;
        ELSIF x =- 954 THEN
            tanh_f := - 891;
        ELSIF x =- 953 THEN
            tanh_f := - 890;
        ELSIF x =- 952 THEN
            tanh_f := - 889;
        ELSIF x =- 951 THEN
            tanh_f := - 888;
        ELSIF x =- 950 THEN
            tanh_f := - 887;
        ELSIF x =- 949 THEN
            tanh_f := - 886;
        ELSIF x =- 948 THEN
            tanh_f := - 886;
        ELSIF x =- 947 THEN
            tanh_f := - 885;
        ELSIF x =- 946 THEN
            tanh_f := - 884;
        ELSIF x =- 945 THEN
            tanh_f := - 883;
        ELSIF x =- 944 THEN
            tanh_f := - 882;
        ELSIF x =- 943 THEN
            tanh_f := - 881;
        ELSIF x =- 942 THEN
            tanh_f := - 881;
        ELSIF x =- 941 THEN
            tanh_f := - 880;
        ELSIF x =- 940 THEN
            tanh_f := - 879;
        ELSIF x =- 939 THEN
            tanh_f := - 878;
        ELSIF x =- 938 THEN
            tanh_f := - 877;
        ELSIF x =- 937 THEN
            tanh_f := - 876;
        ELSIF x =- 936 THEN
            tanh_f := - 876;
        ELSIF x =- 935 THEN
            tanh_f := - 875;
        ELSIF x =- 934 THEN
            tanh_f := - 874;
        ELSIF x =- 933 THEN
            tanh_f := - 873;
        ELSIF x =- 932 THEN
            tanh_f := - 872;
        ELSIF x =- 931 THEN
            tanh_f := - 871;
        ELSIF x =- 930 THEN
            tanh_f := - 871;
        ELSIF x =- 929 THEN
            tanh_f := - 870;
        ELSIF x =- 928 THEN
            tanh_f := - 869;
        ELSIF x =- 927 THEN
            tanh_f := - 868;
        ELSIF x =- 926 THEN
            tanh_f := - 867;
        ELSIF x =- 925 THEN
            tanh_f := - 867;
        ELSIF x =- 924 THEN
            tanh_f := - 866;
        ELSIF x =- 923 THEN
            tanh_f := - 865;
        ELSIF x =- 922 THEN
            tanh_f := - 864;
        ELSIF x =- 921 THEN
            tanh_f := - 863;
        ELSIF x =- 920 THEN
            tanh_f := - 862;
        ELSIF x =- 919 THEN
            tanh_f := - 862;
        ELSIF x =- 918 THEN
            tanh_f := - 861;
        ELSIF x =- 917 THEN
            tanh_f := - 860;
        ELSIF x =- 916 THEN
            tanh_f := - 859;
        ELSIF x =- 915 THEN
            tanh_f := - 858;
        ELSIF x =- 914 THEN
            tanh_f := - 857;
        ELSIF x =- 913 THEN
            tanh_f := - 857;
        ELSIF x =- 912 THEN
            tanh_f := - 856;
        ELSIF x =- 911 THEN
            tanh_f := - 855;
        ELSIF x =- 910 THEN
            tanh_f := - 854;
        ELSIF x =- 909 THEN
            tanh_f := - 853;
        ELSIF x =- 908 THEN
            tanh_f := - 852;
        ELSIF x =- 907 THEN
            tanh_f := - 852;
        ELSIF x =- 906 THEN
            tanh_f := - 851;
        ELSIF x =- 905 THEN
            tanh_f := - 850;
        ELSIF x =- 904 THEN
            tanh_f := - 849;
        ELSIF x =- 903 THEN
            tanh_f := - 848;
        ELSIF x =- 902 THEN
            tanh_f := - 847;
        ELSIF x =- 901 THEN
            tanh_f := - 847;
        ELSIF x =- 900 THEN
            tanh_f := - 846;
        ELSIF x =- 899 THEN
            tanh_f := - 845;
        ELSIF x =- 898 THEN
            tanh_f := - 844;
        ELSIF x =- 897 THEN
            tanh_f := - 843;
        ELSIF x =- 896 THEN
            tanh_f := - 842;
        ELSIF x =- 895 THEN
            tanh_f := - 842;
        ELSIF x =- 894 THEN
            tanh_f := - 841;
        ELSIF x =- 893 THEN
            tanh_f := - 840;
        ELSIF x =- 892 THEN
            tanh_f := - 839;
        ELSIF x =- 891 THEN
            tanh_f := - 838;
        ELSIF x =- 890 THEN
            tanh_f := - 838;
        ELSIF x =- 889 THEN
            tanh_f := - 837;
        ELSIF x =- 888 THEN
            tanh_f := - 836;
        ELSIF x =- 887 THEN
            tanh_f := - 835;
        ELSIF x =- 886 THEN
            tanh_f := - 834;
        ELSIF x =- 885 THEN
            tanh_f := - 833;
        ELSIF x =- 884 THEN
            tanh_f := - 833;
        ELSIF x =- 883 THEN
            tanh_f := - 832;
        ELSIF x =- 882 THEN
            tanh_f := - 831;
        ELSIF x =- 881 THEN
            tanh_f := - 830;
        ELSIF x =- 880 THEN
            tanh_f := - 829;
        ELSIF x =- 879 THEN
            tanh_f := - 828;
        ELSIF x =- 878 THEN
            tanh_f := - 828;
        ELSIF x =- 877 THEN
            tanh_f := - 827;
        ELSIF x =- 876 THEN
            tanh_f := - 826;
        ELSIF x =- 875 THEN
            tanh_f := - 825;
        ELSIF x =- 874 THEN
            tanh_f := - 824;
        ELSIF x =- 873 THEN
            tanh_f := - 823;
        ELSIF x =- 872 THEN
            tanh_f := - 823;
        ELSIF x =- 871 THEN
            tanh_f := - 822;
        ELSIF x =- 870 THEN
            tanh_f := - 821;
        ELSIF x =- 869 THEN
            tanh_f := - 820;
        ELSIF x =- 868 THEN
            tanh_f := - 819;
        ELSIF x =- 867 THEN
            tanh_f := - 818;
        ELSIF x =- 866 THEN
            tanh_f := - 818;
        ELSIF x =- 865 THEN
            tanh_f := - 817;
        ELSIF x =- 864 THEN
            tanh_f := - 816;
        ELSIF x =- 863 THEN
            tanh_f := - 815;
        ELSIF x =- 862 THEN
            tanh_f := - 814;
        ELSIF x =- 861 THEN
            tanh_f := - 814;
        ELSIF x =- 860 THEN
            tanh_f := - 813;
        ELSIF x =- 859 THEN
            tanh_f := - 812;
        ELSIF x =- 858 THEN
            tanh_f := - 811;
        ELSIF x =- 857 THEN
            tanh_f := - 810;
        ELSIF x =- 856 THEN
            tanh_f := - 809;
        ELSIF x =- 855 THEN
            tanh_f := - 809;
        ELSIF x =- 854 THEN
            tanh_f := - 808;
        ELSIF x =- 853 THEN
            tanh_f := - 807;
        ELSIF x =- 852 THEN
            tanh_f := - 806;
        ELSIF x =- 851 THEN
            tanh_f := - 805;
        ELSIF x =- 850 THEN
            tanh_f := - 804;
        ELSIF x =- 849 THEN
            tanh_f := - 804;
        ELSIF x =- 848 THEN
            tanh_f := - 803;
        ELSIF x =- 847 THEN
            tanh_f := - 802;
        ELSIF x =- 846 THEN
            tanh_f := - 801;
        ELSIF x =- 845 THEN
            tanh_f := - 800;
        ELSIF x =- 844 THEN
            tanh_f := - 799;
        ELSIF x =- 843 THEN
            tanh_f := - 799;
        ELSIF x =- 842 THEN
            tanh_f := - 798;
        ELSIF x =- 841 THEN
            tanh_f := - 797;
        ELSIF x =- 840 THEN
            tanh_f := - 796;
        ELSIF x =- 839 THEN
            tanh_f := - 795;
        ELSIF x =- 838 THEN
            tanh_f := - 794;
        ELSIF x =- 837 THEN
            tanh_f := - 794;
        ELSIF x =- 836 THEN
            tanh_f := - 793;
        ELSIF x =- 835 THEN
            tanh_f := - 792;
        ELSIF x =- 834 THEN
            tanh_f := - 791;
        ELSIF x =- 833 THEN
            tanh_f := - 790;
        ELSIF x =- 832 THEN
            tanh_f := - 789;
        ELSIF x =- 831 THEN
            tanh_f := - 789;
        ELSIF x =- 830 THEN
            tanh_f := - 788;
        ELSIF x =- 829 THEN
            tanh_f := - 787;
        ELSIF x =- 828 THEN
            tanh_f := - 786;
        ELSIF x =- 827 THEN
            tanh_f := - 785;
        ELSIF x =- 826 THEN
            tanh_f := - 785;
        ELSIF x =- 825 THEN
            tanh_f := - 784;
        ELSIF x =- 824 THEN
            tanh_f := - 783;
        ELSIF x =- 823 THEN
            tanh_f := - 782;
        ELSIF x =- 822 THEN
            tanh_f := - 781;
        ELSIF x =- 821 THEN
            tanh_f := - 780;
        ELSIF x =- 820 THEN
            tanh_f := - 780;
        ELSIF x =- 819 THEN
            tanh_f := - 779;
        ELSIF x =- 818 THEN
            tanh_f := - 778;
        ELSIF x =- 817 THEN
            tanh_f := - 777;
        ELSIF x =- 816 THEN
            tanh_f := - 776;
        ELSIF x =- 815 THEN
            tanh_f := - 775;
        ELSIF x =- 814 THEN
            tanh_f := - 775;
        ELSIF x =- 813 THEN
            tanh_f := - 774;
        ELSIF x =- 812 THEN
            tanh_f := - 773;
        ELSIF x =- 811 THEN
            tanh_f := - 772;
        ELSIF x =- 810 THEN
            tanh_f := - 771;
        ELSIF x =- 809 THEN
            tanh_f := - 770;
        ELSIF x =- 808 THEN
            tanh_f := - 770;
        ELSIF x =- 807 THEN
            tanh_f := - 769;
        ELSIF x =- 806 THEN
            tanh_f := - 768;
        ELSIF x =- 805 THEN
            tanh_f := - 767;
        ELSIF x =- 804 THEN
            tanh_f := - 766;
        ELSIF x =- 803 THEN
            tanh_f := - 765;
        ELSIF x =- 802 THEN
            tanh_f := - 765;
        ELSIF x =- 801 THEN
            tanh_f := - 764;
        ELSIF x =- 800 THEN
            tanh_f := - 763;
        ELSIF x =- 799 THEN
            tanh_f := - 762;
        ELSIF x =- 798 THEN
            tanh_f := - 761;
        ELSIF x =- 797 THEN
            tanh_f := - 761;
        ELSIF x =- 796 THEN
            tanh_f := - 760;
        ELSIF x =- 795 THEN
            tanh_f := - 759;
        ELSIF x =- 794 THEN
            tanh_f := - 758;
        ELSIF x =- 793 THEN
            tanh_f := - 757;
        ELSIF x =- 792 THEN
            tanh_f := - 756;
        ELSIF x =- 791 THEN
            tanh_f := - 756;
        ELSIF x =- 790 THEN
            tanh_f := - 755;
        ELSIF x =- 789 THEN
            tanh_f := - 754;
        ELSIF x =- 788 THEN
            tanh_f := - 753;
        ELSIF x =- 787 THEN
            tanh_f := - 752;
        ELSIF x =- 786 THEN
            tanh_f := - 751;
        ELSIF x =- 785 THEN
            tanh_f := - 751;
        ELSIF x =- 784 THEN
            tanh_f := - 750;
        ELSIF x =- 783 THEN
            tanh_f := - 749;
        ELSIF x =- 782 THEN
            tanh_f := - 748;
        ELSIF x =- 781 THEN
            tanh_f := - 747;
        ELSIF x =- 780 THEN
            tanh_f := - 746;
        ELSIF x =- 779 THEN
            tanh_f := - 746;
        ELSIF x =- 778 THEN
            tanh_f := - 745;
        ELSIF x =- 777 THEN
            tanh_f := - 744;
        ELSIF x =- 776 THEN
            tanh_f := - 743;
        ELSIF x =- 775 THEN
            tanh_f := - 742;
        ELSIF x =- 774 THEN
            tanh_f := - 741;
        ELSIF x =- 773 THEN
            tanh_f := - 741;
        ELSIF x =- 772 THEN
            tanh_f := - 740;
        ELSIF x =- 771 THEN
            tanh_f := - 739;
        ELSIF x =- 770 THEN
            tanh_f := - 738;
        ELSIF x =- 769 THEN
            tanh_f := - 737;
        ELSIF x =- 768 THEN
            tanh_f := - 736;
        ELSIF x =- 767 THEN
            tanh_f := - 735;
        ELSIF x =- 766 THEN
            tanh_f := - 734;
        ELSIF x =- 765 THEN
            tanh_f := - 733;
        ELSIF x =- 764 THEN
            tanh_f := - 732;
        ELSIF x =- 763 THEN
            tanh_f := - 731;
        ELSIF x =- 762 THEN
            tanh_f := - 731;
        ELSIF x =- 761 THEN
            tanh_f := - 730;
        ELSIF x =- 760 THEN
            tanh_f := - 729;
        ELSIF x =- 759 THEN
            tanh_f := - 728;
        ELSIF x =- 758 THEN
            tanh_f := - 727;
        ELSIF x =- 757 THEN
            tanh_f := - 726;
        ELSIF x =- 756 THEN
            tanh_f := - 725;
        ELSIF x =- 755 THEN
            tanh_f := - 724;
        ELSIF x =- 754 THEN
            tanh_f := - 723;
        ELSIF x =- 753 THEN
            tanh_f := - 722;
        ELSIF x =- 752 THEN
            tanh_f := - 721;
        ELSIF x =- 751 THEN
            tanh_f := - 721;
        ELSIF x =- 750 THEN
            tanh_f := - 720;
        ELSIF x =- 749 THEN
            tanh_f := - 719;
        ELSIF x =- 748 THEN
            tanh_f := - 718;
        ELSIF x =- 747 THEN
            tanh_f := - 717;
        ELSIF x =- 746 THEN
            tanh_f := - 716;
        ELSIF x =- 745 THEN
            tanh_f := - 715;
        ELSIF x =- 744 THEN
            tanh_f := - 714;
        ELSIF x =- 743 THEN
            tanh_f := - 713;
        ELSIF x =- 742 THEN
            tanh_f := - 712;
        ELSIF x =- 741 THEN
            tanh_f := - 711;
        ELSIF x =- 740 THEN
            tanh_f := - 711;
        ELSIF x =- 739 THEN
            tanh_f := - 710;
        ELSIF x =- 738 THEN
            tanh_f := - 709;
        ELSIF x =- 737 THEN
            tanh_f := - 708;
        ELSIF x =- 736 THEN
            tanh_f := - 707;
        ELSIF x =- 735 THEN
            tanh_f := - 706;
        ELSIF x =- 734 THEN
            tanh_f := - 705;
        ELSIF x =- 733 THEN
            tanh_f := - 704;
        ELSIF x =- 732 THEN
            tanh_f := - 703;
        ELSIF x =- 731 THEN
            tanh_f := - 702;
        ELSIF x =- 730 THEN
            tanh_f := - 701;
        ELSIF x =- 729 THEN
            tanh_f := - 701;
        ELSIF x =- 728 THEN
            tanh_f := - 700;
        ELSIF x =- 727 THEN
            tanh_f := - 699;
        ELSIF x =- 726 THEN
            tanh_f := - 698;
        ELSIF x =- 725 THEN
            tanh_f := - 697;
        ELSIF x =- 724 THEN
            tanh_f := - 696;
        ELSIF x =- 723 THEN
            tanh_f := - 695;
        ELSIF x =- 722 THEN
            tanh_f := - 694;
        ELSIF x =- 721 THEN
            tanh_f := - 693;
        ELSIF x =- 720 THEN
            tanh_f := - 692;
        ELSIF x =- 719 THEN
            tanh_f := - 691;
        ELSIF x =- 718 THEN
            tanh_f := - 691;
        ELSIF x =- 717 THEN
            tanh_f := - 690;
        ELSIF x =- 716 THEN
            tanh_f := - 689;
        ELSIF x =- 715 THEN
            tanh_f := - 688;
        ELSIF x =- 714 THEN
            tanh_f := - 687;
        ELSIF x =- 713 THEN
            tanh_f := - 686;
        ELSIF x =- 712 THEN
            tanh_f := - 685;
        ELSIF x =- 711 THEN
            tanh_f := - 684;
        ELSIF x =- 710 THEN
            tanh_f := - 683;
        ELSIF x =- 709 THEN
            tanh_f := - 682;
        ELSIF x =- 708 THEN
            tanh_f := - 682;
        ELSIF x =- 707 THEN
            tanh_f := - 681;
        ELSIF x =- 706 THEN
            tanh_f := - 680;
        ELSIF x =- 705 THEN
            tanh_f := - 679;
        ELSIF x =- 704 THEN
            tanh_f := - 678;
        ELSIF x =- 703 THEN
            tanh_f := - 677;
        ELSIF x =- 702 THEN
            tanh_f := - 676;
        ELSIF x =- 701 THEN
            tanh_f := - 675;
        ELSIF x =- 700 THEN
            tanh_f := - 674;
        ELSIF x =- 699 THEN
            tanh_f := - 673;
        ELSIF x =- 698 THEN
            tanh_f := - 672;
        ELSIF x =- 697 THEN
            tanh_f := - 672;
        ELSIF x =- 696 THEN
            tanh_f := - 671;
        ELSIF x =- 695 THEN
            tanh_f := - 670;
        ELSIF x =- 694 THEN
            tanh_f := - 669;
        ELSIF x =- 693 THEN
            tanh_f := - 668;
        ELSIF x =- 692 THEN
            tanh_f := - 667;
        ELSIF x =- 691 THEN
            tanh_f := - 666;
        ELSIF x =- 690 THEN
            tanh_f := - 665;
        ELSIF x =- 689 THEN
            tanh_f := - 664;
        ELSIF x =- 688 THEN
            tanh_f := - 663;
        ELSIF x =- 687 THEN
            tanh_f := - 662;
        ELSIF x =- 686 THEN
            tanh_f := - 662;
        ELSIF x =- 685 THEN
            tanh_f := - 661;
        ELSIF x =- 684 THEN
            tanh_f := - 660;
        ELSIF x =- 683 THEN
            tanh_f := - 659;
        ELSIF x =- 682 THEN
            tanh_f := - 658;
        ELSIF x =- 681 THEN
            tanh_f := - 657;
        ELSIF x =- 680 THEN
            tanh_f := - 656;
        ELSIF x =- 679 THEN
            tanh_f := - 655;
        ELSIF x =- 678 THEN
            tanh_f := - 654;
        ELSIF x =- 677 THEN
            tanh_f := - 653;
        ELSIF x =- 676 THEN
            tanh_f := - 652;
        ELSIF x =- 675 THEN
            tanh_f := - 652;
        ELSIF x =- 674 THEN
            tanh_f := - 651;
        ELSIF x =- 673 THEN
            tanh_f := - 650;
        ELSIF x =- 672 THEN
            tanh_f := - 649;
        ELSIF x =- 671 THEN
            tanh_f := - 648;
        ELSIF x =- 670 THEN
            tanh_f := - 647;
        ELSIF x =- 669 THEN
            tanh_f := - 646;
        ELSIF x =- 668 THEN
            tanh_f := - 645;
        ELSIF x =- 667 THEN
            tanh_f := - 644;
        ELSIF x =- 666 THEN
            tanh_f := - 643;
        ELSIF x =- 665 THEN
            tanh_f := - 642;
        ELSIF x =- 664 THEN
            tanh_f := - 642;
        ELSIF x =- 663 THEN
            tanh_f := - 641;
        ELSIF x =- 662 THEN
            tanh_f := - 640;
        ELSIF x =- 661 THEN
            tanh_f := - 639;
        ELSIF x =- 660 THEN
            tanh_f := - 638;
        ELSIF x =- 659 THEN
            tanh_f := - 637;
        ELSIF x =- 658 THEN
            tanh_f := - 636;
        ELSIF x =- 657 THEN
            tanh_f := - 635;
        ELSIF x =- 656 THEN
            tanh_f := - 634;
        ELSIF x =- 655 THEN
            tanh_f := - 633;
        ELSIF x =- 654 THEN
            tanh_f := - 632;
        ELSIF x =- 653 THEN
            tanh_f := - 632;
        ELSIF x =- 652 THEN
            tanh_f := - 631;
        ELSIF x =- 651 THEN
            tanh_f := - 630;
        ELSIF x =- 650 THEN
            tanh_f := - 629;
        ELSIF x =- 649 THEN
            tanh_f := - 628;
        ELSIF x =- 648 THEN
            tanh_f := - 627;
        ELSIF x =- 647 THEN
            tanh_f := - 626;
        ELSIF x =- 646 THEN
            tanh_f := - 625;
        ELSIF x =- 645 THEN
            tanh_f := - 624;
        ELSIF x =- 644 THEN
            tanh_f := - 623;
        ELSIF x =- 643 THEN
            tanh_f := - 622;
        ELSIF x =- 642 THEN
            tanh_f := - 622;
        ELSIF x =- 641 THEN
            tanh_f := - 621;
        ELSIF x =- 640 THEN
            tanh_f := - 620;
        ELSIF x =- 639 THEN
            tanh_f := - 619;
        ELSIF x =- 638 THEN
            tanh_f := - 618;
        ELSIF x =- 637 THEN
            tanh_f := - 617;
        ELSIF x =- 636 THEN
            tanh_f := - 616;
        ELSIF x =- 635 THEN
            tanh_f := - 615;
        ELSIF x =- 634 THEN
            tanh_f := - 614;
        ELSIF x =- 633 THEN
            tanh_f := - 613;
        ELSIF x =- 632 THEN
            tanh_f := - 612;
        ELSIF x =- 631 THEN
            tanh_f := - 612;
        ELSIF x =- 630 THEN
            tanh_f := - 611;
        ELSIF x =- 629 THEN
            tanh_f := - 610;
        ELSIF x =- 628 THEN
            tanh_f := - 609;
        ELSIF x =- 627 THEN
            tanh_f := - 608;
        ELSIF x =- 626 THEN
            tanh_f := - 607;
        ELSIF x =- 625 THEN
            tanh_f := - 606;
        ELSIF x =- 624 THEN
            tanh_f := - 605;
        ELSIF x =- 623 THEN
            tanh_f := - 604;
        ELSIF x =- 622 THEN
            tanh_f := - 603;
        ELSIF x =- 621 THEN
            tanh_f := - 602;
        ELSIF x =- 620 THEN
            tanh_f := - 602;
        ELSIF x =- 619 THEN
            tanh_f := - 601;
        ELSIF x =- 618 THEN
            tanh_f := - 600;
        ELSIF x =- 617 THEN
            tanh_f := - 599;
        ELSIF x =- 616 THEN
            tanh_f := - 598;
        ELSIF x =- 615 THEN
            tanh_f := - 597;
        ELSIF x =- 614 THEN
            tanh_f := - 596;
        ELSIF x =- 613 THEN
            tanh_f := - 595;
        ELSIF x =- 612 THEN
            tanh_f := - 594;
        ELSIF x =- 611 THEN
            tanh_f := - 593;
        ELSIF x =- 610 THEN
            tanh_f := - 593;
        ELSIF x =- 609 THEN
            tanh_f := - 592;
        ELSIF x =- 608 THEN
            tanh_f := - 591;
        ELSIF x =- 607 THEN
            tanh_f := - 590;
        ELSIF x =- 606 THEN
            tanh_f := - 589;
        ELSIF x =- 605 THEN
            tanh_f := - 588;
        ELSIF x =- 604 THEN
            tanh_f := - 587;
        ELSIF x =- 603 THEN
            tanh_f := - 586;
        ELSIF x =- 602 THEN
            tanh_f := - 585;
        ELSIF x =- 601 THEN
            tanh_f := - 584;
        ELSIF x =- 600 THEN
            tanh_f := - 583;
        ELSIF x =- 599 THEN
            tanh_f := - 583;
        ELSIF x =- 598 THEN
            tanh_f := - 582;
        ELSIF x =- 597 THEN
            tanh_f := - 581;
        ELSIF x =- 596 THEN
            tanh_f := - 580;
        ELSIF x =- 595 THEN
            tanh_f := - 579;
        ELSIF x =- 594 THEN
            tanh_f := - 578;
        ELSIF x =- 593 THEN
            tanh_f := - 577;
        ELSIF x =- 592 THEN
            tanh_f := - 576;
        ELSIF x =- 591 THEN
            tanh_f := - 575;
        ELSIF x =- 590 THEN
            tanh_f := - 574;
        ELSIF x =- 589 THEN
            tanh_f := - 573;
        ELSIF x =- 588 THEN
            tanh_f := - 573;
        ELSIF x =- 587 THEN
            tanh_f := - 572;
        ELSIF x =- 586 THEN
            tanh_f := - 571;
        ELSIF x =- 585 THEN
            tanh_f := - 570;
        ELSIF x =- 584 THEN
            tanh_f := - 569;
        ELSIF x =- 583 THEN
            tanh_f := - 568;
        ELSIF x =- 582 THEN
            tanh_f := - 567;
        ELSIF x =- 581 THEN
            tanh_f := - 566;
        ELSIF x =- 580 THEN
            tanh_f := - 565;
        ELSIF x =- 579 THEN
            tanh_f := - 564;
        ELSIF x =- 578 THEN
            tanh_f := - 563;
        ELSIF x =- 577 THEN
            tanh_f := - 563;
        ELSIF x =- 576 THEN
            tanh_f := - 562;
        ELSIF x =- 575 THEN
            tanh_f := - 561;
        ELSIF x =- 574 THEN
            tanh_f := - 560;
        ELSIF x =- 573 THEN
            tanh_f := - 559;
        ELSIF x =- 572 THEN
            tanh_f := - 558;
        ELSIF x =- 571 THEN
            tanh_f := - 557;
        ELSIF x =- 570 THEN
            tanh_f := - 556;
        ELSIF x =- 569 THEN
            tanh_f := - 555;
        ELSIF x =- 568 THEN
            tanh_f := - 554;
        ELSIF x =- 567 THEN
            tanh_f := - 553;
        ELSIF x =- 566 THEN
            tanh_f := - 553;
        ELSIF x =- 565 THEN
            tanh_f := - 552;
        ELSIF x =- 564 THEN
            tanh_f := - 551;
        ELSIF x =- 563 THEN
            tanh_f := - 550;
        ELSIF x =- 562 THEN
            tanh_f := - 549;
        ELSIF x =- 561 THEN
            tanh_f := - 548;
        ELSIF x =- 560 THEN
            tanh_f := - 547;
        ELSIF x =- 559 THEN
            tanh_f := - 546;
        ELSIF x =- 558 THEN
            tanh_f := - 545;
        ELSIF x =- 557 THEN
            tanh_f := - 544;
        ELSIF x =- 556 THEN
            tanh_f := - 543;
        ELSIF x =- 555 THEN
            tanh_f := - 543;
        ELSIF x =- 554 THEN
            tanh_f := - 542;
        ELSIF x =- 553 THEN
            tanh_f := - 541;
        ELSIF x =- 552 THEN
            tanh_f := - 540;
        ELSIF x =- 551 THEN
            tanh_f := - 539;
        ELSIF x =- 550 THEN
            tanh_f := - 538;
        ELSIF x =- 549 THEN
            tanh_f := - 537;
        ELSIF x =- 548 THEN
            tanh_f := - 536;
        ELSIF x =- 547 THEN
            tanh_f := - 535;
        ELSIF x =- 546 THEN
            tanh_f := - 534;
        ELSIF x =- 545 THEN
            tanh_f := - 533;
        ELSIF x =- 544 THEN
            tanh_f := - 533;
        ELSIF x =- 543 THEN
            tanh_f := - 532;
        ELSIF x =- 542 THEN
            tanh_f := - 531;
        ELSIF x =- 541 THEN
            tanh_f := - 530;
        ELSIF x =- 540 THEN
            tanh_f := - 529;
        ELSIF x =- 539 THEN
            tanh_f := - 528;
        ELSIF x =- 538 THEN
            tanh_f := - 527;
        ELSIF x =- 537 THEN
            tanh_f := - 526;
        ELSIF x =- 536 THEN
            tanh_f := - 525;
        ELSIF x =- 535 THEN
            tanh_f := - 524;
        ELSIF x =- 534 THEN
            tanh_f := - 523;
        ELSIF x =- 533 THEN
            tanh_f := - 523;
        ELSIF x =- 532 THEN
            tanh_f := - 522;
        ELSIF x =- 531 THEN
            tanh_f := - 521;
        ELSIF x =- 530 THEN
            tanh_f := - 520;
        ELSIF x =- 529 THEN
            tanh_f := - 519;
        ELSIF x =- 528 THEN
            tanh_f := - 518;
        ELSIF x =- 527 THEN
            tanh_f := - 517;
        ELSIF x =- 526 THEN
            tanh_f := - 516;
        ELSIF x =- 525 THEN
            tanh_f := - 515;
        ELSIF x =- 524 THEN
            tanh_f := - 514;
        ELSIF x =- 523 THEN
            tanh_f := - 513;
        ELSIF x =- 522 THEN
            tanh_f := - 513;
        ELSIF x =- 521 THEN
            tanh_f := - 512;
        ELSIF x =- 520 THEN
            tanh_f := - 511;
        ELSIF x =- 519 THEN
            tanh_f := - 510;
        ELSIF x =- 518 THEN
            tanh_f := - 509;
        ELSIF x =- 517 THEN
            tanh_f := - 508;
        ELSIF x =- 516 THEN
            tanh_f := - 507;
        ELSIF x =- 515 THEN
            tanh_f := - 506;
        ELSIF x =- 514 THEN
            tanh_f := - 505;
        ELSIF x =- 513 THEN
            tanh_f := - 504;
        ELSIF x =- 512 THEN
            tanh_f := - 503;
        ELSIF x =- 511 THEN
            tanh_f := - 503;
        ELSIF x =- 510 THEN
            tanh_f := - 502;
        ELSIF x =- 509 THEN
            tanh_f := - 501;
        ELSIF x =- 508 THEN
            tanh_f := - 500;
        ELSIF x =- 507 THEN
            tanh_f := - 499;
        ELSIF x =- 506 THEN
            tanh_f := - 498;
        ELSIF x =- 505 THEN
            tanh_f := - 497;
        ELSIF x =- 504 THEN
            tanh_f := - 496;
        ELSIF x =- 503 THEN
            tanh_f := - 495;
        ELSIF x =- 502 THEN
            tanh_f := - 494;
        ELSIF x =- 501 THEN
            tanh_f := - 493;
        ELSIF x =- 500 THEN
            tanh_f := - 492;
        ELSIF x =- 499 THEN
            tanh_f := - 491;
        ELSIF x =- 498 THEN
            tanh_f := - 490;
        ELSIF x =- 497 THEN
            tanh_f := - 489;
        ELSIF x =- 496 THEN
            tanh_f := - 488;
        ELSIF x =- 495 THEN
            tanh_f := - 487;
        ELSIF x =- 494 THEN
            tanh_f := - 486;
        ELSIF x =- 493 THEN
            tanh_f := - 485;
        ELSIF x =- 492 THEN
            tanh_f := - 484;
        ELSIF x =- 491 THEN
            tanh_f := - 483;
        ELSIF x =- 490 THEN
            tanh_f := - 482;
        ELSIF x =- 489 THEN
            tanh_f := - 481;
        ELSIF x =- 488 THEN
            tanh_f := - 480;
        ELSIF x =- 487 THEN
            tanh_f := - 479;
        ELSIF x =- 486 THEN
            tanh_f := - 478;
        ELSIF x =- 485 THEN
            tanh_f := - 477;
        ELSIF x =- 484 THEN
            tanh_f := - 476;
        ELSIF x =- 483 THEN
            tanh_f := - 475;
        ELSIF x =- 482 THEN
            tanh_f := - 474;
        ELSIF x =- 481 THEN
            tanh_f := - 474;
        ELSIF x =- 480 THEN
            tanh_f := - 473;
        ELSIF x =- 479 THEN
            tanh_f := - 472;
        ELSIF x =- 478 THEN
            tanh_f := - 471;
        ELSIF x =- 477 THEN
            tanh_f := - 470;
        ELSIF x =- 476 THEN
            tanh_f := - 469;
        ELSIF x =- 475 THEN
            tanh_f := - 468;
        ELSIF x =- 474 THEN
            tanh_f := - 467;
        ELSIF x =- 473 THEN
            tanh_f := - 466;
        ELSIF x =- 472 THEN
            tanh_f := - 465;
        ELSIF x =- 471 THEN
            tanh_f := - 464;
        ELSIF x =- 470 THEN
            tanh_f := - 463;
        ELSIF x =- 469 THEN
            tanh_f := - 462;
        ELSIF x =- 468 THEN
            tanh_f := - 461;
        ELSIF x =- 467 THEN
            tanh_f := - 460;
        ELSIF x =- 466 THEN
            tanh_f := - 459;
        ELSIF x =- 465 THEN
            tanh_f := - 458;
        ELSIF x =- 464 THEN
            tanh_f := - 457;
        ELSIF x =- 463 THEN
            tanh_f := - 456;
        ELSIF x =- 462 THEN
            tanh_f := - 455;
        ELSIF x =- 461 THEN
            tanh_f := - 454;
        ELSIF x =- 460 THEN
            tanh_f := - 453;
        ELSIF x =- 459 THEN
            tanh_f := - 452;
        ELSIF x =- 458 THEN
            tanh_f := - 451;
        ELSIF x =- 457 THEN
            tanh_f := - 450;
        ELSIF x =- 456 THEN
            tanh_f := - 449;
        ELSIF x =- 455 THEN
            tanh_f := - 448;
        ELSIF x =- 454 THEN
            tanh_f := - 447;
        ELSIF x =- 453 THEN
            tanh_f := - 446;
        ELSIF x =- 452 THEN
            tanh_f := - 445;
        ELSIF x =- 451 THEN
            tanh_f := - 445;
        ELSIF x =- 450 THEN
            tanh_f := - 444;
        ELSIF x =- 449 THEN
            tanh_f := - 443;
        ELSIF x =- 448 THEN
            tanh_f := - 442;
        ELSIF x =- 447 THEN
            tanh_f := - 441;
        ELSIF x =- 446 THEN
            tanh_f := - 440;
        ELSIF x =- 445 THEN
            tanh_f := - 439;
        ELSIF x =- 444 THEN
            tanh_f := - 438;
        ELSIF x =- 443 THEN
            tanh_f := - 437;
        ELSIF x =- 442 THEN
            tanh_f := - 436;
        ELSIF x =- 441 THEN
            tanh_f := - 435;
        ELSIF x =- 440 THEN
            tanh_f := - 434;
        ELSIF x =- 439 THEN
            tanh_f := - 433;
        ELSIF x =- 438 THEN
            tanh_f := - 432;
        ELSIF x =- 437 THEN
            tanh_f := - 431;
        ELSIF x =- 436 THEN
            tanh_f := - 430;
        ELSIF x =- 435 THEN
            tanh_f := - 429;
        ELSIF x =- 434 THEN
            tanh_f := - 428;
        ELSIF x =- 433 THEN
            tanh_f := - 427;
        ELSIF x =- 432 THEN
            tanh_f := - 426;
        ELSIF x =- 431 THEN
            tanh_f := - 425;
        ELSIF x =- 430 THEN
            tanh_f := - 424;
        ELSIF x =- 429 THEN
            tanh_f := - 423;
        ELSIF x =- 428 THEN
            tanh_f := - 422;
        ELSIF x =- 427 THEN
            tanh_f := - 421;
        ELSIF x =- 426 THEN
            tanh_f := - 420;
        ELSIF x =- 425 THEN
            tanh_f := - 419;
        ELSIF x =- 424 THEN
            tanh_f := - 418;
        ELSIF x =- 423 THEN
            tanh_f := - 417;
        ELSIF x =- 422 THEN
            tanh_f := - 416;
        ELSIF x =- 421 THEN
            tanh_f := - 416;
        ELSIF x =- 420 THEN
            tanh_f := - 415;
        ELSIF x =- 419 THEN
            tanh_f := - 414;
        ELSIF x =- 418 THEN
            tanh_f := - 413;
        ELSIF x =- 417 THEN
            tanh_f := - 412;
        ELSIF x =- 416 THEN
            tanh_f := - 411;
        ELSIF x =- 415 THEN
            tanh_f := - 410;
        ELSIF x =- 414 THEN
            tanh_f := - 409;
        ELSIF x =- 413 THEN
            tanh_f := - 408;
        ELSIF x =- 412 THEN
            tanh_f := - 407;
        ELSIF x =- 411 THEN
            tanh_f := - 406;
        ELSIF x =- 410 THEN
            tanh_f := - 405;
        ELSIF x =- 409 THEN
            tanh_f := - 404;
        ELSIF x =- 408 THEN
            tanh_f := - 403;
        ELSIF x =- 407 THEN
            tanh_f := - 402;
        ELSIF x =- 406 THEN
            tanh_f := - 401;
        ELSIF x =- 405 THEN
            tanh_f := - 400;
        ELSIF x =- 404 THEN
            tanh_f := - 399;
        ELSIF x =- 403 THEN
            tanh_f := - 398;
        ELSIF x =- 402 THEN
            tanh_f := - 397;
        ELSIF x =- 401 THEN
            tanh_f := - 396;
        ELSIF x =- 400 THEN
            tanh_f := - 395;
        ELSIF x =- 399 THEN
            tanh_f := - 394;
        ELSIF x =- 398 THEN
            tanh_f := - 393;
        ELSIF x =- 397 THEN
            tanh_f := - 392;
        ELSIF x =- 396 THEN
            tanh_f := - 391;
        ELSIF x =- 395 THEN
            tanh_f := - 390;
        ELSIF x =- 394 THEN
            tanh_f := - 389;
        ELSIF x =- 393 THEN
            tanh_f := - 388;
        ELSIF x =- 392 THEN
            tanh_f := - 387;
        ELSIF x =- 391 THEN
            tanh_f := - 387;
        ELSIF x =- 390 THEN
            tanh_f := - 386;
        ELSIF x =- 389 THEN
            tanh_f := - 385;
        ELSIF x =- 388 THEN
            tanh_f := - 384;
        ELSIF x =- 387 THEN
            tanh_f := - 383;
        ELSIF x =- 386 THEN
            tanh_f := - 382;
        ELSIF x =- 385 THEN
            tanh_f := - 381;
        ELSIF x =- 384 THEN
            tanh_f := - 380;
        ELSIF x =- 383 THEN
            tanh_f := - 379;
        ELSIF x =- 382 THEN
            tanh_f := - 378;
        ELSIF x =- 381 THEN
            tanh_f := - 377;
        ELSIF x =- 380 THEN
            tanh_f := - 376;
        ELSIF x =- 379 THEN
            tanh_f := - 375;
        ELSIF x =- 378 THEN
            tanh_f := - 374;
        ELSIF x =- 377 THEN
            tanh_f := - 373;
        ELSIF x =- 376 THEN
            tanh_f := - 372;
        ELSIF x =- 375 THEN
            tanh_f := - 371;
        ELSIF x =- 374 THEN
            tanh_f := - 370;
        ELSIF x =- 373 THEN
            tanh_f := - 369;
        ELSIF x =- 372 THEN
            tanh_f := - 368;
        ELSIF x =- 371 THEN
            tanh_f := - 367;
        ELSIF x =- 370 THEN
            tanh_f := - 366;
        ELSIF x =- 369 THEN
            tanh_f := - 365;
        ELSIF x =- 368 THEN
            tanh_f := - 364;
        ELSIF x =- 367 THEN
            tanh_f := - 363;
        ELSIF x =- 366 THEN
            tanh_f := - 362;
        ELSIF x =- 365 THEN
            tanh_f := - 361;
        ELSIF x =- 364 THEN
            tanh_f := - 360;
        ELSIF x =- 363 THEN
            tanh_f := - 359;
        ELSIF x =- 362 THEN
            tanh_f := - 358;
        ELSIF x =- 361 THEN
            tanh_f := - 358;
        ELSIF x =- 360 THEN
            tanh_f := - 357;
        ELSIF x =- 359 THEN
            tanh_f := - 356;
        ELSIF x =- 358 THEN
            tanh_f := - 355;
        ELSIF x =- 357 THEN
            tanh_f := - 354;
        ELSIF x =- 356 THEN
            tanh_f := - 353;
        ELSIF x =- 355 THEN
            tanh_f := - 352;
        ELSIF x =- 354 THEN
            tanh_f := - 351;
        ELSIF x =- 353 THEN
            tanh_f := - 350;
        ELSIF x =- 352 THEN
            tanh_f := - 349;
        ELSIF x =- 351 THEN
            tanh_f := - 348;
        ELSIF x =- 350 THEN
            tanh_f := - 347;
        ELSIF x =- 349 THEN
            tanh_f := - 346;
        ELSIF x =- 348 THEN
            tanh_f := - 345;
        ELSIF x =- 347 THEN
            tanh_f := - 344;
        ELSIF x =- 346 THEN
            tanh_f := - 343;
        ELSIF x =- 345 THEN
            tanh_f := - 342;
        ELSIF x =- 344 THEN
            tanh_f := - 341;
        ELSIF x =- 343 THEN
            tanh_f := - 340;
        ELSIF x =- 342 THEN
            tanh_f := - 339;
        ELSIF x =- 341 THEN
            tanh_f := - 338;
        ELSIF x =- 340 THEN
            tanh_f := - 337;
        ELSIF x =- 339 THEN
            tanh_f := - 336;
        ELSIF x =- 338 THEN
            tanh_f := - 335;
        ELSIF x =- 337 THEN
            tanh_f := - 334;
        ELSIF x =- 336 THEN
            tanh_f := - 333;
        ELSIF x =- 335 THEN
            tanh_f := - 332;
        ELSIF x =- 334 THEN
            tanh_f := - 331;
        ELSIF x =- 333 THEN
            tanh_f := - 330;
        ELSIF x =- 332 THEN
            tanh_f := - 329;
        ELSIF x =- 331 THEN
            tanh_f := - 329;
        ELSIF x =- 330 THEN
            tanh_f := - 328;
        ELSIF x =- 329 THEN
            tanh_f := - 327;
        ELSIF x =- 328 THEN
            tanh_f := - 326;
        ELSIF x =- 327 THEN
            tanh_f := - 325;
        ELSIF x =- 326 THEN
            tanh_f := - 324;
        ELSIF x =- 325 THEN
            tanh_f := - 323;
        ELSIF x =- 324 THEN
            tanh_f := - 322;
        ELSIF x =- 323 THEN
            tanh_f := - 321;
        ELSIF x =- 322 THEN
            tanh_f := - 320;
        ELSIF x =- 321 THEN
            tanh_f := - 319;
        ELSIF x =- 320 THEN
            tanh_f := - 318;
        ELSIF x =- 319 THEN
            tanh_f := - 317;
        ELSIF x =- 318 THEN
            tanh_f := - 316;
        ELSIF x =- 317 THEN
            tanh_f := - 315;
        ELSIF x =- 316 THEN
            tanh_f := - 314;
        ELSIF x =- 315 THEN
            tanh_f := - 313;
        ELSIF x =- 314 THEN
            tanh_f := - 312;
        ELSIF x =- 313 THEN
            tanh_f := - 311;
        ELSIF x =- 312 THEN
            tanh_f := - 310;
        ELSIF x =- 311 THEN
            tanh_f := - 309;
        ELSIF x =- 310 THEN
            tanh_f := - 308;
        ELSIF x =- 309 THEN
            tanh_f := - 307;
        ELSIF x =- 308 THEN
            tanh_f := - 306;
        ELSIF x =- 307 THEN
            tanh_f := - 305;
        ELSIF x =- 306 THEN
            tanh_f := - 304;
        ELSIF x =- 305 THEN
            tanh_f := - 303;
        ELSIF x =- 304 THEN
            tanh_f := - 302;
        ELSIF x =- 303 THEN
            tanh_f := - 301;
        ELSIF x =- 302 THEN
            tanh_f := - 300;
        ELSIF x =- 301 THEN
            tanh_f := - 300;
        ELSIF x =- 300 THEN
            tanh_f := - 299;
        ELSIF x =- 299 THEN
            tanh_f := - 298;
        ELSIF x =- 298 THEN
            tanh_f := - 297;
        ELSIF x =- 297 THEN
            tanh_f := - 296;
        ELSIF x =- 296 THEN
            tanh_f := - 295;
        ELSIF x =- 295 THEN
            tanh_f := - 294;
        ELSIF x =- 294 THEN
            tanh_f := - 293;
        ELSIF x =- 293 THEN
            tanh_f := - 292;
        ELSIF x =- 292 THEN
            tanh_f := - 291;
        ELSIF x =- 291 THEN
            tanh_f := - 290;
        ELSIF x =- 290 THEN
            tanh_f := - 289;
        ELSIF x =- 289 THEN
            tanh_f := - 288;
        ELSIF x =- 288 THEN
            tanh_f := - 287;
        ELSIF x =- 287 THEN
            tanh_f := - 286;
        ELSIF x =- 286 THEN
            tanh_f := - 285;
        ELSIF x =- 285 THEN
            tanh_f := - 284;
        ELSIF x =- 284 THEN
            tanh_f := - 283;
        ELSIF x =- 283 THEN
            tanh_f := - 282;
        ELSIF x =- 282 THEN
            tanh_f := - 281;
        ELSIF x =- 281 THEN
            tanh_f := - 280;
        ELSIF x =- 280 THEN
            tanh_f := - 279;
        ELSIF x =- 279 THEN
            tanh_f := - 278;
        ELSIF x =- 278 THEN
            tanh_f := - 277;
        ELSIF x =- 277 THEN
            tanh_f := - 276;
        ELSIF x =- 276 THEN
            tanh_f := - 275;
        ELSIF x =- 275 THEN
            tanh_f := - 274;
        ELSIF x =- 274 THEN
            tanh_f := - 273;
        ELSIF x =- 273 THEN
            tanh_f := - 272;
        ELSIF x =- 272 THEN
            tanh_f := - 271;
        ELSIF x =- 271 THEN
            tanh_f := - 271;
        ELSIF x =- 270 THEN
            tanh_f := - 270;
        ELSIF x =- 269 THEN
            tanh_f := - 269;
        ELSIF x =- 268 THEN
            tanh_f := - 268;
        ELSIF x =- 267 THEN
            tanh_f := - 267;
        ELSIF x =- 266 THEN
            tanh_f := - 266;
        ELSIF x =- 265 THEN
            tanh_f := - 265;
        ELSIF x =- 264 THEN
            tanh_f := - 264;
        ELSIF x =- 263 THEN
            tanh_f := - 263;
        ELSIF x =- 262 THEN
            tanh_f := - 262;
        ELSIF x =- 261 THEN
            tanh_f := - 261;
        ELSIF x =- 260 THEN
            tanh_f := - 260;
        ELSIF x =- 259 THEN
            tanh_f := - 259;
        ELSIF x =- 258 THEN
            tanh_f := - 258;
        ELSIF x =- 257 THEN
            tanh_f := - 257;
        ELSIF x =- 256 THEN
            tanh_f := - 256;
        ELSIF x =- 255 THEN
            tanh_f := - 255;
        ELSIF x =- 254 THEN
            tanh_f := - 254;
        ELSIF x =- 253 THEN
            tanh_f := - 253;
        ELSIF x =- 252 THEN
            tanh_f := - 252;
        ELSIF x =- 251 THEN
            tanh_f := - 251;
        ELSIF x =- 250 THEN
            tanh_f := - 250;
        ELSIF x =- 249 THEN
            tanh_f := - 249;
        ELSIF x =- 248 THEN
            tanh_f := - 248;
        ELSIF x =- 247 THEN
            tanh_f := - 247;
        ELSIF x =- 246 THEN
            tanh_f := - 246;
        ELSIF x =- 245 THEN
            tanh_f := - 245;
        ELSIF x =- 244 THEN
            tanh_f := - 244;
        ELSIF x =- 243 THEN
            tanh_f := - 243;
        ELSIF x =- 242 THEN
            tanh_f := - 242;
        ELSIF x =- 241 THEN
            tanh_f := - 241;
        ELSIF x =- 240 THEN
            tanh_f := - 240;
        ELSIF x =- 239 THEN
            tanh_f := - 239;
        ELSIF x =- 238 THEN
            tanh_f := - 238;
        ELSIF x =- 237 THEN
            tanh_f := - 237;
        ELSIF x =- 236 THEN
            tanh_f := - 236;
        ELSIF x =- 235 THEN
            tanh_f := - 235;
        ELSIF x =- 234 THEN
            tanh_f := - 234;
        ELSIF x =- 233 THEN
            tanh_f := - 233;
        ELSIF x =- 232 THEN
            tanh_f := - 232;
        ELSIF x =- 231 THEN
            tanh_f := - 231;
        ELSIF x =- 230 THEN
            tanh_f := - 230;
        ELSIF x =- 229 THEN
            tanh_f := - 229;
        ELSIF x =- 228 THEN
            tanh_f := - 228;
        ELSIF x =- 227 THEN
            tanh_f := - 227;
        ELSIF x =- 226 THEN
            tanh_f := - 226;
        ELSIF x =- 225 THEN
            tanh_f := - 225;
        ELSIF x =- 224 THEN
            tanh_f := - 224;
        ELSIF x =- 223 THEN
            tanh_f := - 223;
        ELSIF x =- 222 THEN
            tanh_f := - 222;
        ELSIF x =- 221 THEN
            tanh_f := - 221;
        ELSIF x =- 220 THEN
            tanh_f := - 220;
        ELSIF x =- 219 THEN
            tanh_f := - 219;
        ELSIF x =- 218 THEN
            tanh_f := - 218;
        ELSIF x =- 217 THEN
            tanh_f := - 217;
        ELSIF x =- 216 THEN
            tanh_f := - 216;
        ELSIF x =- 215 THEN
            tanh_f := - 215;
        ELSIF x =- 214 THEN
            tanh_f := - 214;
        ELSIF x =- 213 THEN
            tanh_f := - 213;
        ELSIF x =- 212 THEN
            tanh_f := - 212;
        ELSIF x =- 211 THEN
            tanh_f := - 211;
        ELSIF x =- 210 THEN
            tanh_f := - 210;
        ELSIF x =- 209 THEN
            tanh_f := - 209;
        ELSIF x =- 208 THEN
            tanh_f := - 208;
        ELSIF x =- 207 THEN
            tanh_f := - 207;
        ELSIF x =- 206 THEN
            tanh_f := - 206;
        ELSIF x =- 205 THEN
            tanh_f := - 205;
        ELSIF x =- 204 THEN
            tanh_f := - 204;
        ELSIF x =- 203 THEN
            tanh_f := - 203;
        ELSIF x =- 202 THEN
            tanh_f := - 202;
        ELSIF x =- 201 THEN
            tanh_f := - 201;
        ELSIF x =- 200 THEN
            tanh_f := - 200;
        ELSIF x =- 199 THEN
            tanh_f := - 199;
        ELSIF x =- 198 THEN
            tanh_f := - 198;
        ELSIF x =- 197 THEN
            tanh_f := - 197;
        ELSIF x =- 196 THEN
            tanh_f := - 196;
        ELSIF x =- 195 THEN
            tanh_f := - 195;
        ELSIF x =- 194 THEN
            tanh_f := - 194;
        ELSIF x =- 193 THEN
            tanh_f := - 193;
        ELSIF x =- 192 THEN
            tanh_f := - 192;
        ELSIF x =- 191 THEN
            tanh_f := - 191;
        ELSIF x =- 190 THEN
            tanh_f := - 190;
        ELSIF x =- 189 THEN
            tanh_f := - 189;
        ELSIF x =- 188 THEN
            tanh_f := - 188;
        ELSIF x =- 187 THEN
            tanh_f := - 187;
        ELSIF x =- 186 THEN
            tanh_f := - 186;
        ELSIF x =- 185 THEN
            tanh_f := - 185;
        ELSIF x =- 184 THEN
            tanh_f := - 184;
        ELSIF x =- 183 THEN
            tanh_f := - 183;
        ELSIF x =- 182 THEN
            tanh_f := - 182;
        ELSIF x =- 181 THEN
            tanh_f := - 181;
        ELSIF x =- 180 THEN
            tanh_f := - 180;
        ELSIF x =- 179 THEN
            tanh_f := - 179;
        ELSIF x =- 178 THEN
            tanh_f := - 178;
        ELSIF x =- 177 THEN
            tanh_f := - 177;
        ELSIF x =- 176 THEN
            tanh_f := - 176;
        ELSIF x =- 175 THEN
            tanh_f := - 175;
        ELSIF x =- 174 THEN
            tanh_f := - 174;
        ELSIF x =- 173 THEN
            tanh_f := - 173;
        ELSIF x =- 172 THEN
            tanh_f := - 172;
        ELSIF x =- 171 THEN
            tanh_f := - 171;
        ELSIF x =- 170 THEN
            tanh_f := - 170;
        ELSIF x =- 169 THEN
            tanh_f := - 169;
        ELSIF x =- 168 THEN
            tanh_f := - 168;
        ELSIF x =- 167 THEN
            tanh_f := - 167;
        ELSIF x =- 166 THEN
            tanh_f := - 166;
        ELSIF x =- 165 THEN
            tanh_f := - 165;
        ELSIF x =- 164 THEN
            tanh_f := - 164;
        ELSIF x =- 163 THEN
            tanh_f := - 163;
        ELSIF x =- 162 THEN
            tanh_f := - 162;
        ELSIF x =- 161 THEN
            tanh_f := - 161;
        ELSIF x =- 160 THEN
            tanh_f := - 160;
        ELSIF x =- 159 THEN
            tanh_f := - 159;
        ELSIF x =- 158 THEN
            tanh_f := - 158;
        ELSIF x =- 157 THEN
            tanh_f := - 157;
        ELSIF x =- 156 THEN
            tanh_f := - 156;
        ELSIF x =- 155 THEN
            tanh_f := - 155;
        ELSIF x =- 154 THEN
            tanh_f := - 154;
        ELSIF x =- 153 THEN
            tanh_f := - 153;
        ELSIF x =- 152 THEN
            tanh_f := - 152;
        ELSIF x =- 151 THEN
            tanh_f := - 151;
        ELSIF x =- 150 THEN
            tanh_f := - 150;
        ELSIF x =- 149 THEN
            tanh_f := - 149;
        ELSIF x =- 148 THEN
            tanh_f := - 148;
        ELSIF x =- 147 THEN
            tanh_f := - 147;
        ELSIF x =- 146 THEN
            tanh_f := - 146;
        ELSIF x =- 145 THEN
            tanh_f := - 145;
        ELSIF x =- 144 THEN
            tanh_f := - 144;
        ELSIF x =- 143 THEN
            tanh_f := - 143;
        ELSIF x =- 142 THEN
            tanh_f := - 142;
        ELSIF x =- 141 THEN
            tanh_f := - 141;
        ELSIF x =- 140 THEN
            tanh_f := - 140;
        ELSIF x =- 139 THEN
            tanh_f := - 139;
        ELSIF x =- 138 THEN
            tanh_f := - 138;
        ELSIF x =- 137 THEN
            tanh_f := - 137;
        ELSIF x =- 136 THEN
            tanh_f := - 136;
        ELSIF x =- 135 THEN
            tanh_f := - 135;
        ELSIF x =- 134 THEN
            tanh_f := - 134;
        ELSIF x =- 133 THEN
            tanh_f := - 133;
        ELSIF x =- 132 THEN
            tanh_f := - 132;
        ELSIF x =- 131 THEN
            tanh_f := - 131;
        ELSIF x =- 130 THEN
            tanh_f := - 130;
        ELSIF x =- 129 THEN
            tanh_f := - 129;
        ELSIF x =- 128 THEN
            tanh_f := - 128;
        ELSIF x =- 127 THEN
            tanh_f := - 127;
        ELSIF x =- 126 THEN
            tanh_f := - 126;
        ELSIF x =- 125 THEN
            tanh_f := - 125;
        ELSIF x =- 124 THEN
            tanh_f := - 124;
        ELSIF x =- 123 THEN
            tanh_f := - 123;
        ELSIF x =- 122 THEN
            tanh_f := - 122;
        ELSIF x =- 121 THEN
            tanh_f := - 121;
        ELSIF x =- 120 THEN
            tanh_f := - 120;
        ELSIF x =- 119 THEN
            tanh_f := - 119;
        ELSIF x =- 118 THEN
            tanh_f := - 118;
        ELSIF x =- 117 THEN
            tanh_f := - 117;
        ELSIF x =- 116 THEN
            tanh_f := - 116;
        ELSIF x =- 115 THEN
            tanh_f := - 115;
        ELSIF x =- 114 THEN
            tanh_f := - 114;
        ELSIF x =- 113 THEN
            tanh_f := - 113;
        ELSIF x =- 112 THEN
            tanh_f := - 112;
        ELSIF x =- 111 THEN
            tanh_f := - 111;
        ELSIF x =- 110 THEN
            tanh_f := - 110;
        ELSIF x =- 109 THEN
            tanh_f := - 109;
        ELSIF x =- 108 THEN
            tanh_f := - 108;
        ELSIF x =- 107 THEN
            tanh_f := - 107;
        ELSIF x =- 106 THEN
            tanh_f := - 106;
        ELSIF x =- 105 THEN
            tanh_f := - 105;
        ELSIF x =- 104 THEN
            tanh_f := - 104;
        ELSIF x =- 103 THEN
            tanh_f := - 103;
        ELSIF x =- 102 THEN
            tanh_f := - 102;
        ELSIF x =- 101 THEN
            tanh_f := - 101;
        ELSIF x =- 100 THEN
            tanh_f := - 100;
        ELSIF x =- 99 THEN
            tanh_f := - 99;
        ELSIF x =- 98 THEN
            tanh_f := - 98;
        ELSIF x =- 97 THEN
            tanh_f := - 97;
        ELSIF x =- 96 THEN
            tanh_f := - 96;
        ELSIF x =- 95 THEN
            tanh_f := - 95;
        ELSIF x =- 94 THEN
            tanh_f := - 94;
        ELSIF x =- 93 THEN
            tanh_f := - 93;
        ELSIF x =- 92 THEN
            tanh_f := - 92;
        ELSIF x =- 91 THEN
            tanh_f := - 91;
        ELSIF x =- 90 THEN
            tanh_f := - 90;
        ELSIF x =- 89 THEN
            tanh_f := - 89;
        ELSIF x =- 88 THEN
            tanh_f := - 88;
        ELSIF x =- 87 THEN
            tanh_f := - 87;
        ELSIF x =- 86 THEN
            tanh_f := - 86;
        ELSIF x =- 85 THEN
            tanh_f := - 85;
        ELSIF x =- 84 THEN
            tanh_f := - 84;
        ELSIF x =- 83 THEN
            tanh_f := - 83;
        ELSIF x =- 82 THEN
            tanh_f := - 82;
        ELSIF x =- 81 THEN
            tanh_f := - 81;
        ELSIF x =- 80 THEN
            tanh_f := - 80;
        ELSIF x =- 79 THEN
            tanh_f := - 79;
        ELSIF x =- 78 THEN
            tanh_f := - 78;
        ELSIF x =- 77 THEN
            tanh_f := - 77;
        ELSIF x =- 76 THEN
            tanh_f := - 76;
        ELSIF x =- 75 THEN
            tanh_f := - 75;
        ELSIF x =- 74 THEN
            tanh_f := - 74;
        ELSIF x =- 73 THEN
            tanh_f := - 73;
        ELSIF x =- 72 THEN
            tanh_f := - 72;
        ELSIF x =- 71 THEN
            tanh_f := - 71;
        ELSIF x =- 70 THEN
            tanh_f := - 70;
        ELSIF x =- 69 THEN
            tanh_f := - 69;
        ELSIF x =- 68 THEN
            tanh_f := - 68;
        ELSIF x =- 67 THEN
            tanh_f := - 67;
        ELSIF x =- 66 THEN
            tanh_f := - 66;
        ELSIF x =- 65 THEN
            tanh_f := - 65;
        ELSIF x =- 64 THEN
            tanh_f := - 64;
        ELSIF x =- 63 THEN
            tanh_f := - 63;
        ELSIF x =- 62 THEN
            tanh_f := - 62;
        ELSIF x =- 61 THEN
            tanh_f := - 61;
        ELSIF x =- 60 THEN
            tanh_f := - 60;
        ELSIF x =- 59 THEN
            tanh_f := - 59;
        ELSIF x =- 58 THEN
            tanh_f := - 58;
        ELSIF x =- 57 THEN
            tanh_f := - 57;
        ELSIF x =- 56 THEN
            tanh_f := - 56;
        ELSIF x =- 55 THEN
            tanh_f := - 55;
        ELSIF x =- 54 THEN
            tanh_f := - 54;
        ELSIF x =- 53 THEN
            tanh_f := - 53;
        ELSIF x =- 52 THEN
            tanh_f := - 52;
        ELSIF x =- 51 THEN
            tanh_f := - 51;
        ELSIF x =- 50 THEN
            tanh_f := - 50;
        ELSIF x =- 49 THEN
            tanh_f := - 49;
        ELSIF x =- 48 THEN
            tanh_f := - 48;
        ELSIF x =- 47 THEN
            tanh_f := - 47;
        ELSIF x =- 46 THEN
            tanh_f := - 46;
        ELSIF x =- 45 THEN
            tanh_f := - 45;
        ELSIF x =- 44 THEN
            tanh_f := - 44;
        ELSIF x =- 43 THEN
            tanh_f := - 43;
        ELSIF x =- 42 THEN
            tanh_f := - 42;
        ELSIF x =- 41 THEN
            tanh_f := - 41;
        ELSIF x =- 40 THEN
            tanh_f := - 40;
        ELSIF x =- 39 THEN
            tanh_f := - 39;
        ELSIF x =- 38 THEN
            tanh_f := - 38;
        ELSIF x =- 37 THEN
            tanh_f := - 37;
        ELSIF x =- 36 THEN
            tanh_f := - 36;
        ELSIF x =- 35 THEN
            tanh_f := - 35;
        ELSIF x =- 34 THEN
            tanh_f := - 34;
        ELSIF x =- 33 THEN
            tanh_f := - 33;
        ELSIF x =- 32 THEN
            tanh_f := - 32;
        ELSIF x =- 31 THEN
            tanh_f := - 31;
        ELSIF x =- 30 THEN
            tanh_f := - 30;
        ELSIF x =- 29 THEN
            tanh_f := - 29;
        ELSIF x =- 28 THEN
            tanh_f := - 28;
        ELSIF x =- 27 THEN
            tanh_f := - 27;
        ELSIF x =- 26 THEN
            tanh_f := - 26;
        ELSIF x =- 25 THEN
            tanh_f := - 25;
        ELSIF x =- 24 THEN
            tanh_f := - 24;
        ELSIF x =- 23 THEN
            tanh_f := - 23;
        ELSIF x =- 22 THEN
            tanh_f := - 22;
        ELSIF x =- 21 THEN
            tanh_f := - 21;
        ELSIF x =- 20 THEN
            tanh_f := - 20;
        ELSIF x =- 19 THEN
            tanh_f := - 19;
        ELSIF x =- 18 THEN
            tanh_f := - 18;
        ELSIF x =- 17 THEN
            tanh_f := - 17;
        ELSIF x =- 16 THEN
            tanh_f := - 16;
        ELSIF x =- 15 THEN
            tanh_f := - 15;
        ELSIF x =- 14 THEN
            tanh_f := - 14;
        ELSIF x =- 13 THEN
            tanh_f := - 13;
        ELSIF x =- 12 THEN
            tanh_f := - 12;
        ELSIF x =- 11 THEN
            tanh_f := - 11;
        ELSIF x =- 10 THEN
            tanh_f := - 10;
        ELSIF x =- 9 THEN
            tanh_f := - 9;
        ELSIF x =- 8 THEN
            tanh_f := - 8;
        ELSIF x =- 7 THEN
            tanh_f := - 7;
        ELSIF x =- 6 THEN
            tanh_f := - 6;
        ELSIF x =- 5 THEN
            tanh_f := - 5;
        ELSIF x =- 4 THEN
            tanh_f := - 4;
        ELSIF x =- 3 THEN
            tanh_f := - 3;
        ELSIF x =- 2 THEN
            tanh_f := - 2;
        ELSIF x =- 1 THEN
            tanh_f := - 1;
        ELSIF x = 0 THEN
            tanh_f := 0;
        ELSIF x = 1 THEN
            tanh_f := 1;
        ELSIF x = 2 THEN
            tanh_f := 2;
        ELSIF x = 3 THEN
            tanh_f := 3;
        ELSIF x = 4 THEN
            tanh_f := 4;
        ELSIF x = 5 THEN
            tanh_f := 5;
        ELSIF x = 6 THEN
            tanh_f := 6;
        ELSIF x = 7 THEN
            tanh_f := 7;
        ELSIF x = 8 THEN
            tanh_f := 8;
        ELSIF x = 9 THEN
            tanh_f := 9;
        ELSIF x = 10 THEN
            tanh_f := 10;
        ELSIF x = 11 THEN
            tanh_f := 11;
        ELSIF x = 12 THEN
            tanh_f := 12;
        ELSIF x = 13 THEN
            tanh_f := 13;
        ELSIF x = 14 THEN
            tanh_f := 14;
        ELSIF x = 15 THEN
            tanh_f := 15;
        ELSIF x = 16 THEN
            tanh_f := 16;
        ELSIF x = 17 THEN
            tanh_f := 17;
        ELSIF x = 18 THEN
            tanh_f := 18;
        ELSIF x = 19 THEN
            tanh_f := 19;
        ELSIF x = 20 THEN
            tanh_f := 20;
        ELSIF x = 21 THEN
            tanh_f := 21;
        ELSIF x = 22 THEN
            tanh_f := 22;
        ELSIF x = 23 THEN
            tanh_f := 23;
        ELSIF x = 24 THEN
            tanh_f := 24;
        ELSIF x = 25 THEN
            tanh_f := 25;
        ELSIF x = 26 THEN
            tanh_f := 26;
        ELSIF x = 27 THEN
            tanh_f := 27;
        ELSIF x = 28 THEN
            tanh_f := 28;
        ELSIF x = 29 THEN
            tanh_f := 29;
        ELSIF x = 30 THEN
            tanh_f := 30;
        ELSIF x = 31 THEN
            tanh_f := 31;
        ELSIF x = 32 THEN
            tanh_f := 32;
        ELSIF x = 33 THEN
            tanh_f := 33;
        ELSIF x = 34 THEN
            tanh_f := 34;
        ELSIF x = 35 THEN
            tanh_f := 35;
        ELSIF x = 36 THEN
            tanh_f := 36;
        ELSIF x = 37 THEN
            tanh_f := 37;
        ELSIF x = 38 THEN
            tanh_f := 38;
        ELSIF x = 39 THEN
            tanh_f := 39;
        ELSIF x = 40 THEN
            tanh_f := 40;
        ELSIF x = 41 THEN
            tanh_f := 41;
        ELSIF x = 42 THEN
            tanh_f := 42;
        ELSIF x = 43 THEN
            tanh_f := 43;
        ELSIF x = 44 THEN
            tanh_f := 44;
        ELSIF x = 45 THEN
            tanh_f := 45;
        ELSIF x = 46 THEN
            tanh_f := 46;
        ELSIF x = 47 THEN
            tanh_f := 47;
        ELSIF x = 48 THEN
            tanh_f := 48;
        ELSIF x = 49 THEN
            tanh_f := 49;
        ELSIF x = 50 THEN
            tanh_f := 50;
        ELSIF x = 51 THEN
            tanh_f := 51;
        ELSIF x = 52 THEN
            tanh_f := 52;
        ELSIF x = 53 THEN
            tanh_f := 53;
        ELSIF x = 54 THEN
            tanh_f := 54;
        ELSIF x = 55 THEN
            tanh_f := 55;
        ELSIF x = 56 THEN
            tanh_f := 56;
        ELSIF x = 57 THEN
            tanh_f := 57;
        ELSIF x = 58 THEN
            tanh_f := 58;
        ELSIF x = 59 THEN
            tanh_f := 59;
        ELSIF x = 60 THEN
            tanh_f := 60;
        ELSIF x = 61 THEN
            tanh_f := 61;
        ELSIF x = 62 THEN
            tanh_f := 62;
        ELSIF x = 63 THEN
            tanh_f := 63;
        ELSIF x = 64 THEN
            tanh_f := 64;
        ELSIF x = 65 THEN
            tanh_f := 65;
        ELSIF x = 66 THEN
            tanh_f := 66;
        ELSIF x = 67 THEN
            tanh_f := 67;
        ELSIF x = 68 THEN
            tanh_f := 68;
        ELSIF x = 69 THEN
            tanh_f := 69;
        ELSIF x = 70 THEN
            tanh_f := 70;
        ELSIF x = 71 THEN
            tanh_f := 71;
        ELSIF x = 72 THEN
            tanh_f := 72;
        ELSIF x = 73 THEN
            tanh_f := 73;
        ELSIF x = 74 THEN
            tanh_f := 74;
        ELSIF x = 75 THEN
            tanh_f := 75;
        ELSIF x = 76 THEN
            tanh_f := 76;
        ELSIF x = 77 THEN
            tanh_f := 77;
        ELSIF x = 78 THEN
            tanh_f := 78;
        ELSIF x = 79 THEN
            tanh_f := 79;
        ELSIF x = 80 THEN
            tanh_f := 80;
        ELSIF x = 81 THEN
            tanh_f := 81;
        ELSIF x = 82 THEN
            tanh_f := 82;
        ELSIF x = 83 THEN
            tanh_f := 83;
        ELSIF x = 84 THEN
            tanh_f := 84;
        ELSIF x = 85 THEN
            tanh_f := 85;
        ELSIF x = 86 THEN
            tanh_f := 86;
        ELSIF x = 87 THEN
            tanh_f := 87;
        ELSIF x = 88 THEN
            tanh_f := 88;
        ELSIF x = 89 THEN
            tanh_f := 89;
        ELSIF x = 90 THEN
            tanh_f := 90;
        ELSIF x = 91 THEN
            tanh_f := 91;
        ELSIF x = 92 THEN
            tanh_f := 92;
        ELSIF x = 93 THEN
            tanh_f := 93;
        ELSIF x = 94 THEN
            tanh_f := 94;
        ELSIF x = 95 THEN
            tanh_f := 95;
        ELSIF x = 96 THEN
            tanh_f := 96;
        ELSIF x = 97 THEN
            tanh_f := 97;
        ELSIF x = 98 THEN
            tanh_f := 98;
        ELSIF x = 99 THEN
            tanh_f := 99;
        ELSIF x = 100 THEN
            tanh_f := 100;
        ELSIF x = 101 THEN
            tanh_f := 101;
        ELSIF x = 102 THEN
            tanh_f := 102;
        ELSIF x = 103 THEN
            tanh_f := 103;
        ELSIF x = 104 THEN
            tanh_f := 104;
        ELSIF x = 105 THEN
            tanh_f := 105;
        ELSIF x = 106 THEN
            tanh_f := 106;
        ELSIF x = 107 THEN
            tanh_f := 107;
        ELSIF x = 108 THEN
            tanh_f := 108;
        ELSIF x = 109 THEN
            tanh_f := 109;
        ELSIF x = 110 THEN
            tanh_f := 110;
        ELSIF x = 111 THEN
            tanh_f := 111;
        ELSIF x = 112 THEN
            tanh_f := 112;
        ELSIF x = 113 THEN
            tanh_f := 113;
        ELSIF x = 114 THEN
            tanh_f := 114;
        ELSIF x = 115 THEN
            tanh_f := 115;
        ELSIF x = 116 THEN
            tanh_f := 116;
        ELSIF x = 117 THEN
            tanh_f := 117;
        ELSIF x = 118 THEN
            tanh_f := 118;
        ELSIF x = 119 THEN
            tanh_f := 119;
        ELSIF x = 120 THEN
            tanh_f := 120;
        ELSIF x = 121 THEN
            tanh_f := 121;
        ELSIF x = 122 THEN
            tanh_f := 122;
        ELSIF x = 123 THEN
            tanh_f := 123;
        ELSIF x = 124 THEN
            tanh_f := 124;
        ELSIF x = 125 THEN
            tanh_f := 125;
        ELSIF x = 126 THEN
            tanh_f := 126;
        ELSIF x = 127 THEN
            tanh_f := 127;
        ELSIF x = 128 THEN
            tanh_f := 128;
        ELSIF x = 129 THEN
            tanh_f := 129;
        ELSIF x = 130 THEN
            tanh_f := 130;
        ELSIF x = 131 THEN
            tanh_f := 131;
        ELSIF x = 132 THEN
            tanh_f := 132;
        ELSIF x = 133 THEN
            tanh_f := 133;
        ELSIF x = 134 THEN
            tanh_f := 134;
        ELSIF x = 135 THEN
            tanh_f := 135;
        ELSIF x = 136 THEN
            tanh_f := 136;
        ELSIF x = 137 THEN
            tanh_f := 137;
        ELSIF x = 138 THEN
            tanh_f := 138;
        ELSIF x = 139 THEN
            tanh_f := 139;
        ELSIF x = 140 THEN
            tanh_f := 140;
        ELSIF x = 141 THEN
            tanh_f := 141;
        ELSIF x = 142 THEN
            tanh_f := 142;
        ELSIF x = 143 THEN
            tanh_f := 143;
        ELSIF x = 144 THEN
            tanh_f := 144;
        ELSIF x = 145 THEN
            tanh_f := 145;
        ELSIF x = 146 THEN
            tanh_f := 146;
        ELSIF x = 147 THEN
            tanh_f := 147;
        ELSIF x = 148 THEN
            tanh_f := 148;
        ELSIF x = 149 THEN
            tanh_f := 149;
        ELSIF x = 150 THEN
            tanh_f := 150;
        ELSIF x = 151 THEN
            tanh_f := 151;
        ELSIF x = 152 THEN
            tanh_f := 152;
        ELSIF x = 153 THEN
            tanh_f := 153;
        ELSIF x = 154 THEN
            tanh_f := 154;
        ELSIF x = 155 THEN
            tanh_f := 155;
        ELSIF x = 156 THEN
            tanh_f := 156;
        ELSIF x = 157 THEN
            tanh_f := 157;
        ELSIF x = 158 THEN
            tanh_f := 158;
        ELSIF x = 159 THEN
            tanh_f := 159;
        ELSIF x = 160 THEN
            tanh_f := 160;
        ELSIF x = 161 THEN
            tanh_f := 161;
        ELSIF x = 162 THEN
            tanh_f := 162;
        ELSIF x = 163 THEN
            tanh_f := 163;
        ELSIF x = 164 THEN
            tanh_f := 164;
        ELSIF x = 165 THEN
            tanh_f := 165;
        ELSIF x = 166 THEN
            tanh_f := 166;
        ELSIF x = 167 THEN
            tanh_f := 167;
        ELSIF x = 168 THEN
            tanh_f := 168;
        ELSIF x = 169 THEN
            tanh_f := 169;
        ELSIF x = 170 THEN
            tanh_f := 170;
        ELSIF x = 171 THEN
            tanh_f := 171;
        ELSIF x = 172 THEN
            tanh_f := 172;
        ELSIF x = 173 THEN
            tanh_f := 173;
        ELSIF x = 174 THEN
            tanh_f := 174;
        ELSIF x = 175 THEN
            tanh_f := 175;
        ELSIF x = 176 THEN
            tanh_f := 176;
        ELSIF x = 177 THEN
            tanh_f := 177;
        ELSIF x = 178 THEN
            tanh_f := 178;
        ELSIF x = 179 THEN
            tanh_f := 179;
        ELSIF x = 180 THEN
            tanh_f := 180;
        ELSIF x = 181 THEN
            tanh_f := 181;
        ELSIF x = 182 THEN
            tanh_f := 182;
        ELSIF x = 183 THEN
            tanh_f := 183;
        ELSIF x = 184 THEN
            tanh_f := 184;
        ELSIF x = 185 THEN
            tanh_f := 185;
        ELSIF x = 186 THEN
            tanh_f := 186;
        ELSIF x = 187 THEN
            tanh_f := 187;
        ELSIF x = 188 THEN
            tanh_f := 188;
        ELSIF x = 189 THEN
            tanh_f := 189;
        ELSIF x = 190 THEN
            tanh_f := 190;
        ELSIF x = 191 THEN
            tanh_f := 191;
        ELSIF x = 192 THEN
            tanh_f := 192;
        ELSIF x = 193 THEN
            tanh_f := 193;
        ELSIF x = 194 THEN
            tanh_f := 194;
        ELSIF x = 195 THEN
            tanh_f := 195;
        ELSIF x = 196 THEN
            tanh_f := 196;
        ELSIF x = 197 THEN
            tanh_f := 197;
        ELSIF x = 198 THEN
            tanh_f := 198;
        ELSIF x = 199 THEN
            tanh_f := 199;
        ELSIF x = 200 THEN
            tanh_f := 200;
        ELSIF x = 201 THEN
            tanh_f := 201;
        ELSIF x = 202 THEN
            tanh_f := 202;
        ELSIF x = 203 THEN
            tanh_f := 203;
        ELSIF x = 204 THEN
            tanh_f := 204;
        ELSIF x = 205 THEN
            tanh_f := 205;
        ELSIF x = 206 THEN
            tanh_f := 206;
        ELSIF x = 207 THEN
            tanh_f := 207;
        ELSIF x = 208 THEN
            tanh_f := 208;
        ELSIF x = 209 THEN
            tanh_f := 209;
        ELSIF x = 210 THEN
            tanh_f := 210;
        ELSIF x = 211 THEN
            tanh_f := 211;
        ELSIF x = 212 THEN
            tanh_f := 212;
        ELSIF x = 213 THEN
            tanh_f := 213;
        ELSIF x = 214 THEN
            tanh_f := 214;
        ELSIF x = 215 THEN
            tanh_f := 215;
        ELSIF x = 216 THEN
            tanh_f := 216;
        ELSIF x = 217 THEN
            tanh_f := 217;
        ELSIF x = 218 THEN
            tanh_f := 218;
        ELSIF x = 219 THEN
            tanh_f := 219;
        ELSIF x = 220 THEN
            tanh_f := 220;
        ELSIF x = 221 THEN
            tanh_f := 221;
        ELSIF x = 222 THEN
            tanh_f := 222;
        ELSIF x = 223 THEN
            tanh_f := 223;
        ELSIF x = 224 THEN
            tanh_f := 224;
        ELSIF x = 225 THEN
            tanh_f := 225;
        ELSIF x = 226 THEN
            tanh_f := 226;
        ELSIF x = 227 THEN
            tanh_f := 227;
        ELSIF x = 228 THEN
            tanh_f := 228;
        ELSIF x = 229 THEN
            tanh_f := 229;
        ELSIF x = 230 THEN
            tanh_f := 230;
        ELSIF x = 231 THEN
            tanh_f := 231;
        ELSIF x = 232 THEN
            tanh_f := 232;
        ELSIF x = 233 THEN
            tanh_f := 233;
        ELSIF x = 234 THEN
            tanh_f := 234;
        ELSIF x = 235 THEN
            tanh_f := 235;
        ELSIF x = 236 THEN
            tanh_f := 236;
        ELSIF x = 237 THEN
            tanh_f := 237;
        ELSIF x = 238 THEN
            tanh_f := 238;
        ELSIF x = 239 THEN
            tanh_f := 239;
        ELSIF x = 240 THEN
            tanh_f := 240;
        ELSIF x = 241 THEN
            tanh_f := 241;
        ELSIF x = 242 THEN
            tanh_f := 242;
        ELSIF x = 243 THEN
            tanh_f := 243;
        ELSIF x = 244 THEN
            tanh_f := 244;
        ELSIF x = 245 THEN
            tanh_f := 245;
        ELSIF x = 246 THEN
            tanh_f := 246;
        ELSIF x = 247 THEN
            tanh_f := 247;
        ELSIF x = 248 THEN
            tanh_f := 248;
        ELSIF x = 249 THEN
            tanh_f := 249;
        ELSIF x = 250 THEN
            tanh_f := 250;
        ELSIF x = 251 THEN
            tanh_f := 251;
        ELSIF x = 252 THEN
            tanh_f := 252;
        ELSIF x = 253 THEN
            tanh_f := 253;
        ELSIF x = 254 THEN
            tanh_f := 254;
        ELSIF x = 255 THEN
            tanh_f := 255;
        ELSIF x = 256 THEN
            tanh_f := 255;
        ELSIF x = 257 THEN
            tanh_f := 256;
        ELSIF x = 258 THEN
            tanh_f := 257;
        ELSIF x = 259 THEN
            tanh_f := 258;
        ELSIF x = 260 THEN
            tanh_f := 259;
        ELSIF x = 261 THEN
            tanh_f := 260;
        ELSIF x = 262 THEN
            tanh_f := 261;
        ELSIF x = 263 THEN
            tanh_f := 262;
        ELSIF x = 264 THEN
            tanh_f := 263;
        ELSIF x = 265 THEN
            tanh_f := 264;
        ELSIF x = 266 THEN
            tanh_f := 265;
        ELSIF x = 267 THEN
            tanh_f := 266;
        ELSIF x = 268 THEN
            tanh_f := 267;
        ELSIF x = 269 THEN
            tanh_f := 268;
        ELSIF x = 270 THEN
            tanh_f := 269;
        ELSIF x = 271 THEN
            tanh_f := 270;
        ELSIF x = 272 THEN
            tanh_f := 270;
        ELSIF x = 273 THEN
            tanh_f := 271;
        ELSIF x = 274 THEN
            tanh_f := 272;
        ELSIF x = 275 THEN
            tanh_f := 273;
        ELSIF x = 276 THEN
            tanh_f := 274;
        ELSIF x = 277 THEN
            tanh_f := 275;
        ELSIF x = 278 THEN
            tanh_f := 276;
        ELSIF x = 279 THEN
            tanh_f := 277;
        ELSIF x = 280 THEN
            tanh_f := 278;
        ELSIF x = 281 THEN
            tanh_f := 279;
        ELSIF x = 282 THEN
            tanh_f := 280;
        ELSIF x = 283 THEN
            tanh_f := 281;
        ELSIF x = 284 THEN
            tanh_f := 282;
        ELSIF x = 285 THEN
            tanh_f := 283;
        ELSIF x = 286 THEN
            tanh_f := 284;
        ELSIF x = 287 THEN
            tanh_f := 285;
        ELSIF x = 288 THEN
            tanh_f := 286;
        ELSIF x = 289 THEN
            tanh_f := 287;
        ELSIF x = 290 THEN
            tanh_f := 288;
        ELSIF x = 291 THEN
            tanh_f := 289;
        ELSIF x = 292 THEN
            tanh_f := 290;
        ELSIF x = 293 THEN
            tanh_f := 291;
        ELSIF x = 294 THEN
            tanh_f := 292;
        ELSIF x = 295 THEN
            tanh_f := 293;
        ELSIF x = 296 THEN
            tanh_f := 294;
        ELSIF x = 297 THEN
            tanh_f := 295;
        ELSIF x = 298 THEN
            tanh_f := 296;
        ELSIF x = 299 THEN
            tanh_f := 297;
        ELSIF x = 300 THEN
            tanh_f := 298;
        ELSIF x = 301 THEN
            tanh_f := 299;
        ELSIF x = 302 THEN
            tanh_f := 299;
        ELSIF x = 303 THEN
            tanh_f := 300;
        ELSIF x = 304 THEN
            tanh_f := 301;
        ELSIF x = 305 THEN
            tanh_f := 302;
        ELSIF x = 306 THEN
            tanh_f := 303;
        ELSIF x = 307 THEN
            tanh_f := 304;
        ELSIF x = 308 THEN
            tanh_f := 305;
        ELSIF x = 309 THEN
            tanh_f := 306;
        ELSIF x = 310 THEN
            tanh_f := 307;
        ELSIF x = 311 THEN
            tanh_f := 308;
        ELSIF x = 312 THEN
            tanh_f := 309;
        ELSIF x = 313 THEN
            tanh_f := 310;
        ELSIF x = 314 THEN
            tanh_f := 311;
        ELSIF x = 315 THEN
            tanh_f := 312;
        ELSIF x = 316 THEN
            tanh_f := 313;
        ELSIF x = 317 THEN
            tanh_f := 314;
        ELSIF x = 318 THEN
            tanh_f := 315;
        ELSIF x = 319 THEN
            tanh_f := 316;
        ELSIF x = 320 THEN
            tanh_f := 317;
        ELSIF x = 321 THEN
            tanh_f := 318;
        ELSIF x = 322 THEN
            tanh_f := 319;
        ELSIF x = 323 THEN
            tanh_f := 320;
        ELSIF x = 324 THEN
            tanh_f := 321;
        ELSIF x = 325 THEN
            tanh_f := 322;
        ELSIF x = 326 THEN
            tanh_f := 323;
        ELSIF x = 327 THEN
            tanh_f := 324;
        ELSIF x = 328 THEN
            tanh_f := 325;
        ELSIF x = 329 THEN
            tanh_f := 326;
        ELSIF x = 330 THEN
            tanh_f := 327;
        ELSIF x = 331 THEN
            tanh_f := 328;
        ELSIF x = 332 THEN
            tanh_f := 328;
        ELSIF x = 333 THEN
            tanh_f := 329;
        ELSIF x = 334 THEN
            tanh_f := 330;
        ELSIF x = 335 THEN
            tanh_f := 331;
        ELSIF x = 336 THEN
            tanh_f := 332;
        ELSIF x = 337 THEN
            tanh_f := 333;
        ELSIF x = 338 THEN
            tanh_f := 334;
        ELSIF x = 339 THEN
            tanh_f := 335;
        ELSIF x = 340 THEN
            tanh_f := 336;
        ELSIF x = 341 THEN
            tanh_f := 337;
        ELSIF x = 342 THEN
            tanh_f := 338;
        ELSIF x = 343 THEN
            tanh_f := 339;
        ELSIF x = 344 THEN
            tanh_f := 340;
        ELSIF x = 345 THEN
            tanh_f := 341;
        ELSIF x = 346 THEN
            tanh_f := 342;
        ELSIF x = 347 THEN
            tanh_f := 343;
        ELSIF x = 348 THEN
            tanh_f := 344;
        ELSIF x = 349 THEN
            tanh_f := 345;
        ELSIF x = 350 THEN
            tanh_f := 346;
        ELSIF x = 351 THEN
            tanh_f := 347;
        ELSIF x = 352 THEN
            tanh_f := 348;
        ELSIF x = 353 THEN
            tanh_f := 349;
        ELSIF x = 354 THEN
            tanh_f := 350;
        ELSIF x = 355 THEN
            tanh_f := 351;
        ELSIF x = 356 THEN
            tanh_f := 352;
        ELSIF x = 357 THEN
            tanh_f := 353;
        ELSIF x = 358 THEN
            tanh_f := 354;
        ELSIF x = 359 THEN
            tanh_f := 355;
        ELSIF x = 360 THEN
            tanh_f := 356;
        ELSIF x = 361 THEN
            tanh_f := 357;
        ELSIF x = 362 THEN
            tanh_f := 357;
        ELSIF x = 363 THEN
            tanh_f := 358;
        ELSIF x = 364 THEN
            tanh_f := 359;
        ELSIF x = 365 THEN
            tanh_f := 360;
        ELSIF x = 366 THEN
            tanh_f := 361;
        ELSIF x = 367 THEN
            tanh_f := 362;
        ELSIF x = 368 THEN
            tanh_f := 363;
        ELSIF x = 369 THEN
            tanh_f := 364;
        ELSIF x = 370 THEN
            tanh_f := 365;
        ELSIF x = 371 THEN
            tanh_f := 366;
        ELSIF x = 372 THEN
            tanh_f := 367;
        ELSIF x = 373 THEN
            tanh_f := 368;
        ELSIF x = 374 THEN
            tanh_f := 369;
        ELSIF x = 375 THEN
            tanh_f := 370;
        ELSIF x = 376 THEN
            tanh_f := 371;
        ELSIF x = 377 THEN
            tanh_f := 372;
        ELSIF x = 378 THEN
            tanh_f := 373;
        ELSIF x = 379 THEN
            tanh_f := 374;
        ELSIF x = 380 THEN
            tanh_f := 375;
        ELSIF x = 381 THEN
            tanh_f := 376;
        ELSIF x = 382 THEN
            tanh_f := 377;
        ELSIF x = 383 THEN
            tanh_f := 378;
        ELSIF x = 384 THEN
            tanh_f := 379;
        ELSIF x = 385 THEN
            tanh_f := 380;
        ELSIF x = 386 THEN
            tanh_f := 381;
        ELSIF x = 387 THEN
            tanh_f := 382;
        ELSIF x = 388 THEN
            tanh_f := 383;
        ELSIF x = 389 THEN
            tanh_f := 384;
        ELSIF x = 390 THEN
            tanh_f := 385;
        ELSIF x = 391 THEN
            tanh_f := 386;
        ELSIF x = 392 THEN
            tanh_f := 386;
        ELSIF x = 393 THEN
            tanh_f := 387;
        ELSIF x = 394 THEN
            tanh_f := 388;
        ELSIF x = 395 THEN
            tanh_f := 389;
        ELSIF x = 396 THEN
            tanh_f := 390;
        ELSIF x = 397 THEN
            tanh_f := 391;
        ELSIF x = 398 THEN
            tanh_f := 392;
        ELSIF x = 399 THEN
            tanh_f := 393;
        ELSIF x = 400 THEN
            tanh_f := 394;
        ELSIF x = 401 THEN
            tanh_f := 395;
        ELSIF x = 402 THEN
            tanh_f := 396;
        ELSIF x = 403 THEN
            tanh_f := 397;
        ELSIF x = 404 THEN
            tanh_f := 398;
        ELSIF x = 405 THEN
            tanh_f := 399;
        ELSIF x = 406 THEN
            tanh_f := 400;
        ELSIF x = 407 THEN
            tanh_f := 401;
        ELSIF x = 408 THEN
            tanh_f := 402;
        ELSIF x = 409 THEN
            tanh_f := 403;
        ELSIF x = 410 THEN
            tanh_f := 404;
        ELSIF x = 411 THEN
            tanh_f := 405;
        ELSIF x = 412 THEN
            tanh_f := 406;
        ELSIF x = 413 THEN
            tanh_f := 407;
        ELSIF x = 414 THEN
            tanh_f := 408;
        ELSIF x = 415 THEN
            tanh_f := 409;
        ELSIF x = 416 THEN
            tanh_f := 410;
        ELSIF x = 417 THEN
            tanh_f := 411;
        ELSIF x = 418 THEN
            tanh_f := 412;
        ELSIF x = 419 THEN
            tanh_f := 413;
        ELSIF x = 420 THEN
            tanh_f := 414;
        ELSIF x = 421 THEN
            tanh_f := 415;
        ELSIF x = 422 THEN
            tanh_f := 415;
        ELSIF x = 423 THEN
            tanh_f := 416;
        ELSIF x = 424 THEN
            tanh_f := 417;
        ELSIF x = 425 THEN
            tanh_f := 418;
        ELSIF x = 426 THEN
            tanh_f := 419;
        ELSIF x = 427 THEN
            tanh_f := 420;
        ELSIF x = 428 THEN
            tanh_f := 421;
        ELSIF x = 429 THEN
            tanh_f := 422;
        ELSIF x = 430 THEN
            tanh_f := 423;
        ELSIF x = 431 THEN
            tanh_f := 424;
        ELSIF x = 432 THEN
            tanh_f := 425;
        ELSIF x = 433 THEN
            tanh_f := 426;
        ELSIF x = 434 THEN
            tanh_f := 427;
        ELSIF x = 435 THEN
            tanh_f := 428;
        ELSIF x = 436 THEN
            tanh_f := 429;
        ELSIF x = 437 THEN
            tanh_f := 430;
        ELSIF x = 438 THEN
            tanh_f := 431;
        ELSIF x = 439 THEN
            tanh_f := 432;
        ELSIF x = 440 THEN
            tanh_f := 433;
        ELSIF x = 441 THEN
            tanh_f := 434;
        ELSIF x = 442 THEN
            tanh_f := 435;
        ELSIF x = 443 THEN
            tanh_f := 436;
        ELSIF x = 444 THEN
            tanh_f := 437;
        ELSIF x = 445 THEN
            tanh_f := 438;
        ELSIF x = 446 THEN
            tanh_f := 439;
        ELSIF x = 447 THEN
            tanh_f := 440;
        ELSIF x = 448 THEN
            tanh_f := 441;
        ELSIF x = 449 THEN
            tanh_f := 442;
        ELSIF x = 450 THEN
            tanh_f := 443;
        ELSIF x = 451 THEN
            tanh_f := 444;
        ELSIF x = 452 THEN
            tanh_f := 444;
        ELSIF x = 453 THEN
            tanh_f := 445;
        ELSIF x = 454 THEN
            tanh_f := 446;
        ELSIF x = 455 THEN
            tanh_f := 447;
        ELSIF x = 456 THEN
            tanh_f := 448;
        ELSIF x = 457 THEN
            tanh_f := 449;
        ELSIF x = 458 THEN
            tanh_f := 450;
        ELSIF x = 459 THEN
            tanh_f := 451;
        ELSIF x = 460 THEN
            tanh_f := 452;
        ELSIF x = 461 THEN
            tanh_f := 453;
        ELSIF x = 462 THEN
            tanh_f := 454;
        ELSIF x = 463 THEN
            tanh_f := 455;
        ELSIF x = 464 THEN
            tanh_f := 456;
        ELSIF x = 465 THEN
            tanh_f := 457;
        ELSIF x = 466 THEN
            tanh_f := 458;
        ELSIF x = 467 THEN
            tanh_f := 459;
        ELSIF x = 468 THEN
            tanh_f := 460;
        ELSIF x = 469 THEN
            tanh_f := 461;
        ELSIF x = 470 THEN
            tanh_f := 462;
        ELSIF x = 471 THEN
            tanh_f := 463;
        ELSIF x = 472 THEN
            tanh_f := 464;
        ELSIF x = 473 THEN
            tanh_f := 465;
        ELSIF x = 474 THEN
            tanh_f := 466;
        ELSIF x = 475 THEN
            tanh_f := 467;
        ELSIF x = 476 THEN
            tanh_f := 468;
        ELSIF x = 477 THEN
            tanh_f := 469;
        ELSIF x = 478 THEN
            tanh_f := 470;
        ELSIF x = 479 THEN
            tanh_f := 471;
        ELSIF x = 480 THEN
            tanh_f := 472;
        ELSIF x = 481 THEN
            tanh_f := 473;
        ELSIF x = 482 THEN
            tanh_f := 473;
        ELSIF x = 483 THEN
            tanh_f := 474;
        ELSIF x = 484 THEN
            tanh_f := 475;
        ELSIF x = 485 THEN
            tanh_f := 476;
        ELSIF x = 486 THEN
            tanh_f := 477;
        ELSIF x = 487 THEN
            tanh_f := 478;
        ELSIF x = 488 THEN
            tanh_f := 479;
        ELSIF x = 489 THEN
            tanh_f := 480;
        ELSIF x = 490 THEN
            tanh_f := 481;
        ELSIF x = 491 THEN
            tanh_f := 482;
        ELSIF x = 492 THEN
            tanh_f := 483;
        ELSIF x = 493 THEN
            tanh_f := 484;
        ELSIF x = 494 THEN
            tanh_f := 485;
        ELSIF x = 495 THEN
            tanh_f := 486;
        ELSIF x = 496 THEN
            tanh_f := 487;
        ELSIF x = 497 THEN
            tanh_f := 488;
        ELSIF x = 498 THEN
            tanh_f := 489;
        ELSIF x = 499 THEN
            tanh_f := 490;
        ELSIF x = 500 THEN
            tanh_f := 491;
        ELSIF x = 501 THEN
            tanh_f := 492;
        ELSIF x = 502 THEN
            tanh_f := 493;
        ELSIF x = 503 THEN
            tanh_f := 494;
        ELSIF x = 504 THEN
            tanh_f := 495;
        ELSIF x = 505 THEN
            tanh_f := 496;
        ELSIF x = 506 THEN
            tanh_f := 497;
        ELSIF x = 507 THEN
            tanh_f := 498;
        ELSIF x = 508 THEN
            tanh_f := 499;
        ELSIF x = 509 THEN
            tanh_f := 500;
        ELSIF x = 510 THEN
            tanh_f := 501;
        ELSIF x = 511 THEN
            tanh_f := 502;
        ELSIF x = 512 THEN
            tanh_f := 503;
        ELSIF x = 513 THEN
            tanh_f := 503;
        ELSIF x = 514 THEN
            tanh_f := 504;
        ELSIF x = 515 THEN
            tanh_f := 505;
        ELSIF x = 516 THEN
            tanh_f := 506;
        ELSIF x = 517 THEN
            tanh_f := 507;
        ELSIF x = 518 THEN
            tanh_f := 508;
        ELSIF x = 519 THEN
            tanh_f := 509;
        ELSIF x = 520 THEN
            tanh_f := 510;
        ELSIF x = 521 THEN
            tanh_f := 511;
        ELSIF x = 522 THEN
            tanh_f := 512;
        ELSIF x = 523 THEN
            tanh_f := 512;
        ELSIF x = 524 THEN
            tanh_f := 513;
        ELSIF x = 525 THEN
            tanh_f := 514;
        ELSIF x = 526 THEN
            tanh_f := 515;
        ELSIF x = 527 THEN
            tanh_f := 516;
        ELSIF x = 528 THEN
            tanh_f := 517;
        ELSIF x = 529 THEN
            tanh_f := 518;
        ELSIF x = 530 THEN
            tanh_f := 519;
        ELSIF x = 531 THEN
            tanh_f := 520;
        ELSIF x = 532 THEN
            tanh_f := 521;
        ELSIF x = 533 THEN
            tanh_f := 522;
        ELSIF x = 534 THEN
            tanh_f := 522;
        ELSIF x = 535 THEN
            tanh_f := 523;
        ELSIF x = 536 THEN
            tanh_f := 524;
        ELSIF x = 537 THEN
            tanh_f := 525;
        ELSIF x = 538 THEN
            tanh_f := 526;
        ELSIF x = 539 THEN
            tanh_f := 527;
        ELSIF x = 540 THEN
            tanh_f := 528;
        ELSIF x = 541 THEN
            tanh_f := 529;
        ELSIF x = 542 THEN
            tanh_f := 530;
        ELSIF x = 543 THEN
            tanh_f := 531;
        ELSIF x = 544 THEN
            tanh_f := 532;
        ELSIF x = 545 THEN
            tanh_f := 532;
        ELSIF x = 546 THEN
            tanh_f := 533;
        ELSIF x = 547 THEN
            tanh_f := 534;
        ELSIF x = 548 THEN
            tanh_f := 535;
        ELSIF x = 549 THEN
            tanh_f := 536;
        ELSIF x = 550 THEN
            tanh_f := 537;
        ELSIF x = 551 THEN
            tanh_f := 538;
        ELSIF x = 552 THEN
            tanh_f := 539;
        ELSIF x = 553 THEN
            tanh_f := 540;
        ELSIF x = 554 THEN
            tanh_f := 541;
        ELSIF x = 555 THEN
            tanh_f := 542;
        ELSIF x = 556 THEN
            tanh_f := 542;
        ELSIF x = 557 THEN
            tanh_f := 543;
        ELSIF x = 558 THEN
            tanh_f := 544;
        ELSIF x = 559 THEN
            tanh_f := 545;
        ELSIF x = 560 THEN
            tanh_f := 546;
        ELSIF x = 561 THEN
            tanh_f := 547;
        ELSIF x = 562 THEN
            tanh_f := 548;
        ELSIF x = 563 THEN
            tanh_f := 549;
        ELSIF x = 564 THEN
            tanh_f := 550;
        ELSIF x = 565 THEN
            tanh_f := 551;
        ELSIF x = 566 THEN
            tanh_f := 552;
        ELSIF x = 567 THEN
            tanh_f := 552;
        ELSIF x = 568 THEN
            tanh_f := 553;
        ELSIF x = 569 THEN
            tanh_f := 554;
        ELSIF x = 570 THEN
            tanh_f := 555;
        ELSIF x = 571 THEN
            tanh_f := 556;
        ELSIF x = 572 THEN
            tanh_f := 557;
        ELSIF x = 573 THEN
            tanh_f := 558;
        ELSIF x = 574 THEN
            tanh_f := 559;
        ELSIF x = 575 THEN
            tanh_f := 560;
        ELSIF x = 576 THEN
            tanh_f := 561;
        ELSIF x = 577 THEN
            tanh_f := 562;
        ELSIF x = 578 THEN
            tanh_f := 562;
        ELSIF x = 579 THEN
            tanh_f := 563;
        ELSIF x = 580 THEN
            tanh_f := 564;
        ELSIF x = 581 THEN
            tanh_f := 565;
        ELSIF x = 582 THEN
            tanh_f := 566;
        ELSIF x = 583 THEN
            tanh_f := 567;
        ELSIF x = 584 THEN
            tanh_f := 568;
        ELSIF x = 585 THEN
            tanh_f := 569;
        ELSIF x = 586 THEN
            tanh_f := 570;
        ELSIF x = 587 THEN
            tanh_f := 571;
        ELSIF x = 588 THEN
            tanh_f := 572;
        ELSIF x = 589 THEN
            tanh_f := 572;
        ELSIF x = 590 THEN
            tanh_f := 573;
        ELSIF x = 591 THEN
            tanh_f := 574;
        ELSIF x = 592 THEN
            tanh_f := 575;
        ELSIF x = 593 THEN
            tanh_f := 576;
        ELSIF x = 594 THEN
            tanh_f := 577;
        ELSIF x = 595 THEN
            tanh_f := 578;
        ELSIF x = 596 THEN
            tanh_f := 579;
        ELSIF x = 597 THEN
            tanh_f := 580;
        ELSIF x = 598 THEN
            tanh_f := 581;
        ELSIF x = 599 THEN
            tanh_f := 582;
        ELSIF x = 600 THEN
            tanh_f := 582;
        ELSIF x = 601 THEN
            tanh_f := 583;
        ELSIF x = 602 THEN
            tanh_f := 584;
        ELSIF x = 603 THEN
            tanh_f := 585;
        ELSIF x = 604 THEN
            tanh_f := 586;
        ELSIF x = 605 THEN
            tanh_f := 587;
        ELSIF x = 606 THEN
            tanh_f := 588;
        ELSIF x = 607 THEN
            tanh_f := 589;
        ELSIF x = 608 THEN
            tanh_f := 590;
        ELSIF x = 609 THEN
            tanh_f := 591;
        ELSIF x = 610 THEN
            tanh_f := 592;
        ELSIF x = 611 THEN
            tanh_f := 592;
        ELSIF x = 612 THEN
            tanh_f := 593;
        ELSIF x = 613 THEN
            tanh_f := 594;
        ELSIF x = 614 THEN
            tanh_f := 595;
        ELSIF x = 615 THEN
            tanh_f := 596;
        ELSIF x = 616 THEN
            tanh_f := 597;
        ELSIF x = 617 THEN
            tanh_f := 598;
        ELSIF x = 618 THEN
            tanh_f := 599;
        ELSIF x = 619 THEN
            tanh_f := 600;
        ELSIF x = 620 THEN
            tanh_f := 601;
        ELSIF x = 621 THEN
            tanh_f := 601;
        ELSIF x = 622 THEN
            tanh_f := 602;
        ELSIF x = 623 THEN
            tanh_f := 603;
        ELSIF x = 624 THEN
            tanh_f := 604;
        ELSIF x = 625 THEN
            tanh_f := 605;
        ELSIF x = 626 THEN
            tanh_f := 606;
        ELSIF x = 627 THEN
            tanh_f := 607;
        ELSIF x = 628 THEN
            tanh_f := 608;
        ELSIF x = 629 THEN
            tanh_f := 609;
        ELSIF x = 630 THEN
            tanh_f := 610;
        ELSIF x = 631 THEN
            tanh_f := 611;
        ELSIF x = 632 THEN
            tanh_f := 611;
        ELSIF x = 633 THEN
            tanh_f := 612;
        ELSIF x = 634 THEN
            tanh_f := 613;
        ELSIF x = 635 THEN
            tanh_f := 614;
        ELSIF x = 636 THEN
            tanh_f := 615;
        ELSIF x = 637 THEN
            tanh_f := 616;
        ELSIF x = 638 THEN
            tanh_f := 617;
        ELSIF x = 639 THEN
            tanh_f := 618;
        ELSIF x = 640 THEN
            tanh_f := 619;
        ELSIF x = 641 THEN
            tanh_f := 620;
        ELSIF x = 642 THEN
            tanh_f := 621;
        ELSIF x = 643 THEN
            tanh_f := 621;
        ELSIF x = 644 THEN
            tanh_f := 622;
        ELSIF x = 645 THEN
            tanh_f := 623;
        ELSIF x = 646 THEN
            tanh_f := 624;
        ELSIF x = 647 THEN
            tanh_f := 625;
        ELSIF x = 648 THEN
            tanh_f := 626;
        ELSIF x = 649 THEN
            tanh_f := 627;
        ELSIF x = 650 THEN
            tanh_f := 628;
        ELSIF x = 651 THEN
            tanh_f := 629;
        ELSIF x = 652 THEN
            tanh_f := 630;
        ELSIF x = 653 THEN
            tanh_f := 631;
        ELSIF x = 654 THEN
            tanh_f := 631;
        ELSIF x = 655 THEN
            tanh_f := 632;
        ELSIF x = 656 THEN
            tanh_f := 633;
        ELSIF x = 657 THEN
            tanh_f := 634;
        ELSIF x = 658 THEN
            tanh_f := 635;
        ELSIF x = 659 THEN
            tanh_f := 636;
        ELSIF x = 660 THEN
            tanh_f := 637;
        ELSIF x = 661 THEN
            tanh_f := 638;
        ELSIF x = 662 THEN
            tanh_f := 639;
        ELSIF x = 663 THEN
            tanh_f := 640;
        ELSIF x = 664 THEN
            tanh_f := 641;
        ELSIF x = 665 THEN
            tanh_f := 641;
        ELSIF x = 666 THEN
            tanh_f := 642;
        ELSIF x = 667 THEN
            tanh_f := 643;
        ELSIF x = 668 THEN
            tanh_f := 644;
        ELSIF x = 669 THEN
            tanh_f := 645;
        ELSIF x = 670 THEN
            tanh_f := 646;
        ELSIF x = 671 THEN
            tanh_f := 647;
        ELSIF x = 672 THEN
            tanh_f := 648;
        ELSIF x = 673 THEN
            tanh_f := 649;
        ELSIF x = 674 THEN
            tanh_f := 650;
        ELSIF x = 675 THEN
            tanh_f := 651;
        ELSIF x = 676 THEN
            tanh_f := 651;
        ELSIF x = 677 THEN
            tanh_f := 652;
        ELSIF x = 678 THEN
            tanh_f := 653;
        ELSIF x = 679 THEN
            tanh_f := 654;
        ELSIF x = 680 THEN
            tanh_f := 655;
        ELSIF x = 681 THEN
            tanh_f := 656;
        ELSIF x = 682 THEN
            tanh_f := 657;
        ELSIF x = 683 THEN
            tanh_f := 658;
        ELSIF x = 684 THEN
            tanh_f := 659;
        ELSIF x = 685 THEN
            tanh_f := 660;
        ELSIF x = 686 THEN
            tanh_f := 661;
        ELSIF x = 687 THEN
            tanh_f := 661;
        ELSIF x = 688 THEN
            tanh_f := 662;
        ELSIF x = 689 THEN
            tanh_f := 663;
        ELSIF x = 690 THEN
            tanh_f := 664;
        ELSIF x = 691 THEN
            tanh_f := 665;
        ELSIF x = 692 THEN
            tanh_f := 666;
        ELSIF x = 693 THEN
            tanh_f := 667;
        ELSIF x = 694 THEN
            tanh_f := 668;
        ELSIF x = 695 THEN
            tanh_f := 669;
        ELSIF x = 696 THEN
            tanh_f := 670;
        ELSIF x = 697 THEN
            tanh_f := 671;
        ELSIF x = 698 THEN
            tanh_f := 671;
        ELSIF x = 699 THEN
            tanh_f := 672;
        ELSIF x = 700 THEN
            tanh_f := 673;
        ELSIF x = 701 THEN
            tanh_f := 674;
        ELSIF x = 702 THEN
            tanh_f := 675;
        ELSIF x = 703 THEN
            tanh_f := 676;
        ELSIF x = 704 THEN
            tanh_f := 677;
        ELSIF x = 705 THEN
            tanh_f := 678;
        ELSIF x = 706 THEN
            tanh_f := 679;
        ELSIF x = 707 THEN
            tanh_f := 680;
        ELSIF x = 708 THEN
            tanh_f := 681;
        ELSIF x = 709 THEN
            tanh_f := 681;
        ELSIF x = 710 THEN
            tanh_f := 682;
        ELSIF x = 711 THEN
            tanh_f := 683;
        ELSIF x = 712 THEN
            tanh_f := 684;
        ELSIF x = 713 THEN
            tanh_f := 685;
        ELSIF x = 714 THEN
            tanh_f := 686;
        ELSIF x = 715 THEN
            tanh_f := 687;
        ELSIF x = 716 THEN
            tanh_f := 688;
        ELSIF x = 717 THEN
            tanh_f := 689;
        ELSIF x = 718 THEN
            tanh_f := 690;
        ELSIF x = 719 THEN
            tanh_f := 690;
        ELSIF x = 720 THEN
            tanh_f := 691;
        ELSIF x = 721 THEN
            tanh_f := 692;
        ELSIF x = 722 THEN
            tanh_f := 693;
        ELSIF x = 723 THEN
            tanh_f := 694;
        ELSIF x = 724 THEN
            tanh_f := 695;
        ELSIF x = 725 THEN
            tanh_f := 696;
        ELSIF x = 726 THEN
            tanh_f := 697;
        ELSIF x = 727 THEN
            tanh_f := 698;
        ELSIF x = 728 THEN
            tanh_f := 699;
        ELSIF x = 729 THEN
            tanh_f := 700;
        ELSIF x = 730 THEN
            tanh_f := 700;
        ELSIF x = 731 THEN
            tanh_f := 701;
        ELSIF x = 732 THEN
            tanh_f := 702;
        ELSIF x = 733 THEN
            tanh_f := 703;
        ELSIF x = 734 THEN
            tanh_f := 704;
        ELSIF x = 735 THEN
            tanh_f := 705;
        ELSIF x = 736 THEN
            tanh_f := 706;
        ELSIF x = 737 THEN
            tanh_f := 707;
        ELSIF x = 738 THEN
            tanh_f := 708;
        ELSIF x = 739 THEN
            tanh_f := 709;
        ELSIF x = 740 THEN
            tanh_f := 710;
        ELSIF x = 741 THEN
            tanh_f := 710;
        ELSIF x = 742 THEN
            tanh_f := 711;
        ELSIF x = 743 THEN
            tanh_f := 712;
        ELSIF x = 744 THEN
            tanh_f := 713;
        ELSIF x = 745 THEN
            tanh_f := 714;
        ELSIF x = 746 THEN
            tanh_f := 715;
        ELSIF x = 747 THEN
            tanh_f := 716;
        ELSIF x = 748 THEN
            tanh_f := 717;
        ELSIF x = 749 THEN
            tanh_f := 718;
        ELSIF x = 750 THEN
            tanh_f := 719;
        ELSIF x = 751 THEN
            tanh_f := 720;
        ELSIF x = 752 THEN
            tanh_f := 720;
        ELSIF x = 753 THEN
            tanh_f := 721;
        ELSIF x = 754 THEN
            tanh_f := 722;
        ELSIF x = 755 THEN
            tanh_f := 723;
        ELSIF x = 756 THEN
            tanh_f := 724;
        ELSIF x = 757 THEN
            tanh_f := 725;
        ELSIF x = 758 THEN
            tanh_f := 726;
        ELSIF x = 759 THEN
            tanh_f := 727;
        ELSIF x = 760 THEN
            tanh_f := 728;
        ELSIF x = 761 THEN
            tanh_f := 729;
        ELSIF x = 762 THEN
            tanh_f := 730;
        ELSIF x = 763 THEN
            tanh_f := 730;
        ELSIF x = 764 THEN
            tanh_f := 731;
        ELSIF x = 765 THEN
            tanh_f := 732;
        ELSIF x = 766 THEN
            tanh_f := 733;
        ELSIF x = 767 THEN
            tanh_f := 734;
        ELSIF x = 768 THEN
            tanh_f := 736;
        ELSIF x = 769 THEN
            tanh_f := 736;
        ELSIF x = 770 THEN
            tanh_f := 737;
        ELSIF x = 771 THEN
            tanh_f := 738;
        ELSIF x = 772 THEN
            tanh_f := 739;
        ELSIF x = 773 THEN
            tanh_f := 740;
        ELSIF x = 774 THEN
            tanh_f := 740;
        ELSIF x = 775 THEN
            tanh_f := 741;
        ELSIF x = 776 THEN
            tanh_f := 742;
        ELSIF x = 777 THEN
            tanh_f := 743;
        ELSIF x = 778 THEN
            tanh_f := 744;
        ELSIF x = 779 THEN
            tanh_f := 745;
        ELSIF x = 780 THEN
            tanh_f := 745;
        ELSIF x = 781 THEN
            tanh_f := 746;
        ELSIF x = 782 THEN
            tanh_f := 747;
        ELSIF x = 783 THEN
            tanh_f := 748;
        ELSIF x = 784 THEN
            tanh_f := 749;
        ELSIF x = 785 THEN
            tanh_f := 750;
        ELSIF x = 786 THEN
            tanh_f := 750;
        ELSIF x = 787 THEN
            tanh_f := 751;
        ELSIF x = 788 THEN
            tanh_f := 752;
        ELSIF x = 789 THEN
            tanh_f := 753;
        ELSIF x = 790 THEN
            tanh_f := 754;
        ELSIF x = 791 THEN
            tanh_f := 755;
        ELSIF x = 792 THEN
            tanh_f := 755;
        ELSIF x = 793 THEN
            tanh_f := 756;
        ELSIF x = 794 THEN
            tanh_f := 757;
        ELSIF x = 795 THEN
            tanh_f := 758;
        ELSIF x = 796 THEN
            tanh_f := 759;
        ELSIF x = 797 THEN
            tanh_f := 760;
        ELSIF x = 798 THEN
            tanh_f := 760;
        ELSIF x = 799 THEN
            tanh_f := 761;
        ELSIF x = 800 THEN
            tanh_f := 762;
        ELSIF x = 801 THEN
            tanh_f := 763;
        ELSIF x = 802 THEN
            tanh_f := 764;
        ELSIF x = 803 THEN
            tanh_f := 764;
        ELSIF x = 804 THEN
            tanh_f := 765;
        ELSIF x = 805 THEN
            tanh_f := 766;
        ELSIF x = 806 THEN
            tanh_f := 767;
        ELSIF x = 807 THEN
            tanh_f := 768;
        ELSIF x = 808 THEN
            tanh_f := 769;
        ELSIF x = 809 THEN
            tanh_f := 769;
        ELSIF x = 810 THEN
            tanh_f := 770;
        ELSIF x = 811 THEN
            tanh_f := 771;
        ELSIF x = 812 THEN
            tanh_f := 772;
        ELSIF x = 813 THEN
            tanh_f := 773;
        ELSIF x = 814 THEN
            tanh_f := 774;
        ELSIF x = 815 THEN
            tanh_f := 774;
        ELSIF x = 816 THEN
            tanh_f := 775;
        ELSIF x = 817 THEN
            tanh_f := 776;
        ELSIF x = 818 THEN
            tanh_f := 777;
        ELSIF x = 819 THEN
            tanh_f := 778;
        ELSIF x = 820 THEN
            tanh_f := 779;
        ELSIF x = 821 THEN
            tanh_f := 779;
        ELSIF x = 822 THEN
            tanh_f := 780;
        ELSIF x = 823 THEN
            tanh_f := 781;
        ELSIF x = 824 THEN
            tanh_f := 782;
        ELSIF x = 825 THEN
            tanh_f := 783;
        ELSIF x = 826 THEN
            tanh_f := 784;
        ELSIF x = 827 THEN
            tanh_f := 784;
        ELSIF x = 828 THEN
            tanh_f := 785;
        ELSIF x = 829 THEN
            tanh_f := 786;
        ELSIF x = 830 THEN
            tanh_f := 787;
        ELSIF x = 831 THEN
            tanh_f := 788;
        ELSIF x = 832 THEN
            tanh_f := 789;
        ELSIF x = 833 THEN
            tanh_f := 789;
        ELSIF x = 834 THEN
            tanh_f := 790;
        ELSIF x = 835 THEN
            tanh_f := 791;
        ELSIF x = 836 THEN
            tanh_f := 792;
        ELSIF x = 837 THEN
            tanh_f := 793;
        ELSIF x = 838 THEN
            tanh_f := 793;
        ELSIF x = 839 THEN
            tanh_f := 794;
        ELSIF x = 840 THEN
            tanh_f := 795;
        ELSIF x = 841 THEN
            tanh_f := 796;
        ELSIF x = 842 THEN
            tanh_f := 797;
        ELSIF x = 843 THEN
            tanh_f := 798;
        ELSIF x = 844 THEN
            tanh_f := 798;
        ELSIF x = 845 THEN
            tanh_f := 799;
        ELSIF x = 846 THEN
            tanh_f := 800;
        ELSIF x = 847 THEN
            tanh_f := 801;
        ELSIF x = 848 THEN
            tanh_f := 802;
        ELSIF x = 849 THEN
            tanh_f := 803;
        ELSIF x = 850 THEN
            tanh_f := 803;
        ELSIF x = 851 THEN
            tanh_f := 804;
        ELSIF x = 852 THEN
            tanh_f := 805;
        ELSIF x = 853 THEN
            tanh_f := 806;
        ELSIF x = 854 THEN
            tanh_f := 807;
        ELSIF x = 855 THEN
            tanh_f := 808;
        ELSIF x = 856 THEN
            tanh_f := 808;
        ELSIF x = 857 THEN
            tanh_f := 809;
        ELSIF x = 858 THEN
            tanh_f := 810;
        ELSIF x = 859 THEN
            tanh_f := 811;
        ELSIF x = 860 THEN
            tanh_f := 812;
        ELSIF x = 861 THEN
            tanh_f := 813;
        ELSIF x = 862 THEN
            tanh_f := 813;
        ELSIF x = 863 THEN
            tanh_f := 814;
        ELSIF x = 864 THEN
            tanh_f := 815;
        ELSIF x = 865 THEN
            tanh_f := 816;
        ELSIF x = 866 THEN
            tanh_f := 817;
        ELSIF x = 867 THEN
            tanh_f := 817;
        ELSIF x = 868 THEN
            tanh_f := 818;
        ELSIF x = 869 THEN
            tanh_f := 819;
        ELSIF x = 870 THEN
            tanh_f := 820;
        ELSIF x = 871 THEN
            tanh_f := 821;
        ELSIF x = 872 THEN
            tanh_f := 822;
        ELSIF x = 873 THEN
            tanh_f := 822;
        ELSIF x = 874 THEN
            tanh_f := 823;
        ELSIF x = 875 THEN
            tanh_f := 824;
        ELSIF x = 876 THEN
            tanh_f := 825;
        ELSIF x = 877 THEN
            tanh_f := 826;
        ELSIF x = 878 THEN
            tanh_f := 827;
        ELSIF x = 879 THEN
            tanh_f := 827;
        ELSIF x = 880 THEN
            tanh_f := 828;
        ELSIF x = 881 THEN
            tanh_f := 829;
        ELSIF x = 882 THEN
            tanh_f := 830;
        ELSIF x = 883 THEN
            tanh_f := 831;
        ELSIF x = 884 THEN
            tanh_f := 832;
        ELSIF x = 885 THEN
            tanh_f := 832;
        ELSIF x = 886 THEN
            tanh_f := 833;
        ELSIF x = 887 THEN
            tanh_f := 834;
        ELSIF x = 888 THEN
            tanh_f := 835;
        ELSIF x = 889 THEN
            tanh_f := 836;
        ELSIF x = 890 THEN
            tanh_f := 837;
        ELSIF x = 891 THEN
            tanh_f := 837;
        ELSIF x = 892 THEN
            tanh_f := 838;
        ELSIF x = 893 THEN
            tanh_f := 839;
        ELSIF x = 894 THEN
            tanh_f := 840;
        ELSIF x = 895 THEN
            tanh_f := 841;
        ELSIF x = 896 THEN
            tanh_f := 842;
        ELSIF x = 897 THEN
            tanh_f := 842;
        ELSIF x = 898 THEN
            tanh_f := 843;
        ELSIF x = 899 THEN
            tanh_f := 844;
        ELSIF x = 900 THEN
            tanh_f := 845;
        ELSIF x = 901 THEN
            tanh_f := 846;
        ELSIF x = 902 THEN
            tanh_f := 846;
        ELSIF x = 903 THEN
            tanh_f := 847;
        ELSIF x = 904 THEN
            tanh_f := 848;
        ELSIF x = 905 THEN
            tanh_f := 849;
        ELSIF x = 906 THEN
            tanh_f := 850;
        ELSIF x = 907 THEN
            tanh_f := 851;
        ELSIF x = 908 THEN
            tanh_f := 851;
        ELSIF x = 909 THEN
            tanh_f := 852;
        ELSIF x = 910 THEN
            tanh_f := 853;
        ELSIF x = 911 THEN
            tanh_f := 854;
        ELSIF x = 912 THEN
            tanh_f := 855;
        ELSIF x = 913 THEN
            tanh_f := 856;
        ELSIF x = 914 THEN
            tanh_f := 856;
        ELSIF x = 915 THEN
            tanh_f := 857;
        ELSIF x = 916 THEN
            tanh_f := 858;
        ELSIF x = 917 THEN
            tanh_f := 859;
        ELSIF x = 918 THEN
            tanh_f := 860;
        ELSIF x = 919 THEN
            tanh_f := 861;
        ELSIF x = 920 THEN
            tanh_f := 861;
        ELSIF x = 921 THEN
            tanh_f := 862;
        ELSIF x = 922 THEN
            tanh_f := 863;
        ELSIF x = 923 THEN
            tanh_f := 864;
        ELSIF x = 924 THEN
            tanh_f := 865;
        ELSIF x = 925 THEN
            tanh_f := 866;
        ELSIF x = 926 THEN
            tanh_f := 866;
        ELSIF x = 927 THEN
            tanh_f := 867;
        ELSIF x = 928 THEN
            tanh_f := 868;
        ELSIF x = 929 THEN
            tanh_f := 869;
        ELSIF x = 930 THEN
            tanh_f := 870;
        ELSIF x = 931 THEN
            tanh_f := 870;
        ELSIF x = 932 THEN
            tanh_f := 871;
        ELSIF x = 933 THEN
            tanh_f := 872;
        ELSIF x = 934 THEN
            tanh_f := 873;
        ELSIF x = 935 THEN
            tanh_f := 874;
        ELSIF x = 936 THEN
            tanh_f := 875;
        ELSIF x = 937 THEN
            tanh_f := 875;
        ELSIF x = 938 THEN
            tanh_f := 876;
        ELSIF x = 939 THEN
            tanh_f := 877;
        ELSIF x = 940 THEN
            tanh_f := 878;
        ELSIF x = 941 THEN
            tanh_f := 879;
        ELSIF x = 942 THEN
            tanh_f := 880;
        ELSIF x = 943 THEN
            tanh_f := 880;
        ELSIF x = 944 THEN
            tanh_f := 881;
        ELSIF x = 945 THEN
            tanh_f := 882;
        ELSIF x = 946 THEN
            tanh_f := 883;
        ELSIF x = 947 THEN
            tanh_f := 884;
        ELSIF x = 948 THEN
            tanh_f := 885;
        ELSIF x = 949 THEN
            tanh_f := 885;
        ELSIF x = 950 THEN
            tanh_f := 886;
        ELSIF x = 951 THEN
            tanh_f := 887;
        ELSIF x = 952 THEN
            tanh_f := 888;
        ELSIF x = 953 THEN
            tanh_f := 889;
        ELSIF x = 954 THEN
            tanh_f := 890;
        ELSIF x = 955 THEN
            tanh_f := 890;
        ELSIF x = 956 THEN
            tanh_f := 891;
        ELSIF x = 957 THEN
            tanh_f := 892;
        ELSIF x = 958 THEN
            tanh_f := 893;
        ELSIF x = 959 THEN
            tanh_f := 894;
        ELSIF x = 960 THEN
            tanh_f := 895;
        ELSIF x = 961 THEN
            tanh_f := 895;
        ELSIF x = 962 THEN
            tanh_f := 896;
        ELSIF x = 963 THEN
            tanh_f := 897;
        ELSIF x = 964 THEN
            tanh_f := 898;
        ELSIF x = 965 THEN
            tanh_f := 899;
        ELSIF x = 966 THEN
            tanh_f := 899;
        ELSIF x = 967 THEN
            tanh_f := 900;
        ELSIF x = 968 THEN
            tanh_f := 901;
        ELSIF x = 969 THEN
            tanh_f := 902;
        ELSIF x = 970 THEN
            tanh_f := 903;
        ELSIF x = 971 THEN
            tanh_f := 904;
        ELSIF x = 972 THEN
            tanh_f := 904;
        ELSIF x = 973 THEN
            tanh_f := 905;
        ELSIF x = 974 THEN
            tanh_f := 906;
        ELSIF x = 975 THEN
            tanh_f := 907;
        ELSIF x = 976 THEN
            tanh_f := 908;
        ELSIF x = 977 THEN
            tanh_f := 909;
        ELSIF x = 978 THEN
            tanh_f := 909;
        ELSIF x = 979 THEN
            tanh_f := 910;
        ELSIF x = 980 THEN
            tanh_f := 911;
        ELSIF x = 981 THEN
            tanh_f := 912;
        ELSIF x = 982 THEN
            tanh_f := 913;
        ELSIF x = 983 THEN
            tanh_f := 914;
        ELSIF x = 984 THEN
            tanh_f := 914;
        ELSIF x = 985 THEN
            tanh_f := 915;
        ELSIF x = 986 THEN
            tanh_f := 916;
        ELSIF x = 987 THEN
            tanh_f := 917;
        ELSIF x = 988 THEN
            tanh_f := 918;
        ELSIF x = 989 THEN
            tanh_f := 919;
        ELSIF x = 990 THEN
            tanh_f := 919;
        ELSIF x = 991 THEN
            tanh_f := 920;
        ELSIF x = 992 THEN
            tanh_f := 921;
        ELSIF x = 993 THEN
            tanh_f := 922;
        ELSIF x = 994 THEN
            tanh_f := 923;
        ELSIF x = 995 THEN
            tanh_f := 923;
        ELSIF x = 996 THEN
            tanh_f := 924;
        ELSIF x = 997 THEN
            tanh_f := 925;
        ELSIF x = 998 THEN
            tanh_f := 926;
        ELSIF x = 999 THEN
            tanh_f := 927;
        ELSIF x = 1000 THEN
            tanh_f := 928;
        ELSIF x = 1001 THEN
            tanh_f := 928;
        ELSIF x = 1002 THEN
            tanh_f := 929;
        ELSIF x = 1003 THEN
            tanh_f := 930;
        ELSIF x = 1004 THEN
            tanh_f := 931;
        ELSIF x = 1005 THEN
            tanh_f := 932;
        ELSIF x = 1006 THEN
            tanh_f := 933;
        ELSIF x = 1007 THEN
            tanh_f := 933;
        ELSIF x = 1008 THEN
            tanh_f := 934;
        ELSIF x = 1009 THEN
            tanh_f := 935;
        ELSIF x = 1010 THEN
            tanh_f := 936;
        ELSIF x = 1011 THEN
            tanh_f := 937;
        ELSIF x = 1012 THEN
            tanh_f := 938;
        ELSIF x = 1013 THEN
            tanh_f := 938;
        ELSIF x = 1014 THEN
            tanh_f := 939;
        ELSIF x = 1015 THEN
            tanh_f := 940;
        ELSIF x = 1016 THEN
            tanh_f := 941;
        ELSIF x = 1017 THEN
            tanh_f := 942;
        ELSIF x = 1018 THEN
            tanh_f := 943;
        ELSIF x = 1019 THEN
            tanh_f := 943;
        ELSIF x = 1020 THEN
            tanh_f := 944;
        ELSIF x = 1021 THEN
            tanh_f := 945;
        ELSIF x = 1022 THEN
            tanh_f := 946;
        ELSIF x = 1023 THEN
            tanh_f := 947;
        ELSIF x = 1024 THEN
            tanh_f := 948;
        ELSIF x = 1025 THEN
            tanh_f := 948;
        ELSIF x = 1026 THEN
            tanh_f := 949;
        ELSIF x = 1027 THEN
            tanh_f := 950;
        ELSIF x = 1028 THEN
            tanh_f := 950;
        ELSIF x = 1029 THEN
            tanh_f := 951;
        ELSIF x = 1030 THEN
            tanh_f := 952;
        ELSIF x = 1031 THEN
            tanh_f := 953;
        ELSIF x = 1032 THEN
            tanh_f := 953;
        ELSIF x = 1033 THEN
            tanh_f := 954;
        ELSIF x = 1034 THEN
            tanh_f := 955;
        ELSIF x = 1035 THEN
            tanh_f := 956;
        ELSIF x = 1036 THEN
            tanh_f := 956;
        ELSIF x = 1037 THEN
            tanh_f := 957;
        ELSIF x = 1038 THEN
            tanh_f := 958;
        ELSIF x = 1039 THEN
            tanh_f := 959;
        ELSIF x = 1040 THEN
            tanh_f := 959;
        ELSIF x = 1041 THEN
            tanh_f := 960;
        ELSIF x = 1042 THEN
            tanh_f := 961;
        ELSIF x = 1043 THEN
            tanh_f := 962;
        ELSIF x = 1044 THEN
            tanh_f := 962;
        ELSIF x = 1045 THEN
            tanh_f := 963;
        ELSIF x = 1046 THEN
            tanh_f := 964;
        ELSIF x = 1047 THEN
            tanh_f := 965;
        ELSIF x = 1048 THEN
            tanh_f := 965;
        ELSIF x = 1049 THEN
            tanh_f := 966;
        ELSIF x = 1050 THEN
            tanh_f := 967;
        ELSIF x = 1051 THEN
            tanh_f := 968;
        ELSIF x = 1052 THEN
            tanh_f := 968;
        ELSIF x = 1053 THEN
            tanh_f := 969;
        ELSIF x = 1054 THEN
            tanh_f := 970;
        ELSIF x = 1055 THEN
            tanh_f := 971;
        ELSIF x = 1056 THEN
            tanh_f := 971;
        ELSIF x = 1057 THEN
            tanh_f := 972;
        ELSIF x = 1058 THEN
            tanh_f := 973;
        ELSIF x = 1059 THEN
            tanh_f := 974;
        ELSIF x = 1060 THEN
            tanh_f := 974;
        ELSIF x = 1061 THEN
            tanh_f := 975;
        ELSIF x = 1062 THEN
            tanh_f := 976;
        ELSIF x = 1063 THEN
            tanh_f := 977;
        ELSIF x = 1064 THEN
            tanh_f := 977;
        ELSIF x = 1065 THEN
            tanh_f := 978;
        ELSIF x = 1066 THEN
            tanh_f := 979;
        ELSIF x = 1067 THEN
            tanh_f := 979;
        ELSIF x = 1068 THEN
            tanh_f := 980;
        ELSIF x = 1069 THEN
            tanh_f := 981;
        ELSIF x = 1070 THEN
            tanh_f := 982;
        ELSIF x = 1071 THEN
            tanh_f := 982;
        ELSIF x = 1072 THEN
            tanh_f := 983;
        ELSIF x = 1073 THEN
            tanh_f := 984;
        ELSIF x = 1074 THEN
            tanh_f := 985;
        ELSIF x = 1075 THEN
            tanh_f := 985;
        ELSIF x = 1076 THEN
            tanh_f := 986;
        ELSIF x = 1077 THEN
            tanh_f := 987;
        ELSIF x = 1078 THEN
            tanh_f := 988;
        ELSIF x = 1079 THEN
            tanh_f := 988;
        ELSIF x = 1080 THEN
            tanh_f := 989;
        ELSIF x = 1081 THEN
            tanh_f := 990;
        ELSIF x = 1082 THEN
            tanh_f := 991;
        ELSIF x = 1083 THEN
            tanh_f := 991;
        ELSIF x = 1084 THEN
            tanh_f := 992;
        ELSIF x = 1085 THEN
            tanh_f := 993;
        ELSIF x = 1086 THEN
            tanh_f := 994;
        ELSIF x = 1087 THEN
            tanh_f := 994;
        ELSIF x = 1088 THEN
            tanh_f := 995;
        ELSIF x = 1089 THEN
            tanh_f := 996;
        ELSIF x = 1090 THEN
            tanh_f := 997;
        ELSIF x = 1091 THEN
            tanh_f := 997;
        ELSIF x = 1092 THEN
            tanh_f := 998;
        ELSIF x = 1093 THEN
            tanh_f := 999;
        ELSIF x = 1094 THEN
            tanh_f := 1000;
        ELSIF x = 1095 THEN
            tanh_f := 1000;
        ELSIF x = 1096 THEN
            tanh_f := 1001;
        ELSIF x = 1097 THEN
            tanh_f := 1002;
        ELSIF x = 1098 THEN
            tanh_f := 1003;
        ELSIF x = 1099 THEN
            tanh_f := 1003;
        ELSIF x = 1100 THEN
            tanh_f := 1004;
        ELSIF x = 1101 THEN
            tanh_f := 1005;
        ELSIF x = 1102 THEN
            tanh_f := 1006;
        ELSIF x = 1103 THEN
            tanh_f := 1006;
        ELSIF x = 1104 THEN
            tanh_f := 1007;
        ELSIF x = 1105 THEN
            tanh_f := 1008;
        ELSIF x = 1106 THEN
            tanh_f := 1009;
        ELSIF x = 1107 THEN
            tanh_f := 1009;
        ELSIF x = 1108 THEN
            tanh_f := 1010;
        ELSIF x = 1109 THEN
            tanh_f := 1011;
        ELSIF x = 1110 THEN
            tanh_f := 1011;
        ELSIF x = 1111 THEN
            tanh_f := 1012;
        ELSIF x = 1112 THEN
            tanh_f := 1013;
        ELSIF x = 1113 THEN
            tanh_f := 1014;
        ELSIF x = 1114 THEN
            tanh_f := 1014;
        ELSIF x = 1115 THEN
            tanh_f := 1015;
        ELSIF x = 1116 THEN
            tanh_f := 1016;
        ELSIF x = 1117 THEN
            tanh_f := 1017;
        ELSIF x = 1118 THEN
            tanh_f := 1017;
        ELSIF x = 1119 THEN
            tanh_f := 1018;
        ELSIF x = 1120 THEN
            tanh_f := 1019;
        ELSIF x = 1121 THEN
            tanh_f := 1020;
        ELSIF x = 1122 THEN
            tanh_f := 1020;
        ELSIF x = 1123 THEN
            tanh_f := 1021;
        ELSIF x = 1124 THEN
            tanh_f := 1022;
        ELSIF x = 1125 THEN
            tanh_f := 1023;
        ELSIF x = 1126 THEN
            tanh_f := 1023;
        ELSIF x = 1127 THEN
            tanh_f := 1024;
        ELSIF x = 1128 THEN
            tanh_f := 1025;
        ELSIF x = 1129 THEN
            tanh_f := 1026;
        ELSIF x = 1130 THEN
            tanh_f := 1026;
        ELSIF x = 1131 THEN
            tanh_f := 1027;
        ELSIF x = 1132 THEN
            tanh_f := 1028;
        ELSIF x = 1133 THEN
            tanh_f := 1029;
        ELSIF x = 1134 THEN
            tanh_f := 1029;
        ELSIF x = 1135 THEN
            tanh_f := 1030;
        ELSIF x = 1136 THEN
            tanh_f := 1031;
        ELSIF x = 1137 THEN
            tanh_f := 1032;
        ELSIF x = 1138 THEN
            tanh_f := 1032;
        ELSIF x = 1139 THEN
            tanh_f := 1033;
        ELSIF x = 1140 THEN
            tanh_f := 1034;
        ELSIF x = 1141 THEN
            tanh_f := 1035;
        ELSIF x = 1142 THEN
            tanh_f := 1035;
        ELSIF x = 1143 THEN
            tanh_f := 1036;
        ELSIF x = 1144 THEN
            tanh_f := 1037;
        ELSIF x = 1145 THEN
            tanh_f := 1038;
        ELSIF x = 1146 THEN
            tanh_f := 1038;
        ELSIF x = 1147 THEN
            tanh_f := 1039;
        ELSIF x = 1148 THEN
            tanh_f := 1040;
        ELSIF x = 1149 THEN
            tanh_f := 1041;
        ELSIF x = 1150 THEN
            tanh_f := 1041;
        ELSIF x = 1151 THEN
            tanh_f := 1042;
        ELSIF x = 1152 THEN
            tanh_f := 1043;
        ELSIF x = 1153 THEN
            tanh_f := 1043;
        ELSIF x = 1154 THEN
            tanh_f := 1044;
        ELSIF x = 1155 THEN
            tanh_f := 1045;
        ELSIF x = 1156 THEN
            tanh_f := 1046;
        ELSIF x = 1157 THEN
            tanh_f := 1046;
        ELSIF x = 1158 THEN
            tanh_f := 1047;
        ELSIF x = 1159 THEN
            tanh_f := 1048;
        ELSIF x = 1160 THEN
            tanh_f := 1049;
        ELSIF x = 1161 THEN
            tanh_f := 1049;
        ELSIF x = 1162 THEN
            tanh_f := 1050;
        ELSIF x = 1163 THEN
            tanh_f := 1051;
        ELSIF x = 1164 THEN
            tanh_f := 1052;
        ELSIF x = 1165 THEN
            tanh_f := 1052;
        ELSIF x = 1166 THEN
            tanh_f := 1053;
        ELSIF x = 1167 THEN
            tanh_f := 1054;
        ELSIF x = 1168 THEN
            tanh_f := 1055;
        ELSIF x = 1169 THEN
            tanh_f := 1055;
        ELSIF x = 1170 THEN
            tanh_f := 1056;
        ELSIF x = 1171 THEN
            tanh_f := 1057;
        ELSIF x = 1172 THEN
            tanh_f := 1058;
        ELSIF x = 1173 THEN
            tanh_f := 1058;
        ELSIF x = 1174 THEN
            tanh_f := 1059;
        ELSIF x = 1175 THEN
            tanh_f := 1060;
        ELSIF x = 1176 THEN
            tanh_f := 1061;
        ELSIF x = 1177 THEN
            tanh_f := 1061;
        ELSIF x = 1178 THEN
            tanh_f := 1062;
        ELSIF x = 1179 THEN
            tanh_f := 1063;
        ELSIF x = 1180 THEN
            tanh_f := 1064;
        ELSIF x = 1181 THEN
            tanh_f := 1064;
        ELSIF x = 1182 THEN
            tanh_f := 1065;
        ELSIF x = 1183 THEN
            tanh_f := 1066;
        ELSIF x = 1184 THEN
            tanh_f := 1067;
        ELSIF x = 1185 THEN
            tanh_f := 1067;
        ELSIF x = 1186 THEN
            tanh_f := 1068;
        ELSIF x = 1187 THEN
            tanh_f := 1069;
        ELSIF x = 1188 THEN
            tanh_f := 1070;
        ELSIF x = 1189 THEN
            tanh_f := 1070;
        ELSIF x = 1190 THEN
            tanh_f := 1071;
        ELSIF x = 1191 THEN
            tanh_f := 1072;
        ELSIF x = 1192 THEN
            tanh_f := 1073;
        ELSIF x = 1193 THEN
            tanh_f := 1073;
        ELSIF x = 1194 THEN
            tanh_f := 1074;
        ELSIF x = 1195 THEN
            tanh_f := 1075;
        ELSIF x = 1196 THEN
            tanh_f := 1075;
        ELSIF x = 1197 THEN
            tanh_f := 1076;
        ELSIF x = 1198 THEN
            tanh_f := 1077;
        ELSIF x = 1199 THEN
            tanh_f := 1078;
        ELSIF x = 1200 THEN
            tanh_f := 1078;
        ELSIF x = 1201 THEN
            tanh_f := 1079;
        ELSIF x = 1202 THEN
            tanh_f := 1080;
        ELSIF x = 1203 THEN
            tanh_f := 1081;
        ELSIF x = 1204 THEN
            tanh_f := 1081;
        ELSIF x = 1205 THEN
            tanh_f := 1082;
        ELSIF x = 1206 THEN
            tanh_f := 1083;
        ELSIF x = 1207 THEN
            tanh_f := 1084;
        ELSIF x = 1208 THEN
            tanh_f := 1084;
        ELSIF x = 1209 THEN
            tanh_f := 1085;
        ELSIF x = 1210 THEN
            tanh_f := 1086;
        ELSIF x = 1211 THEN
            tanh_f := 1087;
        ELSIF x = 1212 THEN
            tanh_f := 1087;
        ELSIF x = 1213 THEN
            tanh_f := 1088;
        ELSIF x = 1214 THEN
            tanh_f := 1089;
        ELSIF x = 1215 THEN
            tanh_f := 1090;
        ELSIF x = 1216 THEN
            tanh_f := 1090;
        ELSIF x = 1217 THEN
            tanh_f := 1091;
        ELSIF x = 1218 THEN
            tanh_f := 1092;
        ELSIF x = 1219 THEN
            tanh_f := 1093;
        ELSIF x = 1220 THEN
            tanh_f := 1093;
        ELSIF x = 1221 THEN
            tanh_f := 1094;
        ELSIF x = 1222 THEN
            tanh_f := 1095;
        ELSIF x = 1223 THEN
            tanh_f := 1096;
        ELSIF x = 1224 THEN
            tanh_f := 1096;
        ELSIF x = 1225 THEN
            tanh_f := 1097;
        ELSIF x = 1226 THEN
            tanh_f := 1098;
        ELSIF x = 1227 THEN
            tanh_f := 1099;
        ELSIF x = 1228 THEN
            tanh_f := 1099;
        ELSIF x = 1229 THEN
            tanh_f := 1100;
        ELSIF x = 1230 THEN
            tanh_f := 1101;
        ELSIF x = 1231 THEN
            tanh_f := 1102;
        ELSIF x = 1232 THEN
            tanh_f := 1102;
        ELSIF x = 1233 THEN
            tanh_f := 1103;
        ELSIF x = 1234 THEN
            tanh_f := 1104;
        ELSIF x = 1235 THEN
            tanh_f := 1105;
        ELSIF x = 1236 THEN
            tanh_f := 1105;
        ELSIF x = 1237 THEN
            tanh_f := 1106;
        ELSIF x = 1238 THEN
            tanh_f := 1107;
        ELSIF x = 1239 THEN
            tanh_f := 1107;
        ELSIF x = 1240 THEN
            tanh_f := 1108;
        ELSIF x = 1241 THEN
            tanh_f := 1109;
        ELSIF x = 1242 THEN
            tanh_f := 1110;
        ELSIF x = 1243 THEN
            tanh_f := 1110;
        ELSIF x = 1244 THEN
            tanh_f := 1111;
        ELSIF x = 1245 THEN
            tanh_f := 1112;
        ELSIF x = 1246 THEN
            tanh_f := 1113;
        ELSIF x = 1247 THEN
            tanh_f := 1113;
        ELSIF x = 1248 THEN
            tanh_f := 1114;
        ELSIF x = 1249 THEN
            tanh_f := 1115;
        ELSIF x = 1250 THEN
            tanh_f := 1116;
        ELSIF x = 1251 THEN
            tanh_f := 1116;
        ELSIF x = 1252 THEN
            tanh_f := 1117;
        ELSIF x = 1253 THEN
            tanh_f := 1118;
        ELSIF x = 1254 THEN
            tanh_f := 1119;
        ELSIF x = 1255 THEN
            tanh_f := 1119;
        ELSIF x = 1256 THEN
            tanh_f := 1120;
        ELSIF x = 1257 THEN
            tanh_f := 1121;
        ELSIF x = 1258 THEN
            tanh_f := 1122;
        ELSIF x = 1259 THEN
            tanh_f := 1122;
        ELSIF x = 1260 THEN
            tanh_f := 1123;
        ELSIF x = 1261 THEN
            tanh_f := 1124;
        ELSIF x = 1262 THEN
            tanh_f := 1125;
        ELSIF x = 1263 THEN
            tanh_f := 1125;
        ELSIF x = 1264 THEN
            tanh_f := 1126;
        ELSIF x = 1265 THEN
            tanh_f := 1127;
        ELSIF x = 1266 THEN
            tanh_f := 1128;
        ELSIF x = 1267 THEN
            tanh_f := 1128;
        ELSIF x = 1268 THEN
            tanh_f := 1129;
        ELSIF x = 1269 THEN
            tanh_f := 1130;
        ELSIF x = 1270 THEN
            tanh_f := 1131;
        ELSIF x = 1271 THEN
            tanh_f := 1131;
        ELSIF x = 1272 THEN
            tanh_f := 1132;
        ELSIF x = 1273 THEN
            tanh_f := 1133;
        ELSIF x = 1274 THEN
            tanh_f := 1134;
        ELSIF x = 1275 THEN
            tanh_f := 1134;
        ELSIF x = 1276 THEN
            tanh_f := 1135;
        ELSIF x = 1277 THEN
            tanh_f := 1136;
        ELSIF x = 1278 THEN
            tanh_f := 1137;
        ELSIF x = 1279 THEN
            tanh_f := 1137;
        ELSIF x = 1280 THEN
            tanh_f := 1138;
        ELSIF x = 1281 THEN
            tanh_f := 1139;
        ELSIF x = 1282 THEN
            tanh_f := 1139;
        ELSIF x = 1283 THEN
            tanh_f := 1140;
        ELSIF x = 1284 THEN
            tanh_f := 1141;
        ELSIF x = 1285 THEN
            tanh_f := 1141;
        ELSIF x = 1286 THEN
            tanh_f := 1142;
        ELSIF x = 1287 THEN
            tanh_f := 1142;
        ELSIF x = 1288 THEN
            tanh_f := 1143;
        ELSIF x = 1289 THEN
            tanh_f := 1144;
        ELSIF x = 1290 THEN
            tanh_f := 1144;
        ELSIF x = 1291 THEN
            tanh_f := 1145;
        ELSIF x = 1292 THEN
            tanh_f := 1146;
        ELSIF x = 1293 THEN
            tanh_f := 1146;
        ELSIF x = 1294 THEN
            tanh_f := 1147;
        ELSIF x = 1295 THEN
            tanh_f := 1148;
        ELSIF x = 1296 THEN
            tanh_f := 1148;
        ELSIF x = 1297 THEN
            tanh_f := 1149;
        ELSIF x = 1298 THEN
            tanh_f := 1150;
        ELSIF x = 1299 THEN
            tanh_f := 1150;
        ELSIF x = 1300 THEN
            tanh_f := 1151;
        ELSIF x = 1301 THEN
            tanh_f := 1151;
        ELSIF x = 1302 THEN
            tanh_f := 1152;
        ELSIF x = 1303 THEN
            tanh_f := 1153;
        ELSIF x = 1304 THEN
            tanh_f := 1153;
        ELSIF x = 1305 THEN
            tanh_f := 1154;
        ELSIF x = 1306 THEN
            tanh_f := 1155;
        ELSIF x = 1307 THEN
            tanh_f := 1155;
        ELSIF x = 1308 THEN
            tanh_f := 1156;
        ELSIF x = 1309 THEN
            tanh_f := 1157;
        ELSIF x = 1310 THEN
            tanh_f := 1157;
        ELSIF x = 1311 THEN
            tanh_f := 1158;
        ELSIF x = 1312 THEN
            tanh_f := 1159;
        ELSIF x = 1313 THEN
            tanh_f := 1159;
        ELSIF x = 1314 THEN
            tanh_f := 1160;
        ELSIF x = 1315 THEN
            tanh_f := 1160;
        ELSIF x = 1316 THEN
            tanh_f := 1161;
        ELSIF x = 1317 THEN
            tanh_f := 1162;
        ELSIF x = 1318 THEN
            tanh_f := 1162;
        ELSIF x = 1319 THEN
            tanh_f := 1163;
        ELSIF x = 1320 THEN
            tanh_f := 1164;
        ELSIF x = 1321 THEN
            tanh_f := 1164;
        ELSIF x = 1322 THEN
            tanh_f := 1165;
        ELSIF x = 1323 THEN
            tanh_f := 1166;
        ELSIF x = 1324 THEN
            tanh_f := 1166;
        ELSIF x = 1325 THEN
            tanh_f := 1167;
        ELSIF x = 1326 THEN
            tanh_f := 1168;
        ELSIF x = 1327 THEN
            tanh_f := 1168;
        ELSIF x = 1328 THEN
            tanh_f := 1169;
        ELSIF x = 1329 THEN
            tanh_f := 1169;
        ELSIF x = 1330 THEN
            tanh_f := 1170;
        ELSIF x = 1331 THEN
            tanh_f := 1171;
        ELSIF x = 1332 THEN
            tanh_f := 1171;
        ELSIF x = 1333 THEN
            tanh_f := 1172;
        ELSIF x = 1334 THEN
            tanh_f := 1173;
        ELSIF x = 1335 THEN
            tanh_f := 1173;
        ELSIF x = 1336 THEN
            tanh_f := 1174;
        ELSIF x = 1337 THEN
            tanh_f := 1175;
        ELSIF x = 1338 THEN
            tanh_f := 1175;
        ELSIF x = 1339 THEN
            tanh_f := 1176;
        ELSIF x = 1340 THEN
            tanh_f := 1177;
        ELSIF x = 1341 THEN
            tanh_f := 1177;
        ELSIF x = 1342 THEN
            tanh_f := 1178;
        ELSIF x = 1343 THEN
            tanh_f := 1178;
        ELSIF x = 1344 THEN
            tanh_f := 1179;
        ELSIF x = 1345 THEN
            tanh_f := 1180;
        ELSIF x = 1346 THEN
            tanh_f := 1180;
        ELSIF x = 1347 THEN
            tanh_f := 1181;
        ELSIF x = 1348 THEN
            tanh_f := 1182;
        ELSIF x = 1349 THEN
            tanh_f := 1182;
        ELSIF x = 1350 THEN
            tanh_f := 1183;
        ELSIF x = 1351 THEN
            tanh_f := 1184;
        ELSIF x = 1352 THEN
            tanh_f := 1184;
        ELSIF x = 1353 THEN
            tanh_f := 1185;
        ELSIF x = 1354 THEN
            tanh_f := 1186;
        ELSIF x = 1355 THEN
            tanh_f := 1186;
        ELSIF x = 1356 THEN
            tanh_f := 1187;
        ELSIF x = 1357 THEN
            tanh_f := 1187;
        ELSIF x = 1358 THEN
            tanh_f := 1188;
        ELSIF x = 1359 THEN
            tanh_f := 1189;
        ELSIF x = 1360 THEN
            tanh_f := 1189;
        ELSIF x = 1361 THEN
            tanh_f := 1190;
        ELSIF x = 1362 THEN
            tanh_f := 1191;
        ELSIF x = 1363 THEN
            tanh_f := 1191;
        ELSIF x = 1364 THEN
            tanh_f := 1192;
        ELSIF x = 1365 THEN
            tanh_f := 1193;
        ELSIF x = 1366 THEN
            tanh_f := 1193;
        ELSIF x = 1367 THEN
            tanh_f := 1194;
        ELSIF x = 1368 THEN
            tanh_f := 1195;
        ELSIF x = 1369 THEN
            tanh_f := 1195;
        ELSIF x = 1370 THEN
            tanh_f := 1196;
        ELSIF x = 1371 THEN
            tanh_f := 1196;
        ELSIF x = 1372 THEN
            tanh_f := 1197;
        ELSIF x = 1373 THEN
            tanh_f := 1198;
        ELSIF x = 1374 THEN
            tanh_f := 1198;
        ELSIF x = 1375 THEN
            tanh_f := 1199;
        ELSIF x = 1376 THEN
            tanh_f := 1200;
        ELSIF x = 1377 THEN
            tanh_f := 1200;
        ELSIF x = 1378 THEN
            tanh_f := 1201;
        ELSIF x = 1379 THEN
            tanh_f := 1202;
        ELSIF x = 1380 THEN
            tanh_f := 1202;
        ELSIF x = 1381 THEN
            tanh_f := 1203;
        ELSIF x = 1382 THEN
            tanh_f := 1204;
        ELSIF x = 1383 THEN
            tanh_f := 1204;
        ELSIF x = 1384 THEN
            tanh_f := 1205;
        ELSIF x = 1385 THEN
            tanh_f := 1205;
        ELSIF x = 1386 THEN
            tanh_f := 1206;
        ELSIF x = 1387 THEN
            tanh_f := 1207;
        ELSIF x = 1388 THEN
            tanh_f := 1207;
        ELSIF x = 1389 THEN
            tanh_f := 1208;
        ELSIF x = 1390 THEN
            tanh_f := 1209;
        ELSIF x = 1391 THEN
            tanh_f := 1209;
        ELSIF x = 1392 THEN
            tanh_f := 1210;
        ELSIF x = 1393 THEN
            tanh_f := 1211;
        ELSIF x = 1394 THEN
            tanh_f := 1211;
        ELSIF x = 1395 THEN
            tanh_f := 1212;
        ELSIF x = 1396 THEN
            tanh_f := 1213;
        ELSIF x = 1397 THEN
            tanh_f := 1213;
        ELSIF x = 1398 THEN
            tanh_f := 1214;
        ELSIF x = 1399 THEN
            tanh_f := 1214;
        ELSIF x = 1400 THEN
            tanh_f := 1215;
        ELSIF x = 1401 THEN
            tanh_f := 1216;
        ELSIF x = 1402 THEN
            tanh_f := 1216;
        ELSIF x = 1403 THEN
            tanh_f := 1217;
        ELSIF x = 1404 THEN
            tanh_f := 1218;
        ELSIF x = 1405 THEN
            tanh_f := 1218;
        ELSIF x = 1406 THEN
            tanh_f := 1219;
        ELSIF x = 1407 THEN
            tanh_f := 1220;
        ELSIF x = 1408 THEN
            tanh_f := 1220;
        ELSIF x = 1409 THEN
            tanh_f := 1221;
        ELSIF x = 1410 THEN
            tanh_f := 1222;
        ELSIF x = 1411 THEN
            tanh_f := 1222;
        ELSIF x = 1412 THEN
            tanh_f := 1223;
        ELSIF x = 1413 THEN
            tanh_f := 1223;
        ELSIF x = 1414 THEN
            tanh_f := 1224;
        ELSIF x = 1415 THEN
            tanh_f := 1225;
        ELSIF x = 1416 THEN
            tanh_f := 1225;
        ELSIF x = 1417 THEN
            tanh_f := 1226;
        ELSIF x = 1418 THEN
            tanh_f := 1227;
        ELSIF x = 1419 THEN
            tanh_f := 1227;
        ELSIF x = 1420 THEN
            tanh_f := 1228;
        ELSIF x = 1421 THEN
            tanh_f := 1229;
        ELSIF x = 1422 THEN
            tanh_f := 1229;
        ELSIF x = 1423 THEN
            tanh_f := 1230;
        ELSIF x = 1424 THEN
            tanh_f := 1231;
        ELSIF x = 1425 THEN
            tanh_f := 1231;
        ELSIF x = 1426 THEN
            tanh_f := 1232;
        ELSIF x = 1427 THEN
            tanh_f := 1232;
        ELSIF x = 1428 THEN
            tanh_f := 1233;
        ELSIF x = 1429 THEN
            tanh_f := 1234;
        ELSIF x = 1430 THEN
            tanh_f := 1234;
        ELSIF x = 1431 THEN
            tanh_f := 1235;
        ELSIF x = 1432 THEN
            tanh_f := 1236;
        ELSIF x = 1433 THEN
            tanh_f := 1236;
        ELSIF x = 1434 THEN
            tanh_f := 1237;
        ELSIF x = 1435 THEN
            tanh_f := 1238;
        ELSIF x = 1436 THEN
            tanh_f := 1238;
        ELSIF x = 1437 THEN
            tanh_f := 1239;
        ELSIF x = 1438 THEN
            tanh_f := 1240;
        ELSIF x = 1439 THEN
            tanh_f := 1240;
        ELSIF x = 1440 THEN
            tanh_f := 1241;
        ELSIF x = 1441 THEN
            tanh_f := 1241;
        ELSIF x = 1442 THEN
            tanh_f := 1242;
        ELSIF x = 1443 THEN
            tanh_f := 1243;
        ELSIF x = 1444 THEN
            tanh_f := 1243;
        ELSIF x = 1445 THEN
            tanh_f := 1244;
        ELSIF x = 1446 THEN
            tanh_f := 1245;
        ELSIF x = 1447 THEN
            tanh_f := 1245;
        ELSIF x = 1448 THEN
            tanh_f := 1246;
        ELSIF x = 1449 THEN
            tanh_f := 1247;
        ELSIF x = 1450 THEN
            tanh_f := 1247;
        ELSIF x = 1451 THEN
            tanh_f := 1248;
        ELSIF x = 1452 THEN
            tanh_f := 1249;
        ELSIF x = 1453 THEN
            tanh_f := 1249;
        ELSIF x = 1454 THEN
            tanh_f := 1250;
        ELSIF x = 1455 THEN
            tanh_f := 1250;
        ELSIF x = 1456 THEN
            tanh_f := 1251;
        ELSIF x = 1457 THEN
            tanh_f := 1252;
        ELSIF x = 1458 THEN
            tanh_f := 1252;
        ELSIF x = 1459 THEN
            tanh_f := 1253;
        ELSIF x = 1460 THEN
            tanh_f := 1254;
        ELSIF x = 1461 THEN
            tanh_f := 1254;
        ELSIF x = 1462 THEN
            tanh_f := 1255;
        ELSIF x = 1463 THEN
            tanh_f := 1256;
        ELSIF x = 1464 THEN
            tanh_f := 1256;
        ELSIF x = 1465 THEN
            tanh_f := 1257;
        ELSIF x = 1466 THEN
            tanh_f := 1258;
        ELSIF x = 1467 THEN
            tanh_f := 1258;
        ELSIF x = 1468 THEN
            tanh_f := 1259;
        ELSIF x = 1469 THEN
            tanh_f := 1259;
        ELSIF x = 1470 THEN
            tanh_f := 1260;
        ELSIF x = 1471 THEN
            tanh_f := 1261;
        ELSIF x = 1472 THEN
            tanh_f := 1261;
        ELSIF x = 1473 THEN
            tanh_f := 1262;
        ELSIF x = 1474 THEN
            tanh_f := 1263;
        ELSIF x = 1475 THEN
            tanh_f := 1263;
        ELSIF x = 1476 THEN
            tanh_f := 1264;
        ELSIF x = 1477 THEN
            tanh_f := 1265;
        ELSIF x = 1478 THEN
            tanh_f := 1265;
        ELSIF x = 1479 THEN
            tanh_f := 1266;
        ELSIF x = 1480 THEN
            tanh_f := 1267;
        ELSIF x = 1481 THEN
            tanh_f := 1267;
        ELSIF x = 1482 THEN
            tanh_f := 1268;
        ELSIF x = 1483 THEN
            tanh_f := 1268;
        ELSIF x = 1484 THEN
            tanh_f := 1269;
        ELSIF x = 1485 THEN
            tanh_f := 1270;
        ELSIF x = 1486 THEN
            tanh_f := 1270;
        ELSIF x = 1487 THEN
            tanh_f := 1271;
        ELSIF x = 1488 THEN
            tanh_f := 1272;
        ELSIF x = 1489 THEN
            tanh_f := 1272;
        ELSIF x = 1490 THEN
            tanh_f := 1273;
        ELSIF x = 1491 THEN
            tanh_f := 1274;
        ELSIF x = 1492 THEN
            tanh_f := 1274;
        ELSIF x = 1493 THEN
            tanh_f := 1275;
        ELSIF x = 1494 THEN
            tanh_f := 1276;
        ELSIF x = 1495 THEN
            tanh_f := 1276;
        ELSIF x = 1496 THEN
            tanh_f := 1277;
        ELSIF x = 1497 THEN
            tanh_f := 1277;
        ELSIF x = 1498 THEN
            tanh_f := 1278;
        ELSIF x = 1499 THEN
            tanh_f := 1279;
        ELSIF x = 1500 THEN
            tanh_f := 1279;
        ELSIF x = 1501 THEN
            tanh_f := 1280;
        ELSIF x = 1502 THEN
            tanh_f := 1281;
        ELSIF x = 1503 THEN
            tanh_f := 1281;
        ELSIF x = 1504 THEN
            tanh_f := 1282;
        ELSIF x = 1505 THEN
            tanh_f := 1283;
        ELSIF x = 1506 THEN
            tanh_f := 1283;
        ELSIF x = 1507 THEN
            tanh_f := 1284;
        ELSIF x = 1508 THEN
            tanh_f := 1285;
        ELSIF x = 1509 THEN
            tanh_f := 1285;
        ELSIF x = 1510 THEN
            tanh_f := 1286;
        ELSIF x = 1511 THEN
            tanh_f := 1286;
        ELSIF x = 1512 THEN
            tanh_f := 1287;
        ELSIF x = 1513 THEN
            tanh_f := 1288;
        ELSIF x = 1514 THEN
            tanh_f := 1288;
        ELSIF x = 1515 THEN
            tanh_f := 1289;
        ELSIF x = 1516 THEN
            tanh_f := 1290;
        ELSIF x = 1517 THEN
            tanh_f := 1290;
        ELSIF x = 1518 THEN
            tanh_f := 1291;
        ELSIF x = 1519 THEN
            tanh_f := 1292;
        ELSIF x = 1520 THEN
            tanh_f := 1292;
        ELSIF x = 1521 THEN
            tanh_f := 1293;
        ELSIF x = 1522 THEN
            tanh_f := 1294;
        ELSIF x = 1523 THEN
            tanh_f := 1294;
        ELSIF x = 1524 THEN
            tanh_f := 1295;
        ELSIF x = 1525 THEN
            tanh_f := 1295;
        ELSIF x = 1526 THEN
            tanh_f := 1296;
        ELSIF x = 1527 THEN
            tanh_f := 1297;
        ELSIF x = 1528 THEN
            tanh_f := 1297;
        ELSIF x = 1529 THEN
            tanh_f := 1298;
        ELSIF x = 1530 THEN
            tanh_f := 1299;
        ELSIF x = 1531 THEN
            tanh_f := 1299;
        ELSIF x = 1532 THEN
            tanh_f := 1300;
        ELSIF x = 1533 THEN
            tanh_f := 1301;
        ELSIF x = 1534 THEN
            tanh_f := 1301;
        ELSIF x = 1535 THEN
            tanh_f := 1302;
        ELSIF x = 1536 THEN
            tanh_f := 1303;
        ELSIF x = 1537 THEN
            tanh_f := 1303;
        ELSIF x = 1538 THEN
            tanh_f := 1304;
        ELSIF x = 1539 THEN
            tanh_f := 1304;
        ELSIF x = 1540 THEN
            tanh_f := 1305;
        ELSIF x = 1541 THEN
            tanh_f := 1305;
        ELSIF x = 1542 THEN
            tanh_f := 1306;
        ELSIF x = 1543 THEN
            tanh_f := 1306;
        ELSIF x = 1544 THEN
            tanh_f := 1307;
        ELSIF x = 1545 THEN
            tanh_f := 1307;
        ELSIF x = 1546 THEN
            tanh_f := 1308;
        ELSIF x = 1547 THEN
            tanh_f := 1309;
        ELSIF x = 1548 THEN
            tanh_f := 1309;
        ELSIF x = 1549 THEN
            tanh_f := 1310;
        ELSIF x = 1550 THEN
            tanh_f := 1310;
        ELSIF x = 1551 THEN
            tanh_f := 1311;
        ELSIF x = 1552 THEN
            tanh_f := 1311;
        ELSIF x = 1553 THEN
            tanh_f := 1312;
        ELSIF x = 1554 THEN
            tanh_f := 1312;
        ELSIF x = 1555 THEN
            tanh_f := 1313;
        ELSIF x = 1556 THEN
            tanh_f := 1313;
        ELSIF x = 1557 THEN
            tanh_f := 1314;
        ELSIF x = 1558 THEN
            tanh_f := 1315;
        ELSIF x = 1559 THEN
            tanh_f := 1315;
        ELSIF x = 1560 THEN
            tanh_f := 1316;
        ELSIF x = 1561 THEN
            tanh_f := 1316;
        ELSIF x = 1562 THEN
            tanh_f := 1317;
        ELSIF x = 1563 THEN
            tanh_f := 1317;
        ELSIF x = 1564 THEN
            tanh_f := 1318;
        ELSIF x = 1565 THEN
            tanh_f := 1318;
        ELSIF x = 1566 THEN
            tanh_f := 1319;
        ELSIF x = 1567 THEN
            tanh_f := 1320;
        ELSIF x = 1568 THEN
            tanh_f := 1320;
        ELSIF x = 1569 THEN
            tanh_f := 1321;
        ELSIF x = 1570 THEN
            tanh_f := 1321;
        ELSIF x = 1571 THEN
            tanh_f := 1322;
        ELSIF x = 1572 THEN
            tanh_f := 1322;
        ELSIF x = 1573 THEN
            tanh_f := 1323;
        ELSIF x = 1574 THEN
            tanh_f := 1323;
        ELSIF x = 1575 THEN
            tanh_f := 1324;
        ELSIF x = 1576 THEN
            tanh_f := 1324;
        ELSIF x = 1577 THEN
            tanh_f := 1325;
        ELSIF x = 1578 THEN
            tanh_f := 1326;
        ELSIF x = 1579 THEN
            tanh_f := 1326;
        ELSIF x = 1580 THEN
            tanh_f := 1327;
        ELSIF x = 1581 THEN
            tanh_f := 1327;
        ELSIF x = 1582 THEN
            tanh_f := 1328;
        ELSIF x = 1583 THEN
            tanh_f := 1328;
        ELSIF x = 1584 THEN
            tanh_f := 1329;
        ELSIF x = 1585 THEN
            tanh_f := 1329;
        ELSIF x = 1586 THEN
            tanh_f := 1330;
        ELSIF x = 1587 THEN
            tanh_f := 1330;
        ELSIF x = 1588 THEN
            tanh_f := 1331;
        ELSIF x = 1589 THEN
            tanh_f := 1332;
        ELSIF x = 1590 THEN
            tanh_f := 1332;
        ELSIF x = 1591 THEN
            tanh_f := 1333;
        ELSIF x = 1592 THEN
            tanh_f := 1333;
        ELSIF x = 1593 THEN
            tanh_f := 1334;
        ELSIF x = 1594 THEN
            tanh_f := 1334;
        ELSIF x = 1595 THEN
            tanh_f := 1335;
        ELSIF x = 1596 THEN
            tanh_f := 1335;
        ELSIF x = 1597 THEN
            tanh_f := 1336;
        ELSIF x = 1598 THEN
            tanh_f := 1337;
        ELSIF x = 1599 THEN
            tanh_f := 1337;
        ELSIF x = 1600 THEN
            tanh_f := 1338;
        ELSIF x = 1601 THEN
            tanh_f := 1338;
        ELSIF x = 1602 THEN
            tanh_f := 1339;
        ELSIF x = 1603 THEN
            tanh_f := 1339;
        ELSIF x = 1604 THEN
            tanh_f := 1340;
        ELSIF x = 1605 THEN
            tanh_f := 1340;
        ELSIF x = 1606 THEN
            tanh_f := 1341;
        ELSIF x = 1607 THEN
            tanh_f := 1341;
        ELSIF x = 1608 THEN
            tanh_f := 1342;
        ELSIF x = 1609 THEN
            tanh_f := 1343;
        ELSIF x = 1610 THEN
            tanh_f := 1343;
        ELSIF x = 1611 THEN
            tanh_f := 1344;
        ELSIF x = 1612 THEN
            tanh_f := 1344;
        ELSIF x = 1613 THEN
            tanh_f := 1345;
        ELSIF x = 1614 THEN
            tanh_f := 1345;
        ELSIF x = 1615 THEN
            tanh_f := 1346;
        ELSIF x = 1616 THEN
            tanh_f := 1346;
        ELSIF x = 1617 THEN
            tanh_f := 1347;
        ELSIF x = 1618 THEN
            tanh_f := 1348;
        ELSIF x = 1619 THEN
            tanh_f := 1348;
        ELSIF x = 1620 THEN
            tanh_f := 1349;
        ELSIF x = 1621 THEN
            tanh_f := 1349;
        ELSIF x = 1622 THEN
            tanh_f := 1350;
        ELSIF x = 1623 THEN
            tanh_f := 1350;
        ELSIF x = 1624 THEN
            tanh_f := 1351;
        ELSIF x = 1625 THEN
            tanh_f := 1351;
        ELSIF x = 1626 THEN
            tanh_f := 1352;
        ELSIF x = 1627 THEN
            tanh_f := 1352;
        ELSIF x = 1628 THEN
            tanh_f := 1353;
        ELSIF x = 1629 THEN
            tanh_f := 1354;
        ELSIF x = 1630 THEN
            tanh_f := 1354;
        ELSIF x = 1631 THEN
            tanh_f := 1355;
        ELSIF x = 1632 THEN
            tanh_f := 1355;
        ELSIF x = 1633 THEN
            tanh_f := 1356;
        ELSIF x = 1634 THEN
            tanh_f := 1356;
        ELSIF x = 1635 THEN
            tanh_f := 1357;
        ELSIF x = 1636 THEN
            tanh_f := 1357;
        ELSIF x = 1637 THEN
            tanh_f := 1358;
        ELSIF x = 1638 THEN
            tanh_f := 1358;
        ELSIF x = 1639 THEN
            tanh_f := 1359;
        ELSIF x = 1640 THEN
            tanh_f := 1360;
        ELSIF x = 1641 THEN
            tanh_f := 1360;
        ELSIF x = 1642 THEN
            tanh_f := 1361;
        ELSIF x = 1643 THEN
            tanh_f := 1361;
        ELSIF x = 1644 THEN
            tanh_f := 1362;
        ELSIF x = 1645 THEN
            tanh_f := 1362;
        ELSIF x = 1646 THEN
            tanh_f := 1363;
        ELSIF x = 1647 THEN
            tanh_f := 1363;
        ELSIF x = 1648 THEN
            tanh_f := 1364;
        ELSIF x = 1649 THEN
            tanh_f := 1365;
        ELSIF x = 1650 THEN
            tanh_f := 1365;
        ELSIF x = 1651 THEN
            tanh_f := 1366;
        ELSIF x = 1652 THEN
            tanh_f := 1366;
        ELSIF x = 1653 THEN
            tanh_f := 1367;
        ELSIF x = 1654 THEN
            tanh_f := 1367;
        ELSIF x = 1655 THEN
            tanh_f := 1368;
        ELSIF x = 1656 THEN
            tanh_f := 1368;
        ELSIF x = 1657 THEN
            tanh_f := 1369;
        ELSIF x = 1658 THEN
            tanh_f := 1369;
        ELSIF x = 1659 THEN
            tanh_f := 1370;
        ELSIF x = 1660 THEN
            tanh_f := 1371;
        ELSIF x = 1661 THEN
            tanh_f := 1371;
        ELSIF x = 1662 THEN
            tanh_f := 1372;
        ELSIF x = 1663 THEN
            tanh_f := 1372;
        ELSIF x = 1664 THEN
            tanh_f := 1373;
        ELSIF x = 1665 THEN
            tanh_f := 1373;
        ELSIF x = 1666 THEN
            tanh_f := 1374;
        ELSIF x = 1667 THEN
            tanh_f := 1374;
        ELSIF x = 1668 THEN
            tanh_f := 1375;
        ELSIF x = 1669 THEN
            tanh_f := 1375;
        ELSIF x = 1670 THEN
            tanh_f := 1376;
        ELSIF x = 1671 THEN
            tanh_f := 1377;
        ELSIF x = 1672 THEN
            tanh_f := 1377;
        ELSIF x = 1673 THEN
            tanh_f := 1378;
        ELSIF x = 1674 THEN
            tanh_f := 1378;
        ELSIF x = 1675 THEN
            tanh_f := 1379;
        ELSIF x = 1676 THEN
            tanh_f := 1379;
        ELSIF x = 1677 THEN
            tanh_f := 1380;
        ELSIF x = 1678 THEN
            tanh_f := 1380;
        ELSIF x = 1679 THEN
            tanh_f := 1381;
        ELSIF x = 1680 THEN
            tanh_f := 1382;
        ELSIF x = 1681 THEN
            tanh_f := 1382;
        ELSIF x = 1682 THEN
            tanh_f := 1383;
        ELSIF x = 1683 THEN
            tanh_f := 1383;
        ELSIF x = 1684 THEN
            tanh_f := 1384;
        ELSIF x = 1685 THEN
            tanh_f := 1384;
        ELSIF x = 1686 THEN
            tanh_f := 1385;
        ELSIF x = 1687 THEN
            tanh_f := 1385;
        ELSIF x = 1688 THEN
            tanh_f := 1386;
        ELSIF x = 1689 THEN
            tanh_f := 1386;
        ELSIF x = 1690 THEN
            tanh_f := 1387;
        ELSIF x = 1691 THEN
            tanh_f := 1388;
        ELSIF x = 1692 THEN
            tanh_f := 1388;
        ELSIF x = 1693 THEN
            tanh_f := 1389;
        ELSIF x = 1694 THEN
            tanh_f := 1389;
        ELSIF x = 1695 THEN
            tanh_f := 1390;
        ELSIF x = 1696 THEN
            tanh_f := 1390;
        ELSIF x = 1697 THEN
            tanh_f := 1391;
        ELSIF x = 1698 THEN
            tanh_f := 1391;
        ELSIF x = 1699 THEN
            tanh_f := 1392;
        ELSIF x = 1700 THEN
            tanh_f := 1393;
        ELSIF x = 1701 THEN
            tanh_f := 1393;
        ELSIF x = 1702 THEN
            tanh_f := 1394;
        ELSIF x = 1703 THEN
            tanh_f := 1394;
        ELSIF x = 1704 THEN
            tanh_f := 1395;
        ELSIF x = 1705 THEN
            tanh_f := 1395;
        ELSIF x = 1706 THEN
            tanh_f := 1396;
        ELSIF x = 1707 THEN
            tanh_f := 1396;
        ELSIF x = 1708 THEN
            tanh_f := 1397;
        ELSIF x = 1709 THEN
            tanh_f := 1397;
        ELSIF x = 1710 THEN
            tanh_f := 1398;
        ELSIF x = 1711 THEN
            tanh_f := 1399;
        ELSIF x = 1712 THEN
            tanh_f := 1399;
        ELSIF x = 1713 THEN
            tanh_f := 1400;
        ELSIF x = 1714 THEN
            tanh_f := 1400;
        ELSIF x = 1715 THEN
            tanh_f := 1401;
        ELSIF x = 1716 THEN
            tanh_f := 1401;
        ELSIF x = 1717 THEN
            tanh_f := 1402;
        ELSIF x = 1718 THEN
            tanh_f := 1402;
        ELSIF x = 1719 THEN
            tanh_f := 1403;
        ELSIF x = 1720 THEN
            tanh_f := 1403;
        ELSIF x = 1721 THEN
            tanh_f := 1404;
        ELSIF x = 1722 THEN
            tanh_f := 1405;
        ELSIF x = 1723 THEN
            tanh_f := 1405;
        ELSIF x = 1724 THEN
            tanh_f := 1406;
        ELSIF x = 1725 THEN
            tanh_f := 1406;
        ELSIF x = 1726 THEN
            tanh_f := 1407;
        ELSIF x = 1727 THEN
            tanh_f := 1407;
        ELSIF x = 1728 THEN
            tanh_f := 1408;
        ELSIF x = 1729 THEN
            tanh_f := 1408;
        ELSIF x = 1730 THEN
            tanh_f := 1409;
        ELSIF x = 1731 THEN
            tanh_f := 1410;
        ELSIF x = 1732 THEN
            tanh_f := 1410;
        ELSIF x = 1733 THEN
            tanh_f := 1411;
        ELSIF x = 1734 THEN
            tanh_f := 1411;
        ELSIF x = 1735 THEN
            tanh_f := 1412;
        ELSIF x = 1736 THEN
            tanh_f := 1412;
        ELSIF x = 1737 THEN
            tanh_f := 1413;
        ELSIF x = 1738 THEN
            tanh_f := 1413;
        ELSIF x = 1739 THEN
            tanh_f := 1414;
        ELSIF x = 1740 THEN
            tanh_f := 1414;
        ELSIF x = 1741 THEN
            tanh_f := 1415;
        ELSIF x = 1742 THEN
            tanh_f := 1416;
        ELSIF x = 1743 THEN
            tanh_f := 1416;
        ELSIF x = 1744 THEN
            tanh_f := 1417;
        ELSIF x = 1745 THEN
            tanh_f := 1417;
        ELSIF x = 1746 THEN
            tanh_f := 1418;
        ELSIF x = 1747 THEN
            tanh_f := 1418;
        ELSIF x = 1748 THEN
            tanh_f := 1419;
        ELSIF x = 1749 THEN
            tanh_f := 1419;
        ELSIF x = 1750 THEN
            tanh_f := 1420;
        ELSIF x = 1751 THEN
            tanh_f := 1420;
        ELSIF x = 1752 THEN
            tanh_f := 1421;
        ELSIF x = 1753 THEN
            tanh_f := 1422;
        ELSIF x = 1754 THEN
            tanh_f := 1422;
        ELSIF x = 1755 THEN
            tanh_f := 1423;
        ELSIF x = 1756 THEN
            tanh_f := 1423;
        ELSIF x = 1757 THEN
            tanh_f := 1424;
        ELSIF x = 1758 THEN
            tanh_f := 1424;
        ELSIF x = 1759 THEN
            tanh_f := 1425;
        ELSIF x = 1760 THEN
            tanh_f := 1425;
        ELSIF x = 1761 THEN
            tanh_f := 1426;
        ELSIF x = 1762 THEN
            tanh_f := 1427;
        ELSIF x = 1763 THEN
            tanh_f := 1427;
        ELSIF x = 1764 THEN
            tanh_f := 1428;
        ELSIF x = 1765 THEN
            tanh_f := 1428;
        ELSIF x = 1766 THEN
            tanh_f := 1429;
        ELSIF x = 1767 THEN
            tanh_f := 1429;
        ELSIF x = 1768 THEN
            tanh_f := 1430;
        ELSIF x = 1769 THEN
            tanh_f := 1430;
        ELSIF x = 1770 THEN
            tanh_f := 1431;
        ELSIF x = 1771 THEN
            tanh_f := 1431;
        ELSIF x = 1772 THEN
            tanh_f := 1432;
        ELSIF x = 1773 THEN
            tanh_f := 1433;
        ELSIF x = 1774 THEN
            tanh_f := 1433;
        ELSIF x = 1775 THEN
            tanh_f := 1434;
        ELSIF x = 1776 THEN
            tanh_f := 1434;
        ELSIF x = 1777 THEN
            tanh_f := 1435;
        ELSIF x = 1778 THEN
            tanh_f := 1435;
        ELSIF x = 1779 THEN
            tanh_f := 1436;
        ELSIF x = 1780 THEN
            tanh_f := 1436;
        ELSIF x = 1781 THEN
            tanh_f := 1437;
        ELSIF x = 1782 THEN
            tanh_f := 1438;
        ELSIF x = 1783 THEN
            tanh_f := 1438;
        ELSIF x = 1784 THEN
            tanh_f := 1439;
        ELSIF x = 1785 THEN
            tanh_f := 1439;
        ELSIF x = 1786 THEN
            tanh_f := 1440;
        ELSIF x = 1787 THEN
            tanh_f := 1440;
        ELSIF x = 1788 THEN
            tanh_f := 1441;
        ELSIF x = 1789 THEN
            tanh_f := 1441;
        ELSIF x = 1790 THEN
            tanh_f := 1442;
        ELSIF x = 1791 THEN
            tanh_f := 1442;
        ELSIF x = 1792 THEN
            tanh_f := 1443;
        ELSIF x = 1793 THEN
            tanh_f := 1443;
        ELSIF x = 1794 THEN
            tanh_f := 1443;
        ELSIF x = 1795 THEN
            tanh_f := 1444;
        ELSIF x = 1796 THEN
            tanh_f := 1444;
        ELSIF x = 1797 THEN
            tanh_f := 1445;
        ELSIF x = 1798 THEN
            tanh_f := 1445;
        ELSIF x = 1799 THEN
            tanh_f := 1446;
        ELSIF x = 1800 THEN
            tanh_f := 1446;
        ELSIF x = 1801 THEN
            tanh_f := 1447;
        ELSIF x = 1802 THEN
            tanh_f := 1447;
        ELSIF x = 1803 THEN
            tanh_f := 1448;
        ELSIF x = 1804 THEN
            tanh_f := 1448;
        ELSIF x = 1805 THEN
            tanh_f := 1449;
        ELSIF x = 1806 THEN
            tanh_f := 1449;
        ELSIF x = 1807 THEN
            tanh_f := 1449;
        ELSIF x = 1808 THEN
            tanh_f := 1450;
        ELSIF x = 1809 THEN
            tanh_f := 1450;
        ELSIF x = 1810 THEN
            tanh_f := 1451;
        ELSIF x = 1811 THEN
            tanh_f := 1451;
        ELSIF x = 1812 THEN
            tanh_f := 1452;
        ELSIF x = 1813 THEN
            tanh_f := 1452;
        ELSIF x = 1814 THEN
            tanh_f := 1453;
        ELSIF x = 1815 THEN
            tanh_f := 1453;
        ELSIF x = 1816 THEN
            tanh_f := 1454;
        ELSIF x = 1817 THEN
            tanh_f := 1454;
        ELSIF x = 1818 THEN
            tanh_f := 1455;
        ELSIF x = 1819 THEN
            tanh_f := 1455;
        ELSIF x = 1820 THEN
            tanh_f := 1456;
        ELSIF x = 1821 THEN
            tanh_f := 1456;
        ELSIF x = 1822 THEN
            tanh_f := 1456;
        ELSIF x = 1823 THEN
            tanh_f := 1457;
        ELSIF x = 1824 THEN
            tanh_f := 1457;
        ELSIF x = 1825 THEN
            tanh_f := 1458;
        ELSIF x = 1826 THEN
            tanh_f := 1458;
        ELSIF x = 1827 THEN
            tanh_f := 1459;
        ELSIF x = 1828 THEN
            tanh_f := 1459;
        ELSIF x = 1829 THEN
            tanh_f := 1460;
        ELSIF x = 1830 THEN
            tanh_f := 1460;
        ELSIF x = 1831 THEN
            tanh_f := 1461;
        ELSIF x = 1832 THEN
            tanh_f := 1461;
        ELSIF x = 1833 THEN
            tanh_f := 1462;
        ELSIF x = 1834 THEN
            tanh_f := 1462;
        ELSIF x = 1835 THEN
            tanh_f := 1462;
        ELSIF x = 1836 THEN
            tanh_f := 1463;
        ELSIF x = 1837 THEN
            tanh_f := 1463;
        ELSIF x = 1838 THEN
            tanh_f := 1464;
        ELSIF x = 1839 THEN
            tanh_f := 1464;
        ELSIF x = 1840 THEN
            tanh_f := 1465;
        ELSIF x = 1841 THEN
            tanh_f := 1465;
        ELSIF x = 1842 THEN
            tanh_f := 1466;
        ELSIF x = 1843 THEN
            tanh_f := 1466;
        ELSIF x = 1844 THEN
            tanh_f := 1467;
        ELSIF x = 1845 THEN
            tanh_f := 1467;
        ELSIF x = 1846 THEN
            tanh_f := 1468;
        ELSIF x = 1847 THEN
            tanh_f := 1468;
        ELSIF x = 1848 THEN
            tanh_f := 1469;
        ELSIF x = 1849 THEN
            tanh_f := 1469;
        ELSIF x = 1850 THEN
            tanh_f := 1469;
        ELSIF x = 1851 THEN
            tanh_f := 1470;
        ELSIF x = 1852 THEN
            tanh_f := 1470;
        ELSIF x = 1853 THEN
            tanh_f := 1471;
        ELSIF x = 1854 THEN
            tanh_f := 1471;
        ELSIF x = 1855 THEN
            tanh_f := 1472;
        ELSIF x = 1856 THEN
            tanh_f := 1472;
        ELSIF x = 1857 THEN
            tanh_f := 1473;
        ELSIF x = 1858 THEN
            tanh_f := 1473;
        ELSIF x = 1859 THEN
            tanh_f := 1474;
        ELSIF x = 1860 THEN
            tanh_f := 1474;
        ELSIF x = 1861 THEN
            tanh_f := 1475;
        ELSIF x = 1862 THEN
            tanh_f := 1475;
        ELSIF x = 1863 THEN
            tanh_f := 1476;
        ELSIF x = 1864 THEN
            tanh_f := 1476;
        ELSIF x = 1865 THEN
            tanh_f := 1476;
        ELSIF x = 1866 THEN
            tanh_f := 1477;
        ELSIF x = 1867 THEN
            tanh_f := 1477;
        ELSIF x = 1868 THEN
            tanh_f := 1478;
        ELSIF x = 1869 THEN
            tanh_f := 1478;
        ELSIF x = 1870 THEN
            tanh_f := 1479;
        ELSIF x = 1871 THEN
            tanh_f := 1479;
        ELSIF x = 1872 THEN
            tanh_f := 1480;
        ELSIF x = 1873 THEN
            tanh_f := 1480;
        ELSIF x = 1874 THEN
            tanh_f := 1481;
        ELSIF x = 1875 THEN
            tanh_f := 1481;
        ELSIF x = 1876 THEN
            tanh_f := 1482;
        ELSIF x = 1877 THEN
            tanh_f := 1482;
        ELSIF x = 1878 THEN
            tanh_f := 1482;
        ELSIF x = 1879 THEN
            tanh_f := 1483;
        ELSIF x = 1880 THEN
            tanh_f := 1483;
        ELSIF x = 1881 THEN
            tanh_f := 1484;
        ELSIF x = 1882 THEN
            tanh_f := 1484;
        ELSIF x = 1883 THEN
            tanh_f := 1485;
        ELSIF x = 1884 THEN
            tanh_f := 1485;
        ELSIF x = 1885 THEN
            tanh_f := 1486;
        ELSIF x = 1886 THEN
            tanh_f := 1486;
        ELSIF x = 1887 THEN
            tanh_f := 1487;
        ELSIF x = 1888 THEN
            tanh_f := 1487;
        ELSIF x = 1889 THEN
            tanh_f := 1488;
        ELSIF x = 1890 THEN
            tanh_f := 1488;
        ELSIF x = 1891 THEN
            tanh_f := 1489;
        ELSIF x = 1892 THEN
            tanh_f := 1489;
        ELSIF x = 1893 THEN
            tanh_f := 1489;
        ELSIF x = 1894 THEN
            tanh_f := 1490;
        ELSIF x = 1895 THEN
            tanh_f := 1490;
        ELSIF x = 1896 THEN
            tanh_f := 1491;
        ELSIF x = 1897 THEN
            tanh_f := 1491;
        ELSIF x = 1898 THEN
            tanh_f := 1492;
        ELSIF x = 1899 THEN
            tanh_f := 1492;
        ELSIF x = 1900 THEN
            tanh_f := 1493;
        ELSIF x = 1901 THEN
            tanh_f := 1493;
        ELSIF x = 1902 THEN
            tanh_f := 1494;
        ELSIF x = 1903 THEN
            tanh_f := 1494;
        ELSIF x = 1904 THEN
            tanh_f := 1495;
        ELSIF x = 1905 THEN
            tanh_f := 1495;
        ELSIF x = 1906 THEN
            tanh_f := 1495;
        ELSIF x = 1907 THEN
            tanh_f := 1496;
        ELSIF x = 1908 THEN
            tanh_f := 1496;
        ELSIF x = 1909 THEN
            tanh_f := 1497;
        ELSIF x = 1910 THEN
            tanh_f := 1497;
        ELSIF x = 1911 THEN
            tanh_f := 1498;
        ELSIF x = 1912 THEN
            tanh_f := 1498;
        ELSIF x = 1913 THEN
            tanh_f := 1499;
        ELSIF x = 1914 THEN
            tanh_f := 1499;
        ELSIF x = 1915 THEN
            tanh_f := 1500;
        ELSIF x = 1916 THEN
            tanh_f := 1500;
        ELSIF x = 1917 THEN
            tanh_f := 1501;
        ELSIF x = 1918 THEN
            tanh_f := 1501;
        ELSIF x = 1919 THEN
            tanh_f := 1502;
        ELSIF x = 1920 THEN
            tanh_f := 1502;
        ELSIF x = 1921 THEN
            tanh_f := 1502;
        ELSIF x = 1922 THEN
            tanh_f := 1503;
        ELSIF x = 1923 THEN
            tanh_f := 1503;
        ELSIF x = 1924 THEN
            tanh_f := 1504;
        ELSIF x = 1925 THEN
            tanh_f := 1504;
        ELSIF x = 1926 THEN
            tanh_f := 1505;
        ELSIF x = 1927 THEN
            tanh_f := 1505;
        ELSIF x = 1928 THEN
            tanh_f := 1506;
        ELSIF x = 1929 THEN
            tanh_f := 1506;
        ELSIF x = 1930 THEN
            tanh_f := 1507;
        ELSIF x = 1931 THEN
            tanh_f := 1507;
        ELSIF x = 1932 THEN
            tanh_f := 1508;
        ELSIF x = 1933 THEN
            tanh_f := 1508;
        ELSIF x = 1934 THEN
            tanh_f := 1509;
        ELSIF x = 1935 THEN
            tanh_f := 1509;
        ELSIF x = 1936 THEN
            tanh_f := 1509;
        ELSIF x = 1937 THEN
            tanh_f := 1510;
        ELSIF x = 1938 THEN
            tanh_f := 1510;
        ELSIF x = 1939 THEN
            tanh_f := 1511;
        ELSIF x = 1940 THEN
            tanh_f := 1511;
        ELSIF x = 1941 THEN
            tanh_f := 1512;
        ELSIF x = 1942 THEN
            tanh_f := 1512;
        ELSIF x = 1943 THEN
            tanh_f := 1513;
        ELSIF x = 1944 THEN
            tanh_f := 1513;
        ELSIF x = 1945 THEN
            tanh_f := 1514;
        ELSIF x = 1946 THEN
            tanh_f := 1514;
        ELSIF x = 1947 THEN
            tanh_f := 1515;
        ELSIF x = 1948 THEN
            tanh_f := 1515;
        ELSIF x = 1949 THEN
            tanh_f := 1515;
        ELSIF x = 1950 THEN
            tanh_f := 1516;
        ELSIF x = 1951 THEN
            tanh_f := 1516;
        ELSIF x = 1952 THEN
            tanh_f := 1517;
        ELSIF x = 1953 THEN
            tanh_f := 1517;
        ELSIF x = 1954 THEN
            tanh_f := 1518;
        ELSIF x = 1955 THEN
            tanh_f := 1518;
        ELSIF x = 1956 THEN
            tanh_f := 1519;
        ELSIF x = 1957 THEN
            tanh_f := 1519;
        ELSIF x = 1958 THEN
            tanh_f := 1520;
        ELSIF x = 1959 THEN
            tanh_f := 1520;
        ELSIF x = 1960 THEN
            tanh_f := 1521;
        ELSIF x = 1961 THEN
            tanh_f := 1521;
        ELSIF x = 1962 THEN
            tanh_f := 1522;
        ELSIF x = 1963 THEN
            tanh_f := 1522;
        ELSIF x = 1964 THEN
            tanh_f := 1522;
        ELSIF x = 1965 THEN
            tanh_f := 1523;
        ELSIF x = 1966 THEN
            tanh_f := 1523;
        ELSIF x = 1967 THEN
            tanh_f := 1524;
        ELSIF x = 1968 THEN
            tanh_f := 1524;
        ELSIF x = 1969 THEN
            tanh_f := 1525;
        ELSIF x = 1970 THEN
            tanh_f := 1525;
        ELSIF x = 1971 THEN
            tanh_f := 1526;
        ELSIF x = 1972 THEN
            tanh_f := 1526;
        ELSIF x = 1973 THEN
            tanh_f := 1527;
        ELSIF x = 1974 THEN
            tanh_f := 1527;
        ELSIF x = 1975 THEN
            tanh_f := 1528;
        ELSIF x = 1976 THEN
            tanh_f := 1528;
        ELSIF x = 1977 THEN
            tanh_f := 1528;
        ELSIF x = 1978 THEN
            tanh_f := 1529;
        ELSIF x = 1979 THEN
            tanh_f := 1529;
        ELSIF x = 1980 THEN
            tanh_f := 1530;
        ELSIF x = 1981 THEN
            tanh_f := 1530;
        ELSIF x = 1982 THEN
            tanh_f := 1531;
        ELSIF x = 1983 THEN
            tanh_f := 1531;
        ELSIF x = 1984 THEN
            tanh_f := 1532;
        ELSIF x = 1985 THEN
            tanh_f := 1532;
        ELSIF x = 1986 THEN
            tanh_f := 1533;
        ELSIF x = 1987 THEN
            tanh_f := 1533;
        ELSIF x = 1988 THEN
            tanh_f := 1534;
        ELSIF x = 1989 THEN
            tanh_f := 1534;
        ELSIF x = 1990 THEN
            tanh_f := 1535;
        ELSIF x = 1991 THEN
            tanh_f := 1535;
        ELSIF x = 1992 THEN
            tanh_f := 1535;
        ELSIF x = 1993 THEN
            tanh_f := 1536;
        ELSIF x = 1994 THEN
            tanh_f := 1536;
        ELSIF x = 1995 THEN
            tanh_f := 1537;
        ELSIF x = 1996 THEN
            tanh_f := 1537;
        ELSIF x = 1997 THEN
            tanh_f := 1538;
        ELSIF x = 1998 THEN
            tanh_f := 1538;
        ELSIF x = 1999 THEN
            tanh_f := 1539;
        ELSIF x = 2000 THEN
            tanh_f := 1539;
        ELSIF x = 2001 THEN
            tanh_f := 1540;
        ELSIF x = 2002 THEN
            tanh_f := 1540;
        ELSIF x = 2003 THEN
            tanh_f := 1541;
        ELSIF x = 2004 THEN
            tanh_f := 1541;
        ELSIF x = 2005 THEN
            tanh_f := 1542;
        ELSIF x = 2006 THEN
            tanh_f := 1542;
        ELSIF x = 2007 THEN
            tanh_f := 1542;
        ELSIF x = 2008 THEN
            tanh_f := 1543;
        ELSIF x = 2009 THEN
            tanh_f := 1543;
        ELSIF x = 2010 THEN
            tanh_f := 1544;
        ELSIF x = 2011 THEN
            tanh_f := 1544;
        ELSIF x = 2012 THEN
            tanh_f := 1545;
        ELSIF x = 2013 THEN
            tanh_f := 1545;
        ELSIF x = 2014 THEN
            tanh_f := 1546;
        ELSIF x = 2015 THEN
            tanh_f := 1546;
        ELSIF x = 2016 THEN
            tanh_f := 1547;
        ELSIF x = 2017 THEN
            tanh_f := 1547;
        ELSIF x = 2018 THEN
            tanh_f := 1548;
        ELSIF x = 2019 THEN
            tanh_f := 1548;
        ELSIF x = 2020 THEN
            tanh_f := 1548;
        ELSIF x = 2021 THEN
            tanh_f := 1549;
        ELSIF x = 2022 THEN
            tanh_f := 1549;
        ELSIF x = 2023 THEN
            tanh_f := 1550;
        ELSIF x = 2024 THEN
            tanh_f := 1550;
        ELSIF x = 2025 THEN
            tanh_f := 1551;
        ELSIF x = 2026 THEN
            tanh_f := 1551;
        ELSIF x = 2027 THEN
            tanh_f := 1552;
        ELSIF x = 2028 THEN
            tanh_f := 1552;
        ELSIF x = 2029 THEN
            tanh_f := 1553;
        ELSIF x = 2030 THEN
            tanh_f := 1553;
        ELSIF x = 2031 THEN
            tanh_f := 1554;
        ELSIF x = 2032 THEN
            tanh_f := 1554;
        ELSIF x = 2033 THEN
            tanh_f := 1555;
        ELSIF x = 2034 THEN
            tanh_f := 1555;
        ELSIF x = 2035 THEN
            tanh_f := 1555;
        ELSIF x = 2036 THEN
            tanh_f := 1556;
        ELSIF x = 2037 THEN
            tanh_f := 1556;
        ELSIF x = 2038 THEN
            tanh_f := 1557;
        ELSIF x = 2039 THEN
            tanh_f := 1557;
        ELSIF x = 2040 THEN
            tanh_f := 1558;
        ELSIF x = 2041 THEN
            tanh_f := 1558;
        ELSIF x = 2042 THEN
            tanh_f := 1559;
        ELSIF x = 2043 THEN
            tanh_f := 1559;
        ELSIF x = 2044 THEN
            tanh_f := 1560;
        ELSIF x = 2045 THEN
            tanh_f := 1560;
        ELSIF x = 2046 THEN
            tanh_f := 1561;
        ELSIF x = 2047 THEN
            tanh_f := 1561;
        ELSIF x = 2048 THEN
            tanh_f := 1562;
        ELSIF x = 2049 THEN
            tanh_f := 1562;
        ELSIF x = 2050 THEN
            tanh_f := 1562;
        ELSIF x = 2051 THEN
            tanh_f := 1563;
        ELSIF x = 2052 THEN
            tanh_f := 1563;
        ELSIF x = 2053 THEN
            tanh_f := 1563;
        ELSIF x = 2054 THEN
            tanh_f := 1564;
        ELSIF x = 2055 THEN
            tanh_f := 1564;
        ELSIF x = 2056 THEN
            tanh_f := 1565;
        ELSIF x = 2057 THEN
            tanh_f := 1565;
        ELSIF x = 2058 THEN
            tanh_f := 1565;
        ELSIF x = 2059 THEN
            tanh_f := 1566;
        ELSIF x = 2060 THEN
            tanh_f := 1566;
        ELSIF x = 2061 THEN
            tanh_f := 1566;
        ELSIF x = 2062 THEN
            tanh_f := 1567;
        ELSIF x = 2063 THEN
            tanh_f := 1567;
        ELSIF x = 2064 THEN
            tanh_f := 1568;
        ELSIF x = 2065 THEN
            tanh_f := 1568;
        ELSIF x = 2066 THEN
            tanh_f := 1568;
        ELSIF x = 2067 THEN
            tanh_f := 1569;
        ELSIF x = 2068 THEN
            tanh_f := 1569;
        ELSIF x = 2069 THEN
            tanh_f := 1569;
        ELSIF x = 2070 THEN
            tanh_f := 1570;
        ELSIF x = 2071 THEN
            tanh_f := 1570;
        ELSIF x = 2072 THEN
            tanh_f := 1571;
        ELSIF x = 2073 THEN
            tanh_f := 1571;
        ELSIF x = 2074 THEN
            tanh_f := 1571;
        ELSIF x = 2075 THEN
            tanh_f := 1572;
        ELSIF x = 2076 THEN
            tanh_f := 1572;
        ELSIF x = 2077 THEN
            tanh_f := 1572;
        ELSIF x = 2078 THEN
            tanh_f := 1573;
        ELSIF x = 2079 THEN
            tanh_f := 1573;
        ELSIF x = 2080 THEN
            tanh_f := 1574;
        ELSIF x = 2081 THEN
            tanh_f := 1574;
        ELSIF x = 2082 THEN
            tanh_f := 1574;
        ELSIF x = 2083 THEN
            tanh_f := 1575;
        ELSIF x = 2084 THEN
            tanh_f := 1575;
        ELSIF x = 2085 THEN
            tanh_f := 1575;
        ELSIF x = 2086 THEN
            tanh_f := 1576;
        ELSIF x = 2087 THEN
            tanh_f := 1576;
        ELSIF x = 2088 THEN
            tanh_f := 1577;
        ELSIF x = 2089 THEN
            tanh_f := 1577;
        ELSIF x = 2090 THEN
            tanh_f := 1577;
        ELSIF x = 2091 THEN
            tanh_f := 1578;
        ELSIF x = 2092 THEN
            tanh_f := 1578;
        ELSIF x = 2093 THEN
            tanh_f := 1578;
        ELSIF x = 2094 THEN
            tanh_f := 1579;
        ELSIF x = 2095 THEN
            tanh_f := 1579;
        ELSIF x = 2096 THEN
            tanh_f := 1580;
        ELSIF x = 2097 THEN
            tanh_f := 1580;
        ELSIF x = 2098 THEN
            tanh_f := 1580;
        ELSIF x = 2099 THEN
            tanh_f := 1581;
        ELSIF x = 2100 THEN
            tanh_f := 1581;
        ELSIF x = 2101 THEN
            tanh_f := 1581;
        ELSIF x = 2102 THEN
            tanh_f := 1582;
        ELSIF x = 2103 THEN
            tanh_f := 1582;
        ELSIF x = 2104 THEN
            tanh_f := 1583;
        ELSIF x = 2105 THEN
            tanh_f := 1583;
        ELSIF x = 2106 THEN
            tanh_f := 1583;
        ELSIF x = 2107 THEN
            tanh_f := 1584;
        ELSIF x = 2108 THEN
            tanh_f := 1584;
        ELSIF x = 2109 THEN
            tanh_f := 1584;
        ELSIF x = 2110 THEN
            tanh_f := 1585;
        ELSIF x = 2111 THEN
            tanh_f := 1585;
        ELSIF x = 2112 THEN
            tanh_f := 1586;
        ELSIF x = 2113 THEN
            tanh_f := 1586;
        ELSIF x = 2114 THEN
            tanh_f := 1586;
        ELSIF x = 2115 THEN
            tanh_f := 1587;
        ELSIF x = 2116 THEN
            tanh_f := 1587;
        ELSIF x = 2117 THEN
            tanh_f := 1588;
        ELSIF x = 2118 THEN
            tanh_f := 1588;
        ELSIF x = 2119 THEN
            tanh_f := 1588;
        ELSIF x = 2120 THEN
            tanh_f := 1589;
        ELSIF x = 2121 THEN
            tanh_f := 1589;
        ELSIF x = 2122 THEN
            tanh_f := 1589;
        ELSIF x = 2123 THEN
            tanh_f := 1590;
        ELSIF x = 2124 THEN
            tanh_f := 1590;
        ELSIF x = 2125 THEN
            tanh_f := 1591;
        ELSIF x = 2126 THEN
            tanh_f := 1591;
        ELSIF x = 2127 THEN
            tanh_f := 1591;
        ELSIF x = 2128 THEN
            tanh_f := 1592;
        ELSIF x = 2129 THEN
            tanh_f := 1592;
        ELSIF x = 2130 THEN
            tanh_f := 1592;
        ELSIF x = 2131 THEN
            tanh_f := 1593;
        ELSIF x = 2132 THEN
            tanh_f := 1593;
        ELSIF x = 2133 THEN
            tanh_f := 1594;
        ELSIF x = 2134 THEN
            tanh_f := 1594;
        ELSIF x = 2135 THEN
            tanh_f := 1594;
        ELSIF x = 2136 THEN
            tanh_f := 1595;
        ELSIF x = 2137 THEN
            tanh_f := 1595;
        ELSIF x = 2138 THEN
            tanh_f := 1595;
        ELSIF x = 2139 THEN
            tanh_f := 1596;
        ELSIF x = 2140 THEN
            tanh_f := 1596;
        ELSIF x = 2141 THEN
            tanh_f := 1597;
        ELSIF x = 2142 THEN
            tanh_f := 1597;
        ELSIF x = 2143 THEN
            tanh_f := 1597;
        ELSIF x = 2144 THEN
            tanh_f := 1598;
        ELSIF x = 2145 THEN
            tanh_f := 1598;
        ELSIF x = 2146 THEN
            tanh_f := 1598;
        ELSIF x = 2147 THEN
            tanh_f := 1599;
        ELSIF x = 2148 THEN
            tanh_f := 1599;
        ELSIF x = 2149 THEN
            tanh_f := 1600;
        ELSIF x = 2150 THEN
            tanh_f := 1600;
        ELSIF x = 2151 THEN
            tanh_f := 1600;
        ELSIF x = 2152 THEN
            tanh_f := 1601;
        ELSIF x = 2153 THEN
            tanh_f := 1601;
        ELSIF x = 2154 THEN
            tanh_f := 1601;
        ELSIF x = 2155 THEN
            tanh_f := 1602;
        ELSIF x = 2156 THEN
            tanh_f := 1602;
        ELSIF x = 2157 THEN
            tanh_f := 1603;
        ELSIF x = 2158 THEN
            tanh_f := 1603;
        ELSIF x = 2159 THEN
            tanh_f := 1603;
        ELSIF x = 2160 THEN
            tanh_f := 1604;
        ELSIF x = 2161 THEN
            tanh_f := 1604;
        ELSIF x = 2162 THEN
            tanh_f := 1604;
        ELSIF x = 2163 THEN
            tanh_f := 1605;
        ELSIF x = 2164 THEN
            tanh_f := 1605;
        ELSIF x = 2165 THEN
            tanh_f := 1606;
        ELSIF x = 2166 THEN
            tanh_f := 1606;
        ELSIF x = 2167 THEN
            tanh_f := 1606;
        ELSIF x = 2168 THEN
            tanh_f := 1607;
        ELSIF x = 2169 THEN
            tanh_f := 1607;
        ELSIF x = 2170 THEN
            tanh_f := 1607;
        ELSIF x = 2171 THEN
            tanh_f := 1608;
        ELSIF x = 2172 THEN
            tanh_f := 1608;
        ELSIF x = 2173 THEN
            tanh_f := 1609;
        ELSIF x = 2174 THEN
            tanh_f := 1609;
        ELSIF x = 2175 THEN
            tanh_f := 1609;
        ELSIF x = 2176 THEN
            tanh_f := 1610;
        ELSIF x = 2177 THEN
            tanh_f := 1610;
        ELSIF x = 2178 THEN
            tanh_f := 1611;
        ELSIF x = 2179 THEN
            tanh_f := 1611;
        ELSIF x = 2180 THEN
            tanh_f := 1611;
        ELSIF x = 2181 THEN
            tanh_f := 1612;
        ELSIF x = 2182 THEN
            tanh_f := 1612;
        ELSIF x = 2183 THEN
            tanh_f := 1612;
        ELSIF x = 2184 THEN
            tanh_f := 1613;
        ELSIF x = 2185 THEN
            tanh_f := 1613;
        ELSIF x = 2186 THEN
            tanh_f := 1614;
        ELSIF x = 2187 THEN
            tanh_f := 1614;
        ELSIF x = 2188 THEN
            tanh_f := 1614;
        ELSIF x = 2189 THEN
            tanh_f := 1615;
        ELSIF x = 2190 THEN
            tanh_f := 1615;
        ELSIF x = 2191 THEN
            tanh_f := 1615;
        ELSIF x = 2192 THEN
            tanh_f := 1616;
        ELSIF x = 2193 THEN
            tanh_f := 1616;
        ELSIF x = 2194 THEN
            tanh_f := 1617;
        ELSIF x = 2195 THEN
            tanh_f := 1617;
        ELSIF x = 2196 THEN
            tanh_f := 1617;
        ELSIF x = 2197 THEN
            tanh_f := 1618;
        ELSIF x = 2198 THEN
            tanh_f := 1618;
        ELSIF x = 2199 THEN
            tanh_f := 1618;
        ELSIF x = 2200 THEN
            tanh_f := 1619;
        ELSIF x = 2201 THEN
            tanh_f := 1619;
        ELSIF x = 2202 THEN
            tanh_f := 1620;
        ELSIF x = 2203 THEN
            tanh_f := 1620;
        ELSIF x = 2204 THEN
            tanh_f := 1620;
        ELSIF x = 2205 THEN
            tanh_f := 1621;
        ELSIF x = 2206 THEN
            tanh_f := 1621;
        ELSIF x = 2207 THEN
            tanh_f := 1621;
        ELSIF x = 2208 THEN
            tanh_f := 1622;
        ELSIF x = 2209 THEN
            tanh_f := 1622;
        ELSIF x = 2210 THEN
            tanh_f := 1623;
        ELSIF x = 2211 THEN
            tanh_f := 1623;
        ELSIF x = 2212 THEN
            tanh_f := 1623;
        ELSIF x = 2213 THEN
            tanh_f := 1624;
        ELSIF x = 2214 THEN
            tanh_f := 1624;
        ELSIF x = 2215 THEN
            tanh_f := 1624;
        ELSIF x = 2216 THEN
            tanh_f := 1625;
        ELSIF x = 2217 THEN
            tanh_f := 1625;
        ELSIF x = 2218 THEN
            tanh_f := 1626;
        ELSIF x = 2219 THEN
            tanh_f := 1626;
        ELSIF x = 2220 THEN
            tanh_f := 1626;
        ELSIF x = 2221 THEN
            tanh_f := 1627;
        ELSIF x = 2222 THEN
            tanh_f := 1627;
        ELSIF x = 2223 THEN
            tanh_f := 1627;
        ELSIF x = 2224 THEN
            tanh_f := 1628;
        ELSIF x = 2225 THEN
            tanh_f := 1628;
        ELSIF x = 2226 THEN
            tanh_f := 1629;
        ELSIF x = 2227 THEN
            tanh_f := 1629;
        ELSIF x = 2228 THEN
            tanh_f := 1629;
        ELSIF x = 2229 THEN
            tanh_f := 1630;
        ELSIF x = 2230 THEN
            tanh_f := 1630;
        ELSIF x = 2231 THEN
            tanh_f := 1630;
        ELSIF x = 2232 THEN
            tanh_f := 1631;
        ELSIF x = 2233 THEN
            tanh_f := 1631;
        ELSIF x = 2234 THEN
            tanh_f := 1632;
        ELSIF x = 2235 THEN
            tanh_f := 1632;
        ELSIF x = 2236 THEN
            tanh_f := 1632;
        ELSIF x = 2237 THEN
            tanh_f := 1633;
        ELSIF x = 2238 THEN
            tanh_f := 1633;
        ELSIF x = 2239 THEN
            tanh_f := 1633;
        ELSIF x = 2240 THEN
            tanh_f := 1634;
        ELSIF x = 2241 THEN
            tanh_f := 1634;
        ELSIF x = 2242 THEN
            tanh_f := 1635;
        ELSIF x = 2243 THEN
            tanh_f := 1635;
        ELSIF x = 2244 THEN
            tanh_f := 1635;
        ELSIF x = 2245 THEN
            tanh_f := 1636;
        ELSIF x = 2246 THEN
            tanh_f := 1636;
        ELSIF x = 2247 THEN
            tanh_f := 1637;
        ELSIF x = 2248 THEN
            tanh_f := 1637;
        ELSIF x = 2249 THEN
            tanh_f := 1637;
        ELSIF x = 2250 THEN
            tanh_f := 1638;
        ELSIF x = 2251 THEN
            tanh_f := 1638;
        ELSIF x = 2252 THEN
            tanh_f := 1638;
        ELSIF x = 2253 THEN
            tanh_f := 1639;
        ELSIF x = 2254 THEN
            tanh_f := 1639;
        ELSIF x = 2255 THEN
            tanh_f := 1640;
        ELSIF x = 2256 THEN
            tanh_f := 1640;
        ELSIF x = 2257 THEN
            tanh_f := 1640;
        ELSIF x = 2258 THEN
            tanh_f := 1641;
        ELSIF x = 2259 THEN
            tanh_f := 1641;
        ELSIF x = 2260 THEN
            tanh_f := 1641;
        ELSIF x = 2261 THEN
            tanh_f := 1642;
        ELSIF x = 2262 THEN
            tanh_f := 1642;
        ELSIF x = 2263 THEN
            tanh_f := 1643;
        ELSIF x = 2264 THEN
            tanh_f := 1643;
        ELSIF x = 2265 THEN
            tanh_f := 1643;
        ELSIF x = 2266 THEN
            tanh_f := 1644;
        ELSIF x = 2267 THEN
            tanh_f := 1644;
        ELSIF x = 2268 THEN
            tanh_f := 1644;
        ELSIF x = 2269 THEN
            tanh_f := 1645;
        ELSIF x = 2270 THEN
            tanh_f := 1645;
        ELSIF x = 2271 THEN
            tanh_f := 1646;
        ELSIF x = 2272 THEN
            tanh_f := 1646;
        ELSIF x = 2273 THEN
            tanh_f := 1646;
        ELSIF x = 2274 THEN
            tanh_f := 1647;
        ELSIF x = 2275 THEN
            tanh_f := 1647;
        ELSIF x = 2276 THEN
            tanh_f := 1647;
        ELSIF x = 2277 THEN
            tanh_f := 1648;
        ELSIF x = 2278 THEN
            tanh_f := 1648;
        ELSIF x = 2279 THEN
            tanh_f := 1649;
        ELSIF x = 2280 THEN
            tanh_f := 1649;
        ELSIF x = 2281 THEN
            tanh_f := 1649;
        ELSIF x = 2282 THEN
            tanh_f := 1650;
        ELSIF x = 2283 THEN
            tanh_f := 1650;
        ELSIF x = 2284 THEN
            tanh_f := 1650;
        ELSIF x = 2285 THEN
            tanh_f := 1651;
        ELSIF x = 2286 THEN
            tanh_f := 1651;
        ELSIF x = 2287 THEN
            tanh_f := 1652;
        ELSIF x = 2288 THEN
            tanh_f := 1652;
        ELSIF x = 2289 THEN
            tanh_f := 1652;
        ELSIF x = 2290 THEN
            tanh_f := 1653;
        ELSIF x = 2291 THEN
            tanh_f := 1653;
        ELSIF x = 2292 THEN
            tanh_f := 1653;
        ELSIF x = 2293 THEN
            tanh_f := 1654;
        ELSIF x = 2294 THEN
            tanh_f := 1654;
        ELSIF x = 2295 THEN
            tanh_f := 1655;
        ELSIF x = 2296 THEN
            tanh_f := 1655;
        ELSIF x = 2297 THEN
            tanh_f := 1655;
        ELSIF x = 2298 THEN
            tanh_f := 1656;
        ELSIF x = 2299 THEN
            tanh_f := 1656;
        ELSIF x = 2300 THEN
            tanh_f := 1656;
        ELSIF x = 2301 THEN
            tanh_f := 1657;
        ELSIF x = 2302 THEN
            tanh_f := 1657;
        ELSIF x = 2303 THEN
            tanh_f := 1658;
        ELSIF x = 2304 THEN
            tanh_f := 1658;
        ELSIF x = 2305 THEN
            tanh_f := 1658;
        ELSIF x = 2306 THEN
            tanh_f := 1659;
        ELSIF x = 2307 THEN
            tanh_f := 1659;
        ELSIF x = 2308 THEN
            tanh_f := 1659;
        ELSIF x = 2309 THEN
            tanh_f := 1660;
        ELSIF x = 2310 THEN
            tanh_f := 1660;
        ELSIF x = 2311 THEN
            tanh_f := 1660;
        ELSIF x = 2312 THEN
            tanh_f := 1661;
        ELSIF x = 2313 THEN
            tanh_f := 1661;
        ELSIF x = 2314 THEN
            tanh_f := 1661;
        ELSIF x = 2315 THEN
            tanh_f := 1661;
        ELSIF x = 2316 THEN
            tanh_f := 1662;
        ELSIF x = 2317 THEN
            tanh_f := 1662;
        ELSIF x = 2318 THEN
            tanh_f := 1662;
        ELSIF x = 2319 THEN
            tanh_f := 1663;
        ELSIF x = 2320 THEN
            tanh_f := 1663;
        ELSIF x = 2321 THEN
            tanh_f := 1663;
        ELSIF x = 2322 THEN
            tanh_f := 1664;
        ELSIF x = 2323 THEN
            tanh_f := 1664;
        ELSIF x = 2324 THEN
            tanh_f := 1664;
        ELSIF x = 2325 THEN
            tanh_f := 1665;
        ELSIF x = 2326 THEN
            tanh_f := 1665;
        ELSIF x = 2327 THEN
            tanh_f := 1665;
        ELSIF x = 2328 THEN
            tanh_f := 1666;
        ELSIF x = 2329 THEN
            tanh_f := 1666;
        ELSIF x = 2330 THEN
            tanh_f := 1666;
        ELSIF x = 2331 THEN
            tanh_f := 1666;
        ELSIF x = 2332 THEN
            tanh_f := 1667;
        ELSIF x = 2333 THEN
            tanh_f := 1667;
        ELSIF x = 2334 THEN
            tanh_f := 1667;
        ELSIF x = 2335 THEN
            tanh_f := 1668;
        ELSIF x = 2336 THEN
            tanh_f := 1668;
        ELSIF x = 2337 THEN
            tanh_f := 1668;
        ELSIF x = 2338 THEN
            tanh_f := 1669;
        ELSIF x = 2339 THEN
            tanh_f := 1669;
        ELSIF x = 2340 THEN
            tanh_f := 1669;
        ELSIF x = 2341 THEN
            tanh_f := 1670;
        ELSIF x = 2342 THEN
            tanh_f := 1670;
        ELSIF x = 2343 THEN
            tanh_f := 1670;
        ELSIF x = 2344 THEN
            tanh_f := 1671;
        ELSIF x = 2345 THEN
            tanh_f := 1671;
        ELSIF x = 2346 THEN
            tanh_f := 1671;
        ELSIF x = 2347 THEN
            tanh_f := 1672;
        ELSIF x = 2348 THEN
            tanh_f := 1672;
        ELSIF x = 2349 THEN
            tanh_f := 1672;
        ELSIF x = 2350 THEN
            tanh_f := 1672;
        ELSIF x = 2351 THEN
            tanh_f := 1673;
        ELSIF x = 2352 THEN
            tanh_f := 1673;
        ELSIF x = 2353 THEN
            tanh_f := 1673;
        ELSIF x = 2354 THEN
            tanh_f := 1674;
        ELSIF x = 2355 THEN
            tanh_f := 1674;
        ELSIF x = 2356 THEN
            tanh_f := 1674;
        ELSIF x = 2357 THEN
            tanh_f := 1675;
        ELSIF x = 2358 THEN
            tanh_f := 1675;
        ELSIF x = 2359 THEN
            tanh_f := 1675;
        ELSIF x = 2360 THEN
            tanh_f := 1676;
        ELSIF x = 2361 THEN
            tanh_f := 1676;
        ELSIF x = 2362 THEN
            tanh_f := 1676;
        ELSIF x = 2363 THEN
            tanh_f := 1677;
        ELSIF x = 2364 THEN
            tanh_f := 1677;
        ELSIF x = 2365 THEN
            tanh_f := 1677;
        ELSIF x = 2366 THEN
            tanh_f := 1677;
        ELSIF x = 2367 THEN
            tanh_f := 1678;
        ELSIF x = 2368 THEN
            tanh_f := 1678;
        ELSIF x = 2369 THEN
            tanh_f := 1678;
        ELSIF x = 2370 THEN
            tanh_f := 1679;
        ELSIF x = 2371 THEN
            tanh_f := 1679;
        ELSIF x = 2372 THEN
            tanh_f := 1679;
        ELSIF x = 2373 THEN
            tanh_f := 1680;
        ELSIF x = 2374 THEN
            tanh_f := 1680;
        ELSIF x = 2375 THEN
            tanh_f := 1680;
        ELSIF x = 2376 THEN
            tanh_f := 1681;
        ELSIF x = 2377 THEN
            tanh_f := 1681;
        ELSIF x = 2378 THEN
            tanh_f := 1681;
        ELSIF x = 2379 THEN
            tanh_f := 1682;
        ELSIF x = 2380 THEN
            tanh_f := 1682;
        ELSIF x = 2381 THEN
            tanh_f := 1682;
        ELSIF x = 2382 THEN
            tanh_f := 1683;
        ELSIF x = 2383 THEN
            tanh_f := 1683;
        ELSIF x = 2384 THEN
            tanh_f := 1683;
        ELSIF x = 2385 THEN
            tanh_f := 1683;
        ELSIF x = 2386 THEN
            tanh_f := 1684;
        ELSIF x = 2387 THEN
            tanh_f := 1684;
        ELSIF x = 2388 THEN
            tanh_f := 1684;
        ELSIF x = 2389 THEN
            tanh_f := 1685;
        ELSIF x = 2390 THEN
            tanh_f := 1685;
        ELSIF x = 2391 THEN
            tanh_f := 1685;
        ELSIF x = 2392 THEN
            tanh_f := 1686;
        ELSIF x = 2393 THEN
            tanh_f := 1686;
        ELSIF x = 2394 THEN
            tanh_f := 1686;
        ELSIF x = 2395 THEN
            tanh_f := 1687;
        ELSIF x = 2396 THEN
            tanh_f := 1687;
        ELSIF x = 2397 THEN
            tanh_f := 1687;
        ELSIF x = 2398 THEN
            tanh_f := 1688;
        ELSIF x = 2399 THEN
            tanh_f := 1688;
        ELSIF x = 2400 THEN
            tanh_f := 1688;
        ELSIF x = 2401 THEN
            tanh_f := 1689;
        ELSIF x = 2402 THEN
            tanh_f := 1689;
        ELSIF x = 2403 THEN
            tanh_f := 1689;
        ELSIF x = 2404 THEN
            tanh_f := 1689;
        ELSIF x = 2405 THEN
            tanh_f := 1690;
        ELSIF x = 2406 THEN
            tanh_f := 1690;
        ELSIF x = 2407 THEN
            tanh_f := 1690;
        ELSIF x = 2408 THEN
            tanh_f := 1691;
        ELSIF x = 2409 THEN
            tanh_f := 1691;
        ELSIF x = 2410 THEN
            tanh_f := 1691;
        ELSIF x = 2411 THEN
            tanh_f := 1692;
        ELSIF x = 2412 THEN
            tanh_f := 1692;
        ELSIF x = 2413 THEN
            tanh_f := 1692;
        ELSIF x = 2414 THEN
            tanh_f := 1693;
        ELSIF x = 2415 THEN
            tanh_f := 1693;
        ELSIF x = 2416 THEN
            tanh_f := 1693;
        ELSIF x = 2417 THEN
            tanh_f := 1694;
        ELSIF x = 2418 THEN
            tanh_f := 1694;
        ELSIF x = 2419 THEN
            tanh_f := 1694;
        ELSIF x = 2420 THEN
            tanh_f := 1694;
        ELSIF x = 2421 THEN
            tanh_f := 1695;
        ELSIF x = 2422 THEN
            tanh_f := 1695;
        ELSIF x = 2423 THEN
            tanh_f := 1695;
        ELSIF x = 2424 THEN
            tanh_f := 1696;
        ELSIF x = 2425 THEN
            tanh_f := 1696;
        ELSIF x = 2426 THEN
            tanh_f := 1696;
        ELSIF x = 2427 THEN
            tanh_f := 1697;
        ELSIF x = 2428 THEN
            tanh_f := 1697;
        ELSIF x = 2429 THEN
            tanh_f := 1697;
        ELSIF x = 2430 THEN
            tanh_f := 1698;
        ELSIF x = 2431 THEN
            tanh_f := 1698;
        ELSIF x = 2432 THEN
            tanh_f := 1698;
        ELSIF x = 2433 THEN
            tanh_f := 1699;
        ELSIF x = 2434 THEN
            tanh_f := 1699;
        ELSIF x = 2435 THEN
            tanh_f := 1699;
        ELSIF x = 2436 THEN
            tanh_f := 1700;
        ELSIF x = 2437 THEN
            tanh_f := 1700;
        ELSIF x = 2438 THEN
            tanh_f := 1700;
        ELSIF x = 2439 THEN
            tanh_f := 1700;
        ELSIF x = 2440 THEN
            tanh_f := 1701;
        ELSIF x = 2441 THEN
            tanh_f := 1701;
        ELSIF x = 2442 THEN
            tanh_f := 1701;
        ELSIF x = 2443 THEN
            tanh_f := 1702;
        ELSIF x = 2444 THEN
            tanh_f := 1702;
        ELSIF x = 2445 THEN
            tanh_f := 1702;
        ELSIF x = 2446 THEN
            tanh_f := 1703;
        ELSIF x = 2447 THEN
            tanh_f := 1703;
        ELSIF x = 2448 THEN
            tanh_f := 1703;
        ELSIF x = 2449 THEN
            tanh_f := 1704;
        ELSIF x = 2450 THEN
            tanh_f := 1704;
        ELSIF x = 2451 THEN
            tanh_f := 1704;
        ELSIF x = 2452 THEN
            tanh_f := 1705;
        ELSIF x = 2453 THEN
            tanh_f := 1705;
        ELSIF x = 2454 THEN
            tanh_f := 1705;
        ELSIF x = 2455 THEN
            tanh_f := 1705;
        ELSIF x = 2456 THEN
            tanh_f := 1706;
        ELSIF x = 2457 THEN
            tanh_f := 1706;
        ELSIF x = 2458 THEN
            tanh_f := 1706;
        ELSIF x = 2459 THEN
            tanh_f := 1707;
        ELSIF x = 2460 THEN
            tanh_f := 1707;
        ELSIF x = 2461 THEN
            tanh_f := 1707;
        ELSIF x = 2462 THEN
            tanh_f := 1708;
        ELSIF x = 2463 THEN
            tanh_f := 1708;
        ELSIF x = 2464 THEN
            tanh_f := 1708;
        ELSIF x = 2465 THEN
            tanh_f := 1709;
        ELSIF x = 2466 THEN
            tanh_f := 1709;
        ELSIF x = 2467 THEN
            tanh_f := 1709;
        ELSIF x = 2468 THEN
            tanh_f := 1710;
        ELSIF x = 2469 THEN
            tanh_f := 1710;
        ELSIF x = 2470 THEN
            tanh_f := 1710;
        ELSIF x = 2471 THEN
            tanh_f := 1711;
        ELSIF x = 2472 THEN
            tanh_f := 1711;
        ELSIF x = 2473 THEN
            tanh_f := 1711;
        ELSIF x = 2474 THEN
            tanh_f := 1711;
        ELSIF x = 2475 THEN
            tanh_f := 1712;
        ELSIF x = 2476 THEN
            tanh_f := 1712;
        ELSIF x = 2477 THEN
            tanh_f := 1712;
        ELSIF x = 2478 THEN
            tanh_f := 1713;
        ELSIF x = 2479 THEN
            tanh_f := 1713;
        ELSIF x = 2480 THEN
            tanh_f := 1713;
        ELSIF x = 2481 THEN
            tanh_f := 1714;
        ELSIF x = 2482 THEN
            tanh_f := 1714;
        ELSIF x = 2483 THEN
            tanh_f := 1714;
        ELSIF x = 2484 THEN
            tanh_f := 1715;
        ELSIF x = 2485 THEN
            tanh_f := 1715;
        ELSIF x = 2486 THEN
            tanh_f := 1715;
        ELSIF x = 2487 THEN
            tanh_f := 1716;
        ELSIF x = 2488 THEN
            tanh_f := 1716;
        ELSIF x = 2489 THEN
            tanh_f := 1716;
        ELSIF x = 2490 THEN
            tanh_f := 1716;
        ELSIF x = 2491 THEN
            tanh_f := 1717;
        ELSIF x = 2492 THEN
            tanh_f := 1717;
        ELSIF x = 2493 THEN
            tanh_f := 1717;
        ELSIF x = 2494 THEN
            tanh_f := 1718;
        ELSIF x = 2495 THEN
            tanh_f := 1718;
        ELSIF x = 2496 THEN
            tanh_f := 1718;
        ELSIF x = 2497 THEN
            tanh_f := 1719;
        ELSIF x = 2498 THEN
            tanh_f := 1719;
        ELSIF x = 2499 THEN
            tanh_f := 1719;
        ELSIF x = 2500 THEN
            tanh_f := 1720;
        ELSIF x = 2501 THEN
            tanh_f := 1720;
        ELSIF x = 2502 THEN
            tanh_f := 1720;
        ELSIF x = 2503 THEN
            tanh_f := 1721;
        ELSIF x = 2504 THEN
            tanh_f := 1721;
        ELSIF x = 2505 THEN
            tanh_f := 1721;
        ELSIF x = 2506 THEN
            tanh_f := 1722;
        ELSIF x = 2507 THEN
            tanh_f := 1722;
        ELSIF x = 2508 THEN
            tanh_f := 1722;
        ELSIF x = 2509 THEN
            tanh_f := 1722;
        ELSIF x = 2510 THEN
            tanh_f := 1723;
        ELSIF x = 2511 THEN
            tanh_f := 1723;
        ELSIF x = 2512 THEN
            tanh_f := 1723;
        ELSIF x = 2513 THEN
            tanh_f := 1724;
        ELSIF x = 2514 THEN
            tanh_f := 1724;
        ELSIF x = 2515 THEN
            tanh_f := 1724;
        ELSIF x = 2516 THEN
            tanh_f := 1725;
        ELSIF x = 2517 THEN
            tanh_f := 1725;
        ELSIF x = 2518 THEN
            tanh_f := 1725;
        ELSIF x = 2519 THEN
            tanh_f := 1726;
        ELSIF x = 2520 THEN
            tanh_f := 1726;
        ELSIF x = 2521 THEN
            tanh_f := 1726;
        ELSIF x = 2522 THEN
            tanh_f := 1727;
        ELSIF x = 2523 THEN
            tanh_f := 1727;
        ELSIF x = 2524 THEN
            tanh_f := 1727;
        ELSIF x = 2525 THEN
            tanh_f := 1727;
        ELSIF x = 2526 THEN
            tanh_f := 1728;
        ELSIF x = 2527 THEN
            tanh_f := 1728;
        ELSIF x = 2528 THEN
            tanh_f := 1728;
        ELSIF x = 2529 THEN
            tanh_f := 1729;
        ELSIF x = 2530 THEN
            tanh_f := 1729;
        ELSIF x = 2531 THEN
            tanh_f := 1729;
        ELSIF x = 2532 THEN
            tanh_f := 1730;
        ELSIF x = 2533 THEN
            tanh_f := 1730;
        ELSIF x = 2534 THEN
            tanh_f := 1730;
        ELSIF x = 2535 THEN
            tanh_f := 1731;
        ELSIF x = 2536 THEN
            tanh_f := 1731;
        ELSIF x = 2537 THEN
            tanh_f := 1731;
        ELSIF x = 2538 THEN
            tanh_f := 1732;
        ELSIF x = 2539 THEN
            tanh_f := 1732;
        ELSIF x = 2540 THEN
            tanh_f := 1732;
        ELSIF x = 2541 THEN
            tanh_f := 1733;
        ELSIF x = 2542 THEN
            tanh_f := 1733;
        ELSIF x = 2543 THEN
            tanh_f := 1733;
        ELSIF x = 2544 THEN
            tanh_f := 1733;
        ELSIF x = 2545 THEN
            tanh_f := 1734;
        ELSIF x = 2546 THEN
            tanh_f := 1734;
        ELSIF x = 2547 THEN
            tanh_f := 1734;
        ELSIF x = 2548 THEN
            tanh_f := 1735;
        ELSIF x = 2549 THEN
            tanh_f := 1735;
        ELSIF x = 2550 THEN
            tanh_f := 1735;
        ELSIF x = 2551 THEN
            tanh_f := 1736;
        ELSIF x = 2552 THEN
            tanh_f := 1736;
        ELSIF x = 2553 THEN
            tanh_f := 1736;
        ELSIF x = 2554 THEN
            tanh_f := 1737;
        ELSIF x = 2555 THEN
            tanh_f := 1737;
        ELSIF x = 2556 THEN
            tanh_f := 1737;
        ELSIF x = 2557 THEN
            tanh_f := 1738;
        ELSIF x = 2558 THEN
            tanh_f := 1738;
        ELSIF x = 2559 THEN
            tanh_f := 1738;
        ELSIF x = 2560 THEN
            tanh_f := 1739;
        ELSIF x = 2561 THEN
            tanh_f := 1739;
        ELSIF x = 2562 THEN
            tanh_f := 1739;
        ELSIF x = 2563 THEN
            tanh_f := 1739;
        ELSIF x = 2564 THEN
            tanh_f := 1739;
        ELSIF x = 2565 THEN
            tanh_f := 1740;
        ELSIF x = 2566 THEN
            tanh_f := 1740;
        ELSIF x = 2567 THEN
            tanh_f := 1740;
        ELSIF x = 2568 THEN
            tanh_f := 1740;
        ELSIF x = 2569 THEN
            tanh_f := 1741;
        ELSIF x = 2570 THEN
            tanh_f := 1741;
        ELSIF x = 2571 THEN
            tanh_f := 1741;
        ELSIF x = 2572 THEN
            tanh_f := 1741;
        ELSIF x = 2573 THEN
            tanh_f := 1742;
        ELSIF x = 2574 THEN
            tanh_f := 1742;
        ELSIF x = 2575 THEN
            tanh_f := 1742;
        ELSIF x = 2576 THEN
            tanh_f := 1742;
        ELSIF x = 2577 THEN
            tanh_f := 1743;
        ELSIF x = 2578 THEN
            tanh_f := 1743;
        ELSIF x = 2579 THEN
            tanh_f := 1743;
        ELSIF x = 2580 THEN
            tanh_f := 1743;
        ELSIF x = 2581 THEN
            tanh_f := 1744;
        ELSIF x = 2582 THEN
            tanh_f := 1744;
        ELSIF x = 2583 THEN
            tanh_f := 1744;
        ELSIF x = 2584 THEN
            tanh_f := 1744;
        ELSIF x = 2585 THEN
            tanh_f := 1745;
        ELSIF x = 2586 THEN
            tanh_f := 1745;
        ELSIF x = 2587 THEN
            tanh_f := 1745;
        ELSIF x = 2588 THEN
            tanh_f := 1745;
        ELSIF x = 2589 THEN
            tanh_f := 1746;
        ELSIF x = 2590 THEN
            tanh_f := 1746;
        ELSIF x = 2591 THEN
            tanh_f := 1746;
        ELSIF x = 2592 THEN
            tanh_f := 1746;
        ELSIF x = 2593 THEN
            tanh_f := 1747;
        ELSIF x = 2594 THEN
            tanh_f := 1747;
        ELSIF x = 2595 THEN
            tanh_f := 1747;
        ELSIF x = 2596 THEN
            tanh_f := 1747;
        ELSIF x = 2597 THEN
            tanh_f := 1748;
        ELSIF x = 2598 THEN
            tanh_f := 1748;
        ELSIF x = 2599 THEN
            tanh_f := 1748;
        ELSIF x = 2600 THEN
            tanh_f := 1748;
        ELSIF x = 2601 THEN
            tanh_f := 1749;
        ELSIF x = 2602 THEN
            tanh_f := 1749;
        ELSIF x = 2603 THEN
            tanh_f := 1749;
        ELSIF x = 2604 THEN
            tanh_f := 1749;
        ELSIF x = 2605 THEN
            tanh_f := 1750;
        ELSIF x = 2606 THEN
            tanh_f := 1750;
        ELSIF x = 2607 THEN
            tanh_f := 1750;
        ELSIF x = 2608 THEN
            tanh_f := 1750;
        ELSIF x = 2609 THEN
            tanh_f := 1751;
        ELSIF x = 2610 THEN
            tanh_f := 1751;
        ELSIF x = 2611 THEN
            tanh_f := 1751;
        ELSIF x = 2612 THEN
            tanh_f := 1751;
        ELSIF x = 2613 THEN
            tanh_f := 1752;
        ELSIF x = 2614 THEN
            tanh_f := 1752;
        ELSIF x = 2615 THEN
            tanh_f := 1752;
        ELSIF x = 2616 THEN
            tanh_f := 1752;
        ELSIF x = 2617 THEN
            tanh_f := 1753;
        ELSIF x = 2618 THEN
            tanh_f := 1753;
        ELSIF x = 2619 THEN
            tanh_f := 1753;
        ELSIF x = 2620 THEN
            tanh_f := 1753;
        ELSIF x = 2621 THEN
            tanh_f := 1754;
        ELSIF x = 2622 THEN
            tanh_f := 1754;
        ELSIF x = 2623 THEN
            tanh_f := 1754;
        ELSIF x = 2624 THEN
            tanh_f := 1754;
        ELSIF x = 2625 THEN
            tanh_f := 1755;
        ELSIF x = 2626 THEN
            tanh_f := 1755;
        ELSIF x = 2627 THEN
            tanh_f := 1755;
        ELSIF x = 2628 THEN
            tanh_f := 1755;
        ELSIF x = 2629 THEN
            tanh_f := 1756;
        ELSIF x = 2630 THEN
            tanh_f := 1756;
        ELSIF x = 2631 THEN
            tanh_f := 1756;
        ELSIF x = 2632 THEN
            tanh_f := 1756;
        ELSIF x = 2633 THEN
            tanh_f := 1757;
        ELSIF x = 2634 THEN
            tanh_f := 1757;
        ELSIF x = 2635 THEN
            tanh_f := 1757;
        ELSIF x = 2636 THEN
            tanh_f := 1757;
        ELSIF x = 2637 THEN
            tanh_f := 1758;
        ELSIF x = 2638 THEN
            tanh_f := 1758;
        ELSIF x = 2639 THEN
            tanh_f := 1758;
        ELSIF x = 2640 THEN
            tanh_f := 1758;
        ELSIF x = 2641 THEN
            tanh_f := 1759;
        ELSIF x = 2642 THEN
            tanh_f := 1759;
        ELSIF x = 2643 THEN
            tanh_f := 1759;
        ELSIF x = 2644 THEN
            tanh_f := 1759;
        ELSIF x = 2645 THEN
            tanh_f := 1760;
        ELSIF x = 2646 THEN
            tanh_f := 1760;
        ELSIF x = 2647 THEN
            tanh_f := 1760;
        ELSIF x = 2648 THEN
            tanh_f := 1760;
        ELSIF x = 2649 THEN
            tanh_f := 1761;
        ELSIF x = 2650 THEN
            tanh_f := 1761;
        ELSIF x = 2651 THEN
            tanh_f := 1761;
        ELSIF x = 2652 THEN
            tanh_f := 1761;
        ELSIF x = 2653 THEN
            tanh_f := 1762;
        ELSIF x = 2654 THEN
            tanh_f := 1762;
        ELSIF x = 2655 THEN
            tanh_f := 1762;
        ELSIF x = 2656 THEN
            tanh_f := 1762;
        ELSIF x = 2657 THEN
            tanh_f := 1763;
        ELSIF x = 2658 THEN
            tanh_f := 1763;
        ELSIF x = 2659 THEN
            tanh_f := 1763;
        ELSIF x = 2660 THEN
            tanh_f := 1763;
        ELSIF x = 2661 THEN
            tanh_f := 1764;
        ELSIF x = 2662 THEN
            tanh_f := 1764;
        ELSIF x = 2663 THEN
            tanh_f := 1764;
        ELSIF x = 2664 THEN
            tanh_f := 1764;
        ELSIF x = 2665 THEN
            tanh_f := 1765;
        ELSIF x = 2666 THEN
            tanh_f := 1765;
        ELSIF x = 2667 THEN
            tanh_f := 1765;
        ELSIF x = 2668 THEN
            tanh_f := 1765;
        ELSIF x = 2669 THEN
            tanh_f := 1766;
        ELSIF x = 2670 THEN
            tanh_f := 1766;
        ELSIF x = 2671 THEN
            tanh_f := 1766;
        ELSIF x = 2672 THEN
            tanh_f := 1766;
        ELSIF x = 2673 THEN
            tanh_f := 1767;
        ELSIF x = 2674 THEN
            tanh_f := 1767;
        ELSIF x = 2675 THEN
            tanh_f := 1767;
        ELSIF x = 2676 THEN
            tanh_f := 1767;
        ELSIF x = 2677 THEN
            tanh_f := 1768;
        ELSIF x = 2678 THEN
            tanh_f := 1768;
        ELSIF x = 2679 THEN
            tanh_f := 1768;
        ELSIF x = 2680 THEN
            tanh_f := 1768;
        ELSIF x = 2681 THEN
            tanh_f := 1769;
        ELSIF x = 2682 THEN
            tanh_f := 1769;
        ELSIF x = 2683 THEN
            tanh_f := 1769;
        ELSIF x = 2684 THEN
            tanh_f := 1769;
        ELSIF x = 2685 THEN
            tanh_f := 1770;
        ELSIF x = 2686 THEN
            tanh_f := 1770;
        ELSIF x = 2687 THEN
            tanh_f := 1770;
        ELSIF x = 2688 THEN
            tanh_f := 1770;
        ELSIF x = 2689 THEN
            tanh_f := 1770;
        ELSIF x = 2690 THEN
            tanh_f := 1771;
        ELSIF x = 2691 THEN
            tanh_f := 1771;
        ELSIF x = 2692 THEN
            tanh_f := 1771;
        ELSIF x = 2693 THEN
            tanh_f := 1771;
        ELSIF x = 2694 THEN
            tanh_f := 1772;
        ELSIF x = 2695 THEN
            tanh_f := 1772;
        ELSIF x = 2696 THEN
            tanh_f := 1772;
        ELSIF x = 2697 THEN
            tanh_f := 1772;
        ELSIF x = 2698 THEN
            tanh_f := 1773;
        ELSIF x = 2699 THEN
            tanh_f := 1773;
        ELSIF x = 2700 THEN
            tanh_f := 1773;
        ELSIF x = 2701 THEN
            tanh_f := 1773;
        ELSIF x = 2702 THEN
            tanh_f := 1774;
        ELSIF x = 2703 THEN
            tanh_f := 1774;
        ELSIF x = 2704 THEN
            tanh_f := 1774;
        ELSIF x = 2705 THEN
            tanh_f := 1774;
        ELSIF x = 2706 THEN
            tanh_f := 1775;
        ELSIF x = 2707 THEN
            tanh_f := 1775;
        ELSIF x = 2708 THEN
            tanh_f := 1775;
        ELSIF x = 2709 THEN
            tanh_f := 1775;
        ELSIF x = 2710 THEN
            tanh_f := 1776;
        ELSIF x = 2711 THEN
            tanh_f := 1776;
        ELSIF x = 2712 THEN
            tanh_f := 1776;
        ELSIF x = 2713 THEN
            tanh_f := 1776;
        ELSIF x = 2714 THEN
            tanh_f := 1777;
        ELSIF x = 2715 THEN
            tanh_f := 1777;
        ELSIF x = 2716 THEN
            tanh_f := 1777;
        ELSIF x = 2717 THEN
            tanh_f := 1777;
        ELSIF x = 2718 THEN
            tanh_f := 1778;
        ELSIF x = 2719 THEN
            tanh_f := 1778;
        ELSIF x = 2720 THEN
            tanh_f := 1778;
        ELSIF x = 2721 THEN
            tanh_f := 1778;
        ELSIF x = 2722 THEN
            tanh_f := 1779;
        ELSIF x = 2723 THEN
            tanh_f := 1779;
        ELSIF x = 2724 THEN
            tanh_f := 1779;
        ELSIF x = 2725 THEN
            tanh_f := 1779;
        ELSIF x = 2726 THEN
            tanh_f := 1780;
        ELSIF x = 2727 THEN
            tanh_f := 1780;
        ELSIF x = 2728 THEN
            tanh_f := 1780;
        ELSIF x = 2729 THEN
            tanh_f := 1780;
        ELSIF x = 2730 THEN
            tanh_f := 1781;
        ELSIF x = 2731 THEN
            tanh_f := 1781;
        ELSIF x = 2732 THEN
            tanh_f := 1781;
        ELSIF x = 2733 THEN
            tanh_f := 1781;
        ELSIF x = 2734 THEN
            tanh_f := 1782;
        ELSIF x = 2735 THEN
            tanh_f := 1782;
        ELSIF x = 2736 THEN
            tanh_f := 1782;
        ELSIF x = 2737 THEN
            tanh_f := 1782;
        ELSIF x = 2738 THEN
            tanh_f := 1783;
        ELSIF x = 2739 THEN
            tanh_f := 1783;
        ELSIF x = 2740 THEN
            tanh_f := 1783;
        ELSIF x = 2741 THEN
            tanh_f := 1783;
        ELSIF x = 2742 THEN
            tanh_f := 1784;
        ELSIF x = 2743 THEN
            tanh_f := 1784;
        ELSIF x = 2744 THEN
            tanh_f := 1784;
        ELSIF x = 2745 THEN
            tanh_f := 1784;
        ELSIF x = 2746 THEN
            tanh_f := 1785;
        ELSIF x = 2747 THEN
            tanh_f := 1785;
        ELSIF x = 2748 THEN
            tanh_f := 1785;
        ELSIF x = 2749 THEN
            tanh_f := 1785;
        ELSIF x = 2750 THEN
            tanh_f := 1786;
        ELSIF x = 2751 THEN
            tanh_f := 1786;
        ELSIF x = 2752 THEN
            tanh_f := 1786;
        ELSIF x = 2753 THEN
            tanh_f := 1786;
        ELSIF x = 2754 THEN
            tanh_f := 1787;
        ELSIF x = 2755 THEN
            tanh_f := 1787;
        ELSIF x = 2756 THEN
            tanh_f := 1787;
        ELSIF x = 2757 THEN
            tanh_f := 1787;
        ELSIF x = 2758 THEN
            tanh_f := 1788;
        ELSIF x = 2759 THEN
            tanh_f := 1788;
        ELSIF x = 2760 THEN
            tanh_f := 1788;
        ELSIF x = 2761 THEN
            tanh_f := 1788;
        ELSIF x = 2762 THEN
            tanh_f := 1789;
        ELSIF x = 2763 THEN
            tanh_f := 1789;
        ELSIF x = 2764 THEN
            tanh_f := 1789;
        ELSIF x = 2765 THEN
            tanh_f := 1789;
        ELSIF x = 2766 THEN
            tanh_f := 1790;
        ELSIF x = 2767 THEN
            tanh_f := 1790;
        ELSIF x = 2768 THEN
            tanh_f := 1790;
        ELSIF x = 2769 THEN
            tanh_f := 1790;
        ELSIF x = 2770 THEN
            tanh_f := 1791;
        ELSIF x = 2771 THEN
            tanh_f := 1791;
        ELSIF x = 2772 THEN
            tanh_f := 1791;
        ELSIF x = 2773 THEN
            tanh_f := 1791;
        ELSIF x = 2774 THEN
            tanh_f := 1792;
        ELSIF x = 2775 THEN
            tanh_f := 1792;
        ELSIF x = 2776 THEN
            tanh_f := 1792;
        ELSIF x = 2777 THEN
            tanh_f := 1792;
        ELSIF x = 2778 THEN
            tanh_f := 1793;
        ELSIF x = 2779 THEN
            tanh_f := 1793;
        ELSIF x = 2780 THEN
            tanh_f := 1793;
        ELSIF x = 2781 THEN
            tanh_f := 1793;
        ELSIF x = 2782 THEN
            tanh_f := 1794;
        ELSIF x = 2783 THEN
            tanh_f := 1794;
        ELSIF x = 2784 THEN
            tanh_f := 1794;
        ELSIF x = 2785 THEN
            tanh_f := 1794;
        ELSIF x = 2786 THEN
            tanh_f := 1795;
        ELSIF x = 2787 THEN
            tanh_f := 1795;
        ELSIF x = 2788 THEN
            tanh_f := 1795;
        ELSIF x = 2789 THEN
            tanh_f := 1795;
        ELSIF x = 2790 THEN
            tanh_f := 1796;
        ELSIF x = 2791 THEN
            tanh_f := 1796;
        ELSIF x = 2792 THEN
            tanh_f := 1796;
        ELSIF x = 2793 THEN
            tanh_f := 1796;
        ELSIF x = 2794 THEN
            tanh_f := 1797;
        ELSIF x = 2795 THEN
            tanh_f := 1797;
        ELSIF x = 2796 THEN
            tanh_f := 1797;
        ELSIF x = 2797 THEN
            tanh_f := 1797;
        ELSIF x = 2798 THEN
            tanh_f := 1798;
        ELSIF x = 2799 THEN
            tanh_f := 1798;
        ELSIF x = 2800 THEN
            tanh_f := 1798;
        ELSIF x = 2801 THEN
            tanh_f := 1798;
        ELSIF x = 2802 THEN
            tanh_f := 1799;
        ELSIF x = 2803 THEN
            tanh_f := 1799;
        ELSIF x = 2804 THEN
            tanh_f := 1799;
        ELSIF x = 2805 THEN
            tanh_f := 1799;
        ELSIF x = 2806 THEN
            tanh_f := 1800;
        ELSIF x = 2807 THEN
            tanh_f := 1800;
        ELSIF x = 2808 THEN
            tanh_f := 1800;
        ELSIF x = 2809 THEN
            tanh_f := 1800;
        ELSIF x = 2810 THEN
            tanh_f := 1801;
        ELSIF x = 2811 THEN
            tanh_f := 1801;
        ELSIF x = 2812 THEN
            tanh_f := 1801;
        ELSIF x = 2813 THEN
            tanh_f := 1801;
        ELSIF x = 2814 THEN
            tanh_f := 1802;
        ELSIF x = 2815 THEN
            tanh_f := 1802;
        ELSIF x = 2816 THEN
            tanh_f := 1803;
        ELSIF x = 2817 THEN
            tanh_f := 1803;
        ELSIF x = 2818 THEN
            tanh_f := 1803;
        ELSIF x = 2819 THEN
            tanh_f := 1803;
        ELSIF x = 2820 THEN
            tanh_f := 1803;
        ELSIF x = 2821 THEN
            tanh_f := 1803;
        ELSIF x = 2822 THEN
            tanh_f := 1804;
        ELSIF x = 2823 THEN
            tanh_f := 1804;
        ELSIF x = 2824 THEN
            tanh_f := 1804;
        ELSIF x = 2825 THEN
            tanh_f := 1804;
        ELSIF x = 2826 THEN
            tanh_f := 1804;
        ELSIF x = 2827 THEN
            tanh_f := 1805;
        ELSIF x = 2828 THEN
            tanh_f := 1805;
        ELSIF x = 2829 THEN
            tanh_f := 1805;
        ELSIF x = 2830 THEN
            tanh_f := 1805;
        ELSIF x = 2831 THEN
            tanh_f := 1805;
        ELSIF x = 2832 THEN
            tanh_f := 1806;
        ELSIF x = 2833 THEN
            tanh_f := 1806;
        ELSIF x = 2834 THEN
            tanh_f := 1806;
        ELSIF x = 2835 THEN
            tanh_f := 1806;
        ELSIF x = 2836 THEN
            tanh_f := 1806;
        ELSIF x = 2837 THEN
            tanh_f := 1807;
        ELSIF x = 2838 THEN
            tanh_f := 1807;
        ELSIF x = 2839 THEN
            tanh_f := 1807;
        ELSIF x = 2840 THEN
            tanh_f := 1807;
        ELSIF x = 2841 THEN
            tanh_f := 1807;
        ELSIF x = 2842 THEN
            tanh_f := 1808;
        ELSIF x = 2843 THEN
            tanh_f := 1808;
        ELSIF x = 2844 THEN
            tanh_f := 1808;
        ELSIF x = 2845 THEN
            tanh_f := 1808;
        ELSIF x = 2846 THEN
            tanh_f := 1808;
        ELSIF x = 2847 THEN
            tanh_f := 1809;
        ELSIF x = 2848 THEN
            tanh_f := 1809;
        ELSIF x = 2849 THEN
            tanh_f := 1809;
        ELSIF x = 2850 THEN
            tanh_f := 1809;
        ELSIF x = 2851 THEN
            tanh_f := 1809;
        ELSIF x = 2852 THEN
            tanh_f := 1810;
        ELSIF x = 2853 THEN
            tanh_f := 1810;
        ELSIF x = 2854 THEN
            tanh_f := 1810;
        ELSIF x = 2855 THEN
            tanh_f := 1810;
        ELSIF x = 2856 THEN
            tanh_f := 1810;
        ELSIF x = 2857 THEN
            tanh_f := 1811;
        ELSIF x = 2858 THEN
            tanh_f := 1811;
        ELSIF x = 2859 THEN
            tanh_f := 1811;
        ELSIF x = 2860 THEN
            tanh_f := 1811;
        ELSIF x = 2861 THEN
            tanh_f := 1811;
        ELSIF x = 2862 THEN
            tanh_f := 1812;
        ELSIF x = 2863 THEN
            tanh_f := 1812;
        ELSIF x = 2864 THEN
            tanh_f := 1812;
        ELSIF x = 2865 THEN
            tanh_f := 1812;
        ELSIF x = 2866 THEN
            tanh_f := 1812;
        ELSIF x = 2867 THEN
            tanh_f := 1813;
        ELSIF x = 2868 THEN
            tanh_f := 1813;
        ELSIF x = 2869 THEN
            tanh_f := 1813;
        ELSIF x = 2870 THEN
            tanh_f := 1813;
        ELSIF x = 2871 THEN
            tanh_f := 1813;
        ELSIF x = 2872 THEN
            tanh_f := 1814;
        ELSIF x = 2873 THEN
            tanh_f := 1814;
        ELSIF x = 2874 THEN
            tanh_f := 1814;
        ELSIF x = 2875 THEN
            tanh_f := 1814;
        ELSIF x = 2876 THEN
            tanh_f := 1814;
        ELSIF x = 2877 THEN
            tanh_f := 1815;
        ELSIF x = 2878 THEN
            tanh_f := 1815;
        ELSIF x = 2879 THEN
            tanh_f := 1815;
        ELSIF x = 2880 THEN
            tanh_f := 1815;
        ELSIF x = 2881 THEN
            tanh_f := 1815;
        ELSIF x = 2882 THEN
            tanh_f := 1816;
        ELSIF x = 2883 THEN
            tanh_f := 1816;
        ELSIF x = 2884 THEN
            tanh_f := 1816;
        ELSIF x = 2885 THEN
            tanh_f := 1816;
        ELSIF x = 2886 THEN
            tanh_f := 1816;
        ELSIF x = 2887 THEN
            tanh_f := 1817;
        ELSIF x = 2888 THEN
            tanh_f := 1817;
        ELSIF x = 2889 THEN
            tanh_f := 1817;
        ELSIF x = 2890 THEN
            tanh_f := 1817;
        ELSIF x = 2891 THEN
            tanh_f := 1817;
        ELSIF x = 2892 THEN
            tanh_f := 1818;
        ELSIF x = 2893 THEN
            tanh_f := 1818;
        ELSIF x = 2894 THEN
            tanh_f := 1818;
        ELSIF x = 2895 THEN
            tanh_f := 1818;
        ELSIF x = 2896 THEN
            tanh_f := 1818;
        ELSIF x = 2897 THEN
            tanh_f := 1819;
        ELSIF x = 2898 THEN
            tanh_f := 1819;
        ELSIF x = 2899 THEN
            tanh_f := 1819;
        ELSIF x = 2900 THEN
            tanh_f := 1819;
        ELSIF x = 2901 THEN
            tanh_f := 1819;
        ELSIF x = 2902 THEN
            tanh_f := 1820;
        ELSIF x = 2903 THEN
            tanh_f := 1820;
        ELSIF x = 2904 THEN
            tanh_f := 1820;
        ELSIF x = 2905 THEN
            tanh_f := 1820;
        ELSIF x = 2906 THEN
            tanh_f := 1820;
        ELSIF x = 2907 THEN
            tanh_f := 1821;
        ELSIF x = 2908 THEN
            tanh_f := 1821;
        ELSIF x = 2909 THEN
            tanh_f := 1821;
        ELSIF x = 2910 THEN
            tanh_f := 1821;
        ELSIF x = 2911 THEN
            tanh_f := 1821;
        ELSIF x = 2912 THEN
            tanh_f := 1822;
        ELSIF x = 2913 THEN
            tanh_f := 1822;
        ELSIF x = 2914 THEN
            tanh_f := 1822;
        ELSIF x = 2915 THEN
            tanh_f := 1822;
        ELSIF x = 2916 THEN
            tanh_f := 1822;
        ELSIF x = 2917 THEN
            tanh_f := 1823;
        ELSIF x = 2918 THEN
            tanh_f := 1823;
        ELSIF x = 2919 THEN
            tanh_f := 1823;
        ELSIF x = 2920 THEN
            tanh_f := 1823;
        ELSIF x = 2921 THEN
            tanh_f := 1823;
        ELSIF x = 2922 THEN
            tanh_f := 1824;
        ELSIF x = 2923 THEN
            tanh_f := 1824;
        ELSIF x = 2924 THEN
            tanh_f := 1824;
        ELSIF x = 2925 THEN
            tanh_f := 1824;
        ELSIF x = 2926 THEN
            tanh_f := 1824;
        ELSIF x = 2927 THEN
            tanh_f := 1825;
        ELSIF x = 2928 THEN
            tanh_f := 1825;
        ELSIF x = 2929 THEN
            tanh_f := 1825;
        ELSIF x = 2930 THEN
            tanh_f := 1825;
        ELSIF x = 2931 THEN
            tanh_f := 1825;
        ELSIF x = 2932 THEN
            tanh_f := 1826;
        ELSIF x = 2933 THEN
            tanh_f := 1826;
        ELSIF x = 2934 THEN
            tanh_f := 1826;
        ELSIF x = 2935 THEN
            tanh_f := 1826;
        ELSIF x = 2936 THEN
            tanh_f := 1826;
        ELSIF x = 2937 THEN
            tanh_f := 1827;
        ELSIF x = 2938 THEN
            tanh_f := 1827;
        ELSIF x = 2939 THEN
            tanh_f := 1827;
        ELSIF x = 2940 THEN
            tanh_f := 1827;
        ELSIF x = 2941 THEN
            tanh_f := 1827;
        ELSIF x = 2942 THEN
            tanh_f := 1828;
        ELSIF x = 2943 THEN
            tanh_f := 1828;
        ELSIF x = 2944 THEN
            tanh_f := 1828;
        ELSIF x = 2945 THEN
            tanh_f := 1828;
        ELSIF x = 2946 THEN
            tanh_f := 1828;
        ELSIF x = 2947 THEN
            tanh_f := 1829;
        ELSIF x = 2948 THEN
            tanh_f := 1829;
        ELSIF x = 2949 THEN
            tanh_f := 1829;
        ELSIF x = 2950 THEN
            tanh_f := 1829;
        ELSIF x = 2951 THEN
            tanh_f := 1829;
        ELSIF x = 2952 THEN
            tanh_f := 1830;
        ELSIF x = 2953 THEN
            tanh_f := 1830;
        ELSIF x = 2954 THEN
            tanh_f := 1830;
        ELSIF x = 2955 THEN
            tanh_f := 1830;
        ELSIF x = 2956 THEN
            tanh_f := 1830;
        ELSIF x = 2957 THEN
            tanh_f := 1831;
        ELSIF x = 2958 THEN
            tanh_f := 1831;
        ELSIF x = 2959 THEN
            tanh_f := 1831;
        ELSIF x = 2960 THEN
            tanh_f := 1831;
        ELSIF x = 2961 THEN
            tanh_f := 1831;
        ELSIF x = 2962 THEN
            tanh_f := 1832;
        ELSIF x = 2963 THEN
            tanh_f := 1832;
        ELSIF x = 2964 THEN
            tanh_f := 1832;
        ELSIF x = 2965 THEN
            tanh_f := 1832;
        ELSIF x = 2966 THEN
            tanh_f := 1832;
        ELSIF x = 2967 THEN
            tanh_f := 1833;
        ELSIF x = 2968 THEN
            tanh_f := 1833;
        ELSIF x = 2969 THEN
            tanh_f := 1833;
        ELSIF x = 2970 THEN
            tanh_f := 1833;
        ELSIF x = 2971 THEN
            tanh_f := 1833;
        ELSIF x = 2972 THEN
            tanh_f := 1834;
        ELSIF x = 2973 THEN
            tanh_f := 1834;
        ELSIF x = 2974 THEN
            tanh_f := 1834;
        ELSIF x = 2975 THEN
            tanh_f := 1834;
        ELSIF x = 2976 THEN
            tanh_f := 1834;
        ELSIF x = 2977 THEN
            tanh_f := 1835;
        ELSIF x = 2978 THEN
            tanh_f := 1835;
        ELSIF x = 2979 THEN
            tanh_f := 1835;
        ELSIF x = 2980 THEN
            tanh_f := 1835;
        ELSIF x = 2981 THEN
            tanh_f := 1835;
        ELSIF x = 2982 THEN
            tanh_f := 1836;
        ELSIF x = 2983 THEN
            tanh_f := 1836;
        ELSIF x = 2984 THEN
            tanh_f := 1836;
        ELSIF x = 2985 THEN
            tanh_f := 1836;
        ELSIF x = 2986 THEN
            tanh_f := 1836;
        ELSIF x = 2987 THEN
            tanh_f := 1837;
        ELSIF x = 2988 THEN
            tanh_f := 1837;
        ELSIF x = 2989 THEN
            tanh_f := 1837;
        ELSIF x = 2990 THEN
            tanh_f := 1837;
        ELSIF x = 2991 THEN
            tanh_f := 1837;
        ELSIF x = 2992 THEN
            tanh_f := 1838;
        ELSIF x = 2993 THEN
            tanh_f := 1838;
        ELSIF x = 2994 THEN
            tanh_f := 1838;
        ELSIF x = 2995 THEN
            tanh_f := 1838;
        ELSIF x = 2996 THEN
            tanh_f := 1838;
        ELSIF x = 2997 THEN
            tanh_f := 1839;
        ELSIF x = 2998 THEN
            tanh_f := 1839;
        ELSIF x = 2999 THEN
            tanh_f := 1839;
        ELSIF x = 3000 THEN
            tanh_f := 1839;
        ELSIF x = 3001 THEN
            tanh_f := 1839;
        ELSIF x = 3002 THEN
            tanh_f := 1840;
        ELSIF x = 3003 THEN
            tanh_f := 1840;
        ELSIF x = 3004 THEN
            tanh_f := 1840;
        ELSIF x = 3005 THEN
            tanh_f := 1840;
        ELSIF x = 3006 THEN
            tanh_f := 1840;
        ELSIF x = 3007 THEN
            tanh_f := 1841;
        ELSIF x = 3008 THEN
            tanh_f := 1841;
        ELSIF x = 3009 THEN
            tanh_f := 1841;
        ELSIF x = 3010 THEN
            tanh_f := 1841;
        ELSIF x = 3011 THEN
            tanh_f := 1841;
        ELSIF x = 3012 THEN
            tanh_f := 1842;
        ELSIF x = 3013 THEN
            tanh_f := 1842;
        ELSIF x = 3014 THEN
            tanh_f := 1842;
        ELSIF x = 3015 THEN
            tanh_f := 1842;
        ELSIF x = 3016 THEN
            tanh_f := 1842;
        ELSIF x = 3017 THEN
            tanh_f := 1843;
        ELSIF x = 3018 THEN
            tanh_f := 1843;
        ELSIF x = 3019 THEN
            tanh_f := 1843;
        ELSIF x = 3020 THEN
            tanh_f := 1843;
        ELSIF x = 3021 THEN
            tanh_f := 1843;
        ELSIF x = 3022 THEN
            tanh_f := 1844;
        ELSIF x = 3023 THEN
            tanh_f := 1844;
        ELSIF x = 3024 THEN
            tanh_f := 1844;
        ELSIF x = 3025 THEN
            tanh_f := 1844;
        ELSIF x = 3026 THEN
            tanh_f := 1844;
        ELSIF x = 3027 THEN
            tanh_f := 1845;
        ELSIF x = 3028 THEN
            tanh_f := 1845;
        ELSIF x = 3029 THEN
            tanh_f := 1845;
        ELSIF x = 3030 THEN
            tanh_f := 1845;
        ELSIF x = 3031 THEN
            tanh_f := 1845;
        ELSIF x = 3032 THEN
            tanh_f := 1846;
        ELSIF x = 3033 THEN
            tanh_f := 1846;
        ELSIF x = 3034 THEN
            tanh_f := 1846;
        ELSIF x = 3035 THEN
            tanh_f := 1846;
        ELSIF x = 3036 THEN
            tanh_f := 1846;
        ELSIF x = 3037 THEN
            tanh_f := 1847;
        ELSIF x = 3038 THEN
            tanh_f := 1847;
        ELSIF x = 3039 THEN
            tanh_f := 1847;
        ELSIF x = 3040 THEN
            tanh_f := 1847;
        ELSIF x = 3041 THEN
            tanh_f := 1847;
        ELSIF x = 3042 THEN
            tanh_f := 1848;
        ELSIF x = 3043 THEN
            tanh_f := 1848;
        ELSIF x = 3044 THEN
            tanh_f := 1848;
        ELSIF x = 3045 THEN
            tanh_f := 1848;
        ELSIF x = 3046 THEN
            tanh_f := 1848;
        ELSIF x = 3047 THEN
            tanh_f := 1849;
        ELSIF x = 3048 THEN
            tanh_f := 1849;
        ELSIF x = 3049 THEN
            tanh_f := 1849;
        ELSIF x = 3050 THEN
            tanh_f := 1849;
        ELSIF x = 3051 THEN
            tanh_f := 1849;
        ELSIF x = 3052 THEN
            tanh_f := 1850;
        ELSIF x = 3053 THEN
            tanh_f := 1850;
        ELSIF x = 3054 THEN
            tanh_f := 1850;
        ELSIF x = 3055 THEN
            tanh_f := 1850;
        ELSIF x = 3056 THEN
            tanh_f := 1850;
        ELSIF x = 3057 THEN
            tanh_f := 1851;
        ELSIF x = 3058 THEN
            tanh_f := 1851;
        ELSIF x = 3059 THEN
            tanh_f := 1851;
        ELSIF x = 3060 THEN
            tanh_f := 1851;
        ELSIF x = 3061 THEN
            tanh_f := 1851;
        ELSIF x = 3062 THEN
            tanh_f := 1852;
        ELSIF x = 3063 THEN
            tanh_f := 1852;
        ELSIF x = 3064 THEN
            tanh_f := 1852;
        ELSIF x = 3065 THEN
            tanh_f := 1852;
        ELSIF x = 3066 THEN
            tanh_f := 1852;
        ELSIF x = 3067 THEN
            tanh_f := 1853;
        ELSIF x = 3068 THEN
            tanh_f := 1853;
        ELSIF x = 3069 THEN
            tanh_f := 1853;
        ELSIF x = 3070 THEN
            tanh_f := 1853;
        ELSIF x = 3071 THEN
            tanh_f := 1853;
        ELSIF x = 3072 THEN
            tanh_f := 1854;
        ELSIF x = 3073 THEN
            tanh_f := 1854;
        ELSIF x = 3074 THEN
            tanh_f := 1854;
        ELSIF x = 3075 THEN
            tanh_f := 1854;
        ELSIF x = 3076 THEN
            tanh_f := 1854;
        ELSIF x = 3077 THEN
            tanh_f := 1854;
        ELSIF x = 3078 THEN
            tanh_f := 1854;
        ELSIF x = 3079 THEN
            tanh_f := 1855;
        ELSIF x = 3080 THEN
            tanh_f := 1855;
        ELSIF x = 3081 THEN
            tanh_f := 1855;
        ELSIF x = 3082 THEN
            tanh_f := 1855;
        ELSIF x = 3083 THEN
            tanh_f := 1855;
        ELSIF x = 3084 THEN
            tanh_f := 1855;
        ELSIF x = 3085 THEN
            tanh_f := 1856;
        ELSIF x = 3086 THEN
            tanh_f := 1856;
        ELSIF x = 3087 THEN
            tanh_f := 1856;
        ELSIF x = 3088 THEN
            tanh_f := 1856;
        ELSIF x = 3089 THEN
            tanh_f := 1856;
        ELSIF x = 3090 THEN
            tanh_f := 1856;
        ELSIF x = 3091 THEN
            tanh_f := 1857;
        ELSIF x = 3092 THEN
            tanh_f := 1857;
        ELSIF x = 3093 THEN
            tanh_f := 1857;
        ELSIF x = 3094 THEN
            tanh_f := 1857;
        ELSIF x = 3095 THEN
            tanh_f := 1857;
        ELSIF x = 3096 THEN
            tanh_f := 1857;
        ELSIF x = 3097 THEN
            tanh_f := 1858;
        ELSIF x = 3098 THEN
            tanh_f := 1858;
        ELSIF x = 3099 THEN
            tanh_f := 1858;
        ELSIF x = 3100 THEN
            tanh_f := 1858;
        ELSIF x = 3101 THEN
            tanh_f := 1858;
        ELSIF x = 3102 THEN
            tanh_f := 1858;
        ELSIF x = 3103 THEN
            tanh_f := 1859;
        ELSIF x = 3104 THEN
            tanh_f := 1859;
        ELSIF x = 3105 THEN
            tanh_f := 1859;
        ELSIF x = 3106 THEN
            tanh_f := 1859;
        ELSIF x = 3107 THEN
            tanh_f := 1859;
        ELSIF x = 3108 THEN
            tanh_f := 1859;
        ELSIF x = 3109 THEN
            tanh_f := 1860;
        ELSIF x = 3110 THEN
            tanh_f := 1860;
        ELSIF x = 3111 THEN
            tanh_f := 1860;
        ELSIF x = 3112 THEN
            tanh_f := 1860;
        ELSIF x = 3113 THEN
            tanh_f := 1860;
        ELSIF x = 3114 THEN
            tanh_f := 1860;
        ELSIF x = 3115 THEN
            tanh_f := 1861;
        ELSIF x = 3116 THEN
            tanh_f := 1861;
        ELSIF x = 3117 THEN
            tanh_f := 1861;
        ELSIF x = 3118 THEN
            tanh_f := 1861;
        ELSIF x = 3119 THEN
            tanh_f := 1861;
        ELSIF x = 3120 THEN
            tanh_f := 1861;
        ELSIF x = 3121 THEN
            tanh_f := 1862;
        ELSIF x = 3122 THEN
            tanh_f := 1862;
        ELSIF x = 3123 THEN
            tanh_f := 1862;
        ELSIF x = 3124 THEN
            tanh_f := 1862;
        ELSIF x = 3125 THEN
            tanh_f := 1862;
        ELSIF x = 3126 THEN
            tanh_f := 1862;
        ELSIF x = 3127 THEN
            tanh_f := 1863;
        ELSIF x = 3128 THEN
            tanh_f := 1863;
        ELSIF x = 3129 THEN
            tanh_f := 1863;
        ELSIF x = 3130 THEN
            tanh_f := 1863;
        ELSIF x = 3131 THEN
            tanh_f := 1863;
        ELSIF x = 3132 THEN
            tanh_f := 1863;
        ELSIF x = 3133 THEN
            tanh_f := 1864;
        ELSIF x = 3134 THEN
            tanh_f := 1864;
        ELSIF x = 3135 THEN
            tanh_f := 1864;
        ELSIF x = 3136 THEN
            tanh_f := 1864;
        ELSIF x = 3137 THEN
            tanh_f := 1864;
        ELSIF x = 3138 THEN
            tanh_f := 1864;
        ELSIF x = 3139 THEN
            tanh_f := 1864;
        ELSIF x = 3140 THEN
            tanh_f := 1865;
        ELSIF x = 3141 THEN
            tanh_f := 1865;
        ELSIF x = 3142 THEN
            tanh_f := 1865;
        ELSIF x = 3143 THEN
            tanh_f := 1865;
        ELSIF x = 3144 THEN
            tanh_f := 1865;
        ELSIF x = 3145 THEN
            tanh_f := 1865;
        ELSIF x = 3146 THEN
            tanh_f := 1866;
        ELSIF x = 3147 THEN
            tanh_f := 1866;
        ELSIF x = 3148 THEN
            tanh_f := 1866;
        ELSIF x = 3149 THEN
            tanh_f := 1866;
        ELSIF x = 3150 THEN
            tanh_f := 1866;
        ELSIF x = 3151 THEN
            tanh_f := 1866;
        ELSIF x = 3152 THEN
            tanh_f := 1867;
        ELSIF x = 3153 THEN
            tanh_f := 1867;
        ELSIF x = 3154 THEN
            tanh_f := 1867;
        ELSIF x = 3155 THEN
            tanh_f := 1867;
        ELSIF x = 3156 THEN
            tanh_f := 1867;
        ELSIF x = 3157 THEN
            tanh_f := 1867;
        ELSIF x = 3158 THEN
            tanh_f := 1868;
        ELSIF x = 3159 THEN
            tanh_f := 1868;
        ELSIF x = 3160 THEN
            tanh_f := 1868;
        ELSIF x = 3161 THEN
            tanh_f := 1868;
        ELSIF x = 3162 THEN
            tanh_f := 1868;
        ELSIF x = 3163 THEN
            tanh_f := 1868;
        ELSIF x = 3164 THEN
            tanh_f := 1869;
        ELSIF x = 3165 THEN
            tanh_f := 1869;
        ELSIF x = 3166 THEN
            tanh_f := 1869;
        ELSIF x = 3167 THEN
            tanh_f := 1869;
        ELSIF x = 3168 THEN
            tanh_f := 1869;
        ELSIF x = 3169 THEN
            tanh_f := 1869;
        ELSIF x = 3170 THEN
            tanh_f := 1870;
        ELSIF x = 3171 THEN
            tanh_f := 1870;
        ELSIF x = 3172 THEN
            tanh_f := 1870;
        ELSIF x = 3173 THEN
            tanh_f := 1870;
        ELSIF x = 3174 THEN
            tanh_f := 1870;
        ELSIF x = 3175 THEN
            tanh_f := 1870;
        ELSIF x = 3176 THEN
            tanh_f := 1871;
        ELSIF x = 3177 THEN
            tanh_f := 1871;
        ELSIF x = 3178 THEN
            tanh_f := 1871;
        ELSIF x = 3179 THEN
            tanh_f := 1871;
        ELSIF x = 3180 THEN
            tanh_f := 1871;
        ELSIF x = 3181 THEN
            tanh_f := 1871;
        ELSIF x = 3182 THEN
            tanh_f := 1872;
        ELSIF x = 3183 THEN
            tanh_f := 1872;
        ELSIF x = 3184 THEN
            tanh_f := 1872;
        ELSIF x = 3185 THEN
            tanh_f := 1872;
        ELSIF x = 3186 THEN
            tanh_f := 1872;
        ELSIF x = 3187 THEN
            tanh_f := 1872;
        ELSIF x = 3188 THEN
            tanh_f := 1873;
        ELSIF x = 3189 THEN
            tanh_f := 1873;
        ELSIF x = 3190 THEN
            tanh_f := 1873;
        ELSIF x = 3191 THEN
            tanh_f := 1873;
        ELSIF x = 3192 THEN
            tanh_f := 1873;
        ELSIF x = 3193 THEN
            tanh_f := 1873;
        ELSIF x = 3194 THEN
            tanh_f := 1874;
        ELSIF x = 3195 THEN
            tanh_f := 1874;
        ELSIF x = 3196 THEN
            tanh_f := 1874;
        ELSIF x = 3197 THEN
            tanh_f := 1874;
        ELSIF x = 3198 THEN
            tanh_f := 1874;
        ELSIF x = 3199 THEN
            tanh_f := 1874;
        ELSIF x = 3200 THEN
            tanh_f := 1875;
        ELSIF x = 3201 THEN
            tanh_f := 1875;
        ELSIF x = 3202 THEN
            tanh_f := 1875;
        ELSIF x = 3203 THEN
            tanh_f := 1875;
        ELSIF x = 3204 THEN
            tanh_f := 1875;
        ELSIF x = 3205 THEN
            tanh_f := 1875;
        ELSIF x = 3206 THEN
            tanh_f := 1875;
        ELSIF x = 3207 THEN
            tanh_f := 1876;
        ELSIF x = 3208 THEN
            tanh_f := 1876;
        ELSIF x = 3209 THEN
            tanh_f := 1876;
        ELSIF x = 3210 THEN
            tanh_f := 1876;
        ELSIF x = 3211 THEN
            tanh_f := 1876;
        ELSIF x = 3212 THEN
            tanh_f := 1876;
        ELSIF x = 3213 THEN
            tanh_f := 1877;
        ELSIF x = 3214 THEN
            tanh_f := 1877;
        ELSIF x = 3215 THEN
            tanh_f := 1877;
        ELSIF x = 3216 THEN
            tanh_f := 1877;
        ELSIF x = 3217 THEN
            tanh_f := 1877;
        ELSIF x = 3218 THEN
            tanh_f := 1877;
        ELSIF x = 3219 THEN
            tanh_f := 1878;
        ELSIF x = 3220 THEN
            tanh_f := 1878;
        ELSIF x = 3221 THEN
            tanh_f := 1878;
        ELSIF x = 3222 THEN
            tanh_f := 1878;
        ELSIF x = 3223 THEN
            tanh_f := 1878;
        ELSIF x = 3224 THEN
            tanh_f := 1878;
        ELSIF x = 3225 THEN
            tanh_f := 1879;
        ELSIF x = 3226 THEN
            tanh_f := 1879;
        ELSIF x = 3227 THEN
            tanh_f := 1879;
        ELSIF x = 3228 THEN
            tanh_f := 1879;
        ELSIF x = 3229 THEN
            tanh_f := 1879;
        ELSIF x = 3230 THEN
            tanh_f := 1879;
        ELSIF x = 3231 THEN
            tanh_f := 1880;
        ELSIF x = 3232 THEN
            tanh_f := 1880;
        ELSIF x = 3233 THEN
            tanh_f := 1880;
        ELSIF x = 3234 THEN
            tanh_f := 1880;
        ELSIF x = 3235 THEN
            tanh_f := 1880;
        ELSIF x = 3236 THEN
            tanh_f := 1880;
        ELSIF x = 3237 THEN
            tanh_f := 1881;
        ELSIF x = 3238 THEN
            tanh_f := 1881;
        ELSIF x = 3239 THEN
            tanh_f := 1881;
        ELSIF x = 3240 THEN
            tanh_f := 1881;
        ELSIF x = 3241 THEN
            tanh_f := 1881;
        ELSIF x = 3242 THEN
            tanh_f := 1881;
        ELSIF x = 3243 THEN
            tanh_f := 1882;
        ELSIF x = 3244 THEN
            tanh_f := 1882;
        ELSIF x = 3245 THEN
            tanh_f := 1882;
        ELSIF x = 3246 THEN
            tanh_f := 1882;
        ELSIF x = 3247 THEN
            tanh_f := 1882;
        ELSIF x = 3248 THEN
            tanh_f := 1882;
        ELSIF x = 3249 THEN
            tanh_f := 1883;
        ELSIF x = 3250 THEN
            tanh_f := 1883;
        ELSIF x = 3251 THEN
            tanh_f := 1883;
        ELSIF x = 3252 THEN
            tanh_f := 1883;
        ELSIF x = 3253 THEN
            tanh_f := 1883;
        ELSIF x = 3254 THEN
            tanh_f := 1883;
        ELSIF x = 3255 THEN
            tanh_f := 1884;
        ELSIF x = 3256 THEN
            tanh_f := 1884;
        ELSIF x = 3257 THEN
            tanh_f := 1884;
        ELSIF x = 3258 THEN
            tanh_f := 1884;
        ELSIF x = 3259 THEN
            tanh_f := 1884;
        ELSIF x = 3260 THEN
            tanh_f := 1884;
        ELSIF x = 3261 THEN
            tanh_f := 1885;
        ELSIF x = 3262 THEN
            tanh_f := 1885;
        ELSIF x = 3263 THEN
            tanh_f := 1885;
        ELSIF x = 3264 THEN
            tanh_f := 1885;
        ELSIF x = 3265 THEN
            tanh_f := 1885;
        ELSIF x = 3266 THEN
            tanh_f := 1885;
        ELSIF x = 3267 THEN
            tanh_f := 1885;
        ELSIF x = 3268 THEN
            tanh_f := 1886;
        ELSIF x = 3269 THEN
            tanh_f := 1886;
        ELSIF x = 3270 THEN
            tanh_f := 1886;
        ELSIF x = 3271 THEN
            tanh_f := 1886;
        ELSIF x = 3272 THEN
            tanh_f := 1886;
        ELSIF x = 3273 THEN
            tanh_f := 1886;
        ELSIF x = 3274 THEN
            tanh_f := 1887;
        ELSIF x = 3275 THEN
            tanh_f := 1887;
        ELSIF x = 3276 THEN
            tanh_f := 1887;
        ELSIF x = 3277 THEN
            tanh_f := 1887;
        ELSIF x = 3278 THEN
            tanh_f := 1887;
        ELSIF x = 3279 THEN
            tanh_f := 1887;
        ELSIF x = 3280 THEN
            tanh_f := 1888;
        ELSIF x = 3281 THEN
            tanh_f := 1888;
        ELSIF x = 3282 THEN
            tanh_f := 1888;
        ELSIF x = 3283 THEN
            tanh_f := 1888;
        ELSIF x = 3284 THEN
            tanh_f := 1888;
        ELSIF x = 3285 THEN
            tanh_f := 1888;
        ELSIF x = 3286 THEN
            tanh_f := 1889;
        ELSIF x = 3287 THEN
            tanh_f := 1889;
        ELSIF x = 3288 THEN
            tanh_f := 1889;
        ELSIF x = 3289 THEN
            tanh_f := 1889;
        ELSIF x = 3290 THEN
            tanh_f := 1889;
        ELSIF x = 3291 THEN
            tanh_f := 1889;
        ELSIF x = 3292 THEN
            tanh_f := 1890;
        ELSIF x = 3293 THEN
            tanh_f := 1890;
        ELSIF x = 3294 THEN
            tanh_f := 1890;
        ELSIF x = 3295 THEN
            tanh_f := 1890;
        ELSIF x = 3296 THEN
            tanh_f := 1890;
        ELSIF x = 3297 THEN
            tanh_f := 1890;
        ELSIF x = 3298 THEN
            tanh_f := 1891;
        ELSIF x = 3299 THEN
            tanh_f := 1891;
        ELSIF x = 3300 THEN
            tanh_f := 1891;
        ELSIF x = 3301 THEN
            tanh_f := 1891;
        ELSIF x = 3302 THEN
            tanh_f := 1891;
        ELSIF x = 3303 THEN
            tanh_f := 1891;
        ELSIF x = 3304 THEN
            tanh_f := 1892;
        ELSIF x = 3305 THEN
            tanh_f := 1892;
        ELSIF x = 3306 THEN
            tanh_f := 1892;
        ELSIF x = 3307 THEN
            tanh_f := 1892;
        ELSIF x = 3308 THEN
            tanh_f := 1892;
        ELSIF x = 3309 THEN
            tanh_f := 1892;
        ELSIF x = 3310 THEN
            tanh_f := 1893;
        ELSIF x = 3311 THEN
            tanh_f := 1893;
        ELSIF x = 3312 THEN
            tanh_f := 1893;
        ELSIF x = 3313 THEN
            tanh_f := 1893;
        ELSIF x = 3314 THEN
            tanh_f := 1893;
        ELSIF x = 3315 THEN
            tanh_f := 1893;
        ELSIF x = 3316 THEN
            tanh_f := 1894;
        ELSIF x = 3317 THEN
            tanh_f := 1894;
        ELSIF x = 3318 THEN
            tanh_f := 1894;
        ELSIF x = 3319 THEN
            tanh_f := 1894;
        ELSIF x = 3320 THEN
            tanh_f := 1894;
        ELSIF x = 3321 THEN
            tanh_f := 1894;
        ELSIF x = 3322 THEN
            tanh_f := 1895;
        ELSIF x = 3323 THEN
            tanh_f := 1895;
        ELSIF x = 3324 THEN
            tanh_f := 1895;
        ELSIF x = 3325 THEN
            tanh_f := 1895;
        ELSIF x = 3326 THEN
            tanh_f := 1895;
        ELSIF x = 3327 THEN
            tanh_f := 1895;
        ELSIF x = 3328 THEN
            tanh_f := 1896;
        ELSIF x = 3329 THEN
            tanh_f := 1896;
        ELSIF x = 3330 THEN
            tanh_f := 1896;
        ELSIF x = 3331 THEN
            tanh_f := 1896;
        ELSIF x = 3332 THEN
            tanh_f := 1896;
        ELSIF x = 3333 THEN
            tanh_f := 1896;
        ELSIF x = 3334 THEN
            tanh_f := 1896;
        ELSIF x = 3335 THEN
            tanh_f := 1896;
        ELSIF x = 3336 THEN
            tanh_f := 1897;
        ELSIF x = 3337 THEN
            tanh_f := 1897;
        ELSIF x = 3338 THEN
            tanh_f := 1897;
        ELSIF x = 3339 THEN
            tanh_f := 1897;
        ELSIF x = 3340 THEN
            tanh_f := 1897;
        ELSIF x = 3341 THEN
            tanh_f := 1897;
        ELSIF x = 3342 THEN
            tanh_f := 1897;
        ELSIF x = 3343 THEN
            tanh_f := 1897;
        ELSIF x = 3344 THEN
            tanh_f := 1898;
        ELSIF x = 3345 THEN
            tanh_f := 1898;
        ELSIF x = 3346 THEN
            tanh_f := 1898;
        ELSIF x = 3347 THEN
            tanh_f := 1898;
        ELSIF x = 3348 THEN
            tanh_f := 1898;
        ELSIF x = 3349 THEN
            tanh_f := 1898;
        ELSIF x = 3350 THEN
            tanh_f := 1898;
        ELSIF x = 3351 THEN
            tanh_f := 1898;
        ELSIF x = 3352 THEN
            tanh_f := 1899;
        ELSIF x = 3353 THEN
            tanh_f := 1899;
        ELSIF x = 3354 THEN
            tanh_f := 1899;
        ELSIF x = 3355 THEN
            tanh_f := 1899;
        ELSIF x = 3356 THEN
            tanh_f := 1899;
        ELSIF x = 3357 THEN
            tanh_f := 1899;
        ELSIF x = 3358 THEN
            tanh_f := 1899;
        ELSIF x = 3359 THEN
            tanh_f := 1899;
        ELSIF x = 3360 THEN
            tanh_f := 1900;
        ELSIF x = 3361 THEN
            tanh_f := 1900;
        ELSIF x = 3362 THEN
            tanh_f := 1900;
        ELSIF x = 3363 THEN
            tanh_f := 1900;
        ELSIF x = 3364 THEN
            tanh_f := 1900;
        ELSIF x = 3365 THEN
            tanh_f := 1900;
        ELSIF x = 3366 THEN
            tanh_f := 1900;
        ELSIF x = 3367 THEN
            tanh_f := 1900;
        ELSIF x = 3368 THEN
            tanh_f := 1901;
        ELSIF x = 3369 THEN
            tanh_f := 1901;
        ELSIF x = 3370 THEN
            tanh_f := 1901;
        ELSIF x = 3371 THEN
            tanh_f := 1901;
        ELSIF x = 3372 THEN
            tanh_f := 1901;
        ELSIF x = 3373 THEN
            tanh_f := 1901;
        ELSIF x = 3374 THEN
            tanh_f := 1901;
        ELSIF x = 3375 THEN
            tanh_f := 1901;
        ELSIF x = 3376 THEN
            tanh_f := 1902;
        ELSIF x = 3377 THEN
            tanh_f := 1902;
        ELSIF x = 3378 THEN
            tanh_f := 1902;
        ELSIF x = 3379 THEN
            tanh_f := 1902;
        ELSIF x = 3380 THEN
            tanh_f := 1902;
        ELSIF x = 3381 THEN
            tanh_f := 1902;
        ELSIF x = 3382 THEN
            tanh_f := 1902;
        ELSIF x = 3383 THEN
            tanh_f := 1902;
        ELSIF x = 3384 THEN
            tanh_f := 1903;
        ELSIF x = 3385 THEN
            tanh_f := 1903;
        ELSIF x = 3386 THEN
            tanh_f := 1903;
        ELSIF x = 3387 THEN
            tanh_f := 1903;
        ELSIF x = 3388 THEN
            tanh_f := 1903;
        ELSIF x = 3389 THEN
            tanh_f := 1903;
        ELSIF x = 3390 THEN
            tanh_f := 1903;
        ELSIF x = 3391 THEN
            tanh_f := 1903;
        ELSIF x = 3392 THEN
            tanh_f := 1904;
        ELSIF x = 3393 THEN
            tanh_f := 1904;
        ELSIF x = 3394 THEN
            tanh_f := 1904;
        ELSIF x = 3395 THEN
            tanh_f := 1904;
        ELSIF x = 3396 THEN
            tanh_f := 1904;
        ELSIF x = 3397 THEN
            tanh_f := 1904;
        ELSIF x = 3398 THEN
            tanh_f := 1904;
        ELSIF x = 3399 THEN
            tanh_f := 1904;
        ELSIF x = 3400 THEN
            tanh_f := 1905;
        ELSIF x = 3401 THEN
            tanh_f := 1905;
        ELSIF x = 3402 THEN
            tanh_f := 1905;
        ELSIF x = 3403 THEN
            tanh_f := 1905;
        ELSIF x = 3404 THEN
            tanh_f := 1905;
        ELSIF x = 3405 THEN
            tanh_f := 1905;
        ELSIF x = 3406 THEN
            tanh_f := 1905;
        ELSIF x = 3407 THEN
            tanh_f := 1905;
        ELSIF x = 3408 THEN
            tanh_f := 1906;
        ELSIF x = 3409 THEN
            tanh_f := 1906;
        ELSIF x = 3410 THEN
            tanh_f := 1906;
        ELSIF x = 3411 THEN
            tanh_f := 1906;
        ELSIF x = 3412 THEN
            tanh_f := 1906;
        ELSIF x = 3413 THEN
            tanh_f := 1906;
        ELSIF x = 3414 THEN
            tanh_f := 1906;
        ELSIF x = 3415 THEN
            tanh_f := 1906;
        ELSIF x = 3416 THEN
            tanh_f := 1907;
        ELSIF x = 3417 THEN
            tanh_f := 1907;
        ELSIF x = 3418 THEN
            tanh_f := 1907;
        ELSIF x = 3419 THEN
            tanh_f := 1907;
        ELSIF x = 3420 THEN
            tanh_f := 1907;
        ELSIF x = 3421 THEN
            tanh_f := 1907;
        ELSIF x = 3422 THEN
            tanh_f := 1907;
        ELSIF x = 3423 THEN
            tanh_f := 1907;
        ELSIF x = 3424 THEN
            tanh_f := 1908;
        ELSIF x = 3425 THEN
            tanh_f := 1908;
        ELSIF x = 3426 THEN
            tanh_f := 1908;
        ELSIF x = 3427 THEN
            tanh_f := 1908;
        ELSIF x = 3428 THEN
            tanh_f := 1908;
        ELSIF x = 3429 THEN
            tanh_f := 1908;
        ELSIF x = 3430 THEN
            tanh_f := 1908;
        ELSIF x = 3431 THEN
            tanh_f := 1908;
        ELSIF x = 3432 THEN
            tanh_f := 1909;
        ELSIF x = 3433 THEN
            tanh_f := 1909;
        ELSIF x = 3434 THEN
            tanh_f := 1909;
        ELSIF x = 3435 THEN
            tanh_f := 1909;
        ELSIF x = 3436 THEN
            tanh_f := 1909;
        ELSIF x = 3437 THEN
            tanh_f := 1909;
        ELSIF x = 3438 THEN
            tanh_f := 1909;
        ELSIF x = 3439 THEN
            tanh_f := 1909;
        ELSIF x = 3440 THEN
            tanh_f := 1910;
        ELSIF x = 3441 THEN
            tanh_f := 1910;
        ELSIF x = 3442 THEN
            tanh_f := 1910;
        ELSIF x = 3443 THEN
            tanh_f := 1910;
        ELSIF x = 3444 THEN
            tanh_f := 1910;
        ELSIF x = 3445 THEN
            tanh_f := 1910;
        ELSIF x = 3446 THEN
            tanh_f := 1910;
        ELSIF x = 3447 THEN
            tanh_f := 1910;
        ELSIF x = 3448 THEN
            tanh_f := 1911;
        ELSIF x = 3449 THEN
            tanh_f := 1911;
        ELSIF x = 3450 THEN
            tanh_f := 1911;
        ELSIF x = 3451 THEN
            tanh_f := 1911;
        ELSIF x = 3452 THEN
            tanh_f := 1911;
        ELSIF x = 3453 THEN
            tanh_f := 1911;
        ELSIF x = 3454 THEN
            tanh_f := 1911;
        ELSIF x = 3455 THEN
            tanh_f := 1911;
        ELSIF x = 3456 THEN
            tanh_f := 1912;
        ELSIF x = 3457 THEN
            tanh_f := 1912;
        ELSIF x = 3458 THEN
            tanh_f := 1912;
        ELSIF x = 3459 THEN
            tanh_f := 1912;
        ELSIF x = 3460 THEN
            tanh_f := 1912;
        ELSIF x = 3461 THEN
            tanh_f := 1912;
        ELSIF x = 3462 THEN
            tanh_f := 1912;
        ELSIF x = 3463 THEN
            tanh_f := 1912;
        ELSIF x = 3464 THEN
            tanh_f := 1913;
        ELSIF x = 3465 THEN
            tanh_f := 1913;
        ELSIF x = 3466 THEN
            tanh_f := 1913;
        ELSIF x = 3467 THEN
            tanh_f := 1913;
        ELSIF x = 3468 THEN
            tanh_f := 1913;
        ELSIF x = 3469 THEN
            tanh_f := 1913;
        ELSIF x = 3470 THEN
            tanh_f := 1913;
        ELSIF x = 3471 THEN
            tanh_f := 1913;
        ELSIF x = 3472 THEN
            tanh_f := 1914;
        ELSIF x = 3473 THEN
            tanh_f := 1914;
        ELSIF x = 3474 THEN
            tanh_f := 1914;
        ELSIF x = 3475 THEN
            tanh_f := 1914;
        ELSIF x = 3476 THEN
            tanh_f := 1914;
        ELSIF x = 3477 THEN
            tanh_f := 1914;
        ELSIF x = 3478 THEN
            tanh_f := 1914;
        ELSIF x = 3479 THEN
            tanh_f := 1914;
        ELSIF x = 3480 THEN
            tanh_f := 1915;
        ELSIF x = 3481 THEN
            tanh_f := 1915;
        ELSIF x = 3482 THEN
            tanh_f := 1915;
        ELSIF x = 3483 THEN
            tanh_f := 1915;
        ELSIF x = 3484 THEN
            tanh_f := 1915;
        ELSIF x = 3485 THEN
            tanh_f := 1915;
        ELSIF x = 3486 THEN
            tanh_f := 1915;
        ELSIF x = 3487 THEN
            tanh_f := 1915;
        ELSIF x = 3488 THEN
            tanh_f := 1916;
        ELSIF x = 3489 THEN
            tanh_f := 1916;
        ELSIF x = 3490 THEN
            tanh_f := 1916;
        ELSIF x = 3491 THEN
            tanh_f := 1916;
        ELSIF x = 3492 THEN
            tanh_f := 1916;
        ELSIF x = 3493 THEN
            tanh_f := 1916;
        ELSIF x = 3494 THEN
            tanh_f := 1916;
        ELSIF x = 3495 THEN
            tanh_f := 1916;
        ELSIF x = 3496 THEN
            tanh_f := 1917;
        ELSIF x = 3497 THEN
            tanh_f := 1917;
        ELSIF x = 3498 THEN
            tanh_f := 1917;
        ELSIF x = 3499 THEN
            tanh_f := 1917;
        ELSIF x = 3500 THEN
            tanh_f := 1917;
        ELSIF x = 3501 THEN
            tanh_f := 1917;
        ELSIF x = 3502 THEN
            tanh_f := 1917;
        ELSIF x = 3503 THEN
            tanh_f := 1917;
        ELSIF x = 3504 THEN
            tanh_f := 1918;
        ELSIF x = 3505 THEN
            tanh_f := 1918;
        ELSIF x = 3506 THEN
            tanh_f := 1918;
        ELSIF x = 3507 THEN
            tanh_f := 1918;
        ELSIF x = 3508 THEN
            tanh_f := 1918;
        ELSIF x = 3509 THEN
            tanh_f := 1918;
        ELSIF x = 3510 THEN
            tanh_f := 1918;
        ELSIF x = 3511 THEN
            tanh_f := 1918;
        ELSIF x = 3512 THEN
            tanh_f := 1919;
        ELSIF x = 3513 THEN
            tanh_f := 1919;
        ELSIF x = 3514 THEN
            tanh_f := 1919;
        ELSIF x = 3515 THEN
            tanh_f := 1919;
        ELSIF x = 3516 THEN
            tanh_f := 1919;
        ELSIF x = 3517 THEN
            tanh_f := 1919;
        ELSIF x = 3518 THEN
            tanh_f := 1919;
        ELSIF x = 3519 THEN
            tanh_f := 1919;
        ELSIF x = 3520 THEN
            tanh_f := 1920;
        ELSIF x = 3521 THEN
            tanh_f := 1920;
        ELSIF x = 3522 THEN
            tanh_f := 1920;
        ELSIF x = 3523 THEN
            tanh_f := 1920;
        ELSIF x = 3524 THEN
            tanh_f := 1920;
        ELSIF x = 3525 THEN
            tanh_f := 1920;
        ELSIF x = 3526 THEN
            tanh_f := 1920;
        ELSIF x = 3527 THEN
            tanh_f := 1920;
        ELSIF x = 3528 THEN
            tanh_f := 1921;
        ELSIF x = 3529 THEN
            tanh_f := 1921;
        ELSIF x = 3530 THEN
            tanh_f := 1921;
        ELSIF x = 3531 THEN
            tanh_f := 1921;
        ELSIF x = 3532 THEN
            tanh_f := 1921;
        ELSIF x = 3533 THEN
            tanh_f := 1921;
        ELSIF x = 3534 THEN
            tanh_f := 1921;
        ELSIF x = 3535 THEN
            tanh_f := 1921;
        ELSIF x = 3536 THEN
            tanh_f := 1922;
        ELSIF x = 3537 THEN
            tanh_f := 1922;
        ELSIF x = 3538 THEN
            tanh_f := 1922;
        ELSIF x = 3539 THEN
            tanh_f := 1922;
        ELSIF x = 3540 THEN
            tanh_f := 1922;
        ELSIF x = 3541 THEN
            tanh_f := 1922;
        ELSIF x = 3542 THEN
            tanh_f := 1922;
        ELSIF x = 3543 THEN
            tanh_f := 1922;
        ELSIF x = 3544 THEN
            tanh_f := 1923;
        ELSIF x = 3545 THEN
            tanh_f := 1923;
        ELSIF x = 3546 THEN
            tanh_f := 1923;
        ELSIF x = 3547 THEN
            tanh_f := 1923;
        ELSIF x = 3548 THEN
            tanh_f := 1923;
        ELSIF x = 3549 THEN
            tanh_f := 1923;
        ELSIF x = 3550 THEN
            tanh_f := 1923;
        ELSIF x = 3551 THEN
            tanh_f := 1923;
        ELSIF x = 3552 THEN
            tanh_f := 1924;
        ELSIF x = 3553 THEN
            tanh_f := 1924;
        ELSIF x = 3554 THEN
            tanh_f := 1924;
        ELSIF x = 3555 THEN
            tanh_f := 1924;
        ELSIF x = 3556 THEN
            tanh_f := 1924;
        ELSIF x = 3557 THEN
            tanh_f := 1924;
        ELSIF x = 3558 THEN
            tanh_f := 1924;
        ELSIF x = 3559 THEN
            tanh_f := 1924;
        ELSIF x = 3560 THEN
            tanh_f := 1925;
        ELSIF x = 3561 THEN
            tanh_f := 1925;
        ELSIF x = 3562 THEN
            tanh_f := 1925;
        ELSIF x = 3563 THEN
            tanh_f := 1925;
        ELSIF x = 3564 THEN
            tanh_f := 1925;
        ELSIF x = 3565 THEN
            tanh_f := 1925;
        ELSIF x = 3566 THEN
            tanh_f := 1925;
        ELSIF x = 3567 THEN
            tanh_f := 1925;
        ELSIF x = 3568 THEN
            tanh_f := 1926;
        ELSIF x = 3569 THEN
            tanh_f := 1926;
        ELSIF x = 3570 THEN
            tanh_f := 1926;
        ELSIF x = 3571 THEN
            tanh_f := 1926;
        ELSIF x = 3572 THEN
            tanh_f := 1926;
        ELSIF x = 3573 THEN
            tanh_f := 1926;
        ELSIF x = 3574 THEN
            tanh_f := 1926;
        ELSIF x = 3575 THEN
            tanh_f := 1926;
        ELSIF x = 3576 THEN
            tanh_f := 1927;
        ELSIF x = 3577 THEN
            tanh_f := 1927;
        ELSIF x = 3578 THEN
            tanh_f := 1927;
        ELSIF x = 3579 THEN
            tanh_f := 1927;
        ELSIF x = 3580 THEN
            tanh_f := 1927;
        ELSIF x = 3581 THEN
            tanh_f := 1927;
        ELSIF x = 3582 THEN
            tanh_f := 1927;
        ELSIF x = 3583 THEN
            tanh_f := 1927;
        ELSIF x = 3584 THEN
            tanh_f := 1928;
        ELSIF x = 3585 THEN
            tanh_f := 1928;
        ELSIF x = 3586 THEN
            tanh_f := 1928;
        ELSIF x = 3587 THEN
            tanh_f := 1928;
        ELSIF x = 3588 THEN
            tanh_f := 1928;
        ELSIF x = 3589 THEN
            tanh_f := 1928;
        ELSIF x = 3590 THEN
            tanh_f := 1928;
        ELSIF x = 3591 THEN
            tanh_f := 1928;
        ELSIF x = 3592 THEN
            tanh_f := 1928;
        ELSIF x = 3593 THEN
            tanh_f := 1928;
        ELSIF x = 3594 THEN
            tanh_f := 1929;
        ELSIF x = 3595 THEN
            tanh_f := 1929;
        ELSIF x = 3596 THEN
            tanh_f := 1929;
        ELSIF x = 3597 THEN
            tanh_f := 1929;
        ELSIF x = 3598 THEN
            tanh_f := 1929;
        ELSIF x = 3599 THEN
            tanh_f := 1929;
        ELSIF x = 3600 THEN
            tanh_f := 1929;
        ELSIF x = 3601 THEN
            tanh_f := 1929;
        ELSIF x = 3602 THEN
            tanh_f := 1929;
        ELSIF x = 3603 THEN
            tanh_f := 1930;
        ELSIF x = 3604 THEN
            tanh_f := 1930;
        ELSIF x = 3605 THEN
            tanh_f := 1930;
        ELSIF x = 3606 THEN
            tanh_f := 1930;
        ELSIF x = 3607 THEN
            tanh_f := 1930;
        ELSIF x = 3608 THEN
            tanh_f := 1930;
        ELSIF x = 3609 THEN
            tanh_f := 1930;
        ELSIF x = 3610 THEN
            tanh_f := 1930;
        ELSIF x = 3611 THEN
            tanh_f := 1930;
        ELSIF x = 3612 THEN
            tanh_f := 1930;
        ELSIF x = 3613 THEN
            tanh_f := 1931;
        ELSIF x = 3614 THEN
            tanh_f := 1931;
        ELSIF x = 3615 THEN
            tanh_f := 1931;
        ELSIF x = 3616 THEN
            tanh_f := 1931;
        ELSIF x = 3617 THEN
            tanh_f := 1931;
        ELSIF x = 3618 THEN
            tanh_f := 1931;
        ELSIF x = 3619 THEN
            tanh_f := 1931;
        ELSIF x = 3620 THEN
            tanh_f := 1931;
        ELSIF x = 3621 THEN
            tanh_f := 1931;
        ELSIF x = 3622 THEN
            tanh_f := 1932;
        ELSIF x = 3623 THEN
            tanh_f := 1932;
        ELSIF x = 3624 THEN
            tanh_f := 1932;
        ELSIF x = 3625 THEN
            tanh_f := 1932;
        ELSIF x = 3626 THEN
            tanh_f := 1932;
        ELSIF x = 3627 THEN
            tanh_f := 1932;
        ELSIF x = 3628 THEN
            tanh_f := 1932;
        ELSIF x = 3629 THEN
            tanh_f := 1932;
        ELSIF x = 3630 THEN
            tanh_f := 1932;
        ELSIF x = 3631 THEN
            tanh_f := 1932;
        ELSIF x = 3632 THEN
            tanh_f := 1933;
        ELSIF x = 3633 THEN
            tanh_f := 1933;
        ELSIF x = 3634 THEN
            tanh_f := 1933;
        ELSIF x = 3635 THEN
            tanh_f := 1933;
        ELSIF x = 3636 THEN
            tanh_f := 1933;
        ELSIF x = 3637 THEN
            tanh_f := 1933;
        ELSIF x = 3638 THEN
            tanh_f := 1933;
        ELSIF x = 3639 THEN
            tanh_f := 1933;
        ELSIF x = 3640 THEN
            tanh_f := 1933;
        ELSIF x = 3641 THEN
            tanh_f := 1934;
        ELSIF x = 3642 THEN
            tanh_f := 1934;
        ELSIF x = 3643 THEN
            tanh_f := 1934;
        ELSIF x = 3644 THEN
            tanh_f := 1934;
        ELSIF x = 3645 THEN
            tanh_f := 1934;
        ELSIF x = 3646 THEN
            tanh_f := 1934;
        ELSIF x = 3647 THEN
            tanh_f := 1934;
        ELSIF x = 3648 THEN
            tanh_f := 1934;
        ELSIF x = 3649 THEN
            tanh_f := 1934;
        ELSIF x = 3650 THEN
            tanh_f := 1934;
        ELSIF x = 3651 THEN
            tanh_f := 1935;
        ELSIF x = 3652 THEN
            tanh_f := 1935;
        ELSIF x = 3653 THEN
            tanh_f := 1935;
        ELSIF x = 3654 THEN
            tanh_f := 1935;
        ELSIF x = 3655 THEN
            tanh_f := 1935;
        ELSIF x = 3656 THEN
            tanh_f := 1935;
        ELSIF x = 3657 THEN
            tanh_f := 1935;
        ELSIF x = 3658 THEN
            tanh_f := 1935;
        ELSIF x = 3659 THEN
            tanh_f := 1935;
        ELSIF x = 3660 THEN
            tanh_f := 1936;
        ELSIF x = 3661 THEN
            tanh_f := 1936;
        ELSIF x = 3662 THEN
            tanh_f := 1936;
        ELSIF x = 3663 THEN
            tanh_f := 1936;
        ELSIF x = 3664 THEN
            tanh_f := 1936;
        ELSIF x = 3665 THEN
            tanh_f := 1936;
        ELSIF x = 3666 THEN
            tanh_f := 1936;
        ELSIF x = 3667 THEN
            tanh_f := 1936;
        ELSIF x = 3668 THEN
            tanh_f := 1936;
        ELSIF x = 3669 THEN
            tanh_f := 1936;
        ELSIF x = 3670 THEN
            tanh_f := 1937;
        ELSIF x = 3671 THEN
            tanh_f := 1937;
        ELSIF x = 3672 THEN
            tanh_f := 1937;
        ELSIF x = 3673 THEN
            tanh_f := 1937;
        ELSIF x = 3674 THEN
            tanh_f := 1937;
        ELSIF x = 3675 THEN
            tanh_f := 1937;
        ELSIF x = 3676 THEN
            tanh_f := 1937;
        ELSIF x = 3677 THEN
            tanh_f := 1937;
        ELSIF x = 3678 THEN
            tanh_f := 1937;
        ELSIF x = 3679 THEN
            tanh_f := 1938;
        ELSIF x = 3680 THEN
            tanh_f := 1938;
        ELSIF x = 3681 THEN
            tanh_f := 1938;
        ELSIF x = 3682 THEN
            tanh_f := 1938;
        ELSIF x = 3683 THEN
            tanh_f := 1938;
        ELSIF x = 3684 THEN
            tanh_f := 1938;
        ELSIF x = 3685 THEN
            tanh_f := 1938;
        ELSIF x = 3686 THEN
            tanh_f := 1938;
        ELSIF x = 3687 THEN
            tanh_f := 1938;
        ELSIF x = 3688 THEN
            tanh_f := 1938;
        ELSIF x = 3689 THEN
            tanh_f := 1939;
        ELSIF x = 3690 THEN
            tanh_f := 1939;
        ELSIF x = 3691 THEN
            tanh_f := 1939;
        ELSIF x = 3692 THEN
            tanh_f := 1939;
        ELSIF x = 3693 THEN
            tanh_f := 1939;
        ELSIF x = 3694 THEN
            tanh_f := 1939;
        ELSIF x = 3695 THEN
            tanh_f := 1939;
        ELSIF x = 3696 THEN
            tanh_f := 1939;
        ELSIF x = 3697 THEN
            tanh_f := 1939;
        ELSIF x = 3698 THEN
            tanh_f := 1940;
        ELSIF x = 3699 THEN
            tanh_f := 1940;
        ELSIF x = 3700 THEN
            tanh_f := 1940;
        ELSIF x = 3701 THEN
            tanh_f := 1940;
        ELSIF x = 3702 THEN
            tanh_f := 1940;
        ELSIF x = 3703 THEN
            tanh_f := 1940;
        ELSIF x = 3704 THEN
            tanh_f := 1940;
        ELSIF x = 3705 THEN
            tanh_f := 1940;
        ELSIF x = 3706 THEN
            tanh_f := 1940;
        ELSIF x = 3707 THEN
            tanh_f := 1940;
        ELSIF x = 3708 THEN
            tanh_f := 1941;
        ELSIF x = 3709 THEN
            tanh_f := 1941;
        ELSIF x = 3710 THEN
            tanh_f := 1941;
        ELSIF x = 3711 THEN
            tanh_f := 1941;
        ELSIF x = 3712 THEN
            tanh_f := 1941;
        ELSIF x = 3713 THEN
            tanh_f := 1941;
        ELSIF x = 3714 THEN
            tanh_f := 1941;
        ELSIF x = 3715 THEN
            tanh_f := 1941;
        ELSIF x = 3716 THEN
            tanh_f := 1941;
        ELSIF x = 3717 THEN
            tanh_f := 1942;
        ELSIF x = 3718 THEN
            tanh_f := 1942;
        ELSIF x = 3719 THEN
            tanh_f := 1942;
        ELSIF x = 3720 THEN
            tanh_f := 1942;
        ELSIF x = 3721 THEN
            tanh_f := 1942;
        ELSIF x = 3722 THEN
            tanh_f := 1942;
        ELSIF x = 3723 THEN
            tanh_f := 1942;
        ELSIF x = 3724 THEN
            tanh_f := 1942;
        ELSIF x = 3725 THEN
            tanh_f := 1942;
        ELSIF x = 3726 THEN
            tanh_f := 1942;
        ELSIF x = 3727 THEN
            tanh_f := 1943;
        ELSIF x = 3728 THEN
            tanh_f := 1943;
        ELSIF x = 3729 THEN
            tanh_f := 1943;
        ELSIF x = 3730 THEN
            tanh_f := 1943;
        ELSIF x = 3731 THEN
            tanh_f := 1943;
        ELSIF x = 3732 THEN
            tanh_f := 1943;
        ELSIF x = 3733 THEN
            tanh_f := 1943;
        ELSIF x = 3734 THEN
            tanh_f := 1943;
        ELSIF x = 3735 THEN
            tanh_f := 1943;
        ELSIF x = 3736 THEN
            tanh_f := 1944;
        ELSIF x = 3737 THEN
            tanh_f := 1944;
        ELSIF x = 3738 THEN
            tanh_f := 1944;
        ELSIF x = 3739 THEN
            tanh_f := 1944;
        ELSIF x = 3740 THEN
            tanh_f := 1944;
        ELSIF x = 3741 THEN
            tanh_f := 1944;
        ELSIF x = 3742 THEN
            tanh_f := 1944;
        ELSIF x = 3743 THEN
            tanh_f := 1944;
        ELSIF x = 3744 THEN
            tanh_f := 1944;
        ELSIF x = 3745 THEN
            tanh_f := 1944;
        ELSIF x = 3746 THEN
            tanh_f := 1945;
        ELSIF x = 3747 THEN
            tanh_f := 1945;
        ELSIF x = 3748 THEN
            tanh_f := 1945;
        ELSIF x = 3749 THEN
            tanh_f := 1945;
        ELSIF x = 3750 THEN
            tanh_f := 1945;
        ELSIF x = 3751 THEN
            tanh_f := 1945;
        ELSIF x = 3752 THEN
            tanh_f := 1945;
        ELSIF x = 3753 THEN
            tanh_f := 1945;
        ELSIF x = 3754 THEN
            tanh_f := 1945;
        ELSIF x = 3755 THEN
            tanh_f := 1946;
        ELSIF x = 3756 THEN
            tanh_f := 1946;
        ELSIF x = 3757 THEN
            tanh_f := 1946;
        ELSIF x = 3758 THEN
            tanh_f := 1946;
        ELSIF x = 3759 THEN
            tanh_f := 1946;
        ELSIF x = 3760 THEN
            tanh_f := 1946;
        ELSIF x = 3761 THEN
            tanh_f := 1946;
        ELSIF x = 3762 THEN
            tanh_f := 1946;
        ELSIF x = 3763 THEN
            tanh_f := 1946;
        ELSIF x = 3764 THEN
            tanh_f := 1946;
        ELSIF x = 3765 THEN
            tanh_f := 1947;
        ELSIF x = 3766 THEN
            tanh_f := 1947;
        ELSIF x = 3767 THEN
            tanh_f := 1947;
        ELSIF x = 3768 THEN
            tanh_f := 1947;
        ELSIF x = 3769 THEN
            tanh_f := 1947;
        ELSIF x = 3770 THEN
            tanh_f := 1947;
        ELSIF x = 3771 THEN
            tanh_f := 1947;
        ELSIF x = 3772 THEN
            tanh_f := 1947;
        ELSIF x = 3773 THEN
            tanh_f := 1947;
        ELSIF x = 3774 THEN
            tanh_f := 1948;
        ELSIF x = 3775 THEN
            tanh_f := 1948;
        ELSIF x = 3776 THEN
            tanh_f := 1948;
        ELSIF x = 3777 THEN
            tanh_f := 1948;
        ELSIF x = 3778 THEN
            tanh_f := 1948;
        ELSIF x = 3779 THEN
            tanh_f := 1948;
        ELSIF x = 3780 THEN
            tanh_f := 1948;
        ELSIF x = 3781 THEN
            tanh_f := 1948;
        ELSIF x = 3782 THEN
            tanh_f := 1948;
        ELSIF x = 3783 THEN
            tanh_f := 1948;
        ELSIF x = 3784 THEN
            tanh_f := 1949;
        ELSIF x = 3785 THEN
            tanh_f := 1949;
        ELSIF x = 3786 THEN
            tanh_f := 1949;
        ELSIF x = 3787 THEN
            tanh_f := 1949;
        ELSIF x = 3788 THEN
            tanh_f := 1949;
        ELSIF x = 3789 THEN
            tanh_f := 1949;
        ELSIF x = 3790 THEN
            tanh_f := 1949;
        ELSIF x = 3791 THEN
            tanh_f := 1949;
        ELSIF x = 3792 THEN
            tanh_f := 1949;
        ELSIF x = 3793 THEN
            tanh_f := 1950;
        ELSIF x = 3794 THEN
            tanh_f := 1950;
        ELSIF x = 3795 THEN
            tanh_f := 1950;
        ELSIF x = 3796 THEN
            tanh_f := 1950;
        ELSIF x = 3797 THEN
            tanh_f := 1950;
        ELSIF x = 3798 THEN
            tanh_f := 1950;
        ELSIF x = 3799 THEN
            tanh_f := 1950;
        ELSIF x = 3800 THEN
            tanh_f := 1950;
        ELSIF x = 3801 THEN
            tanh_f := 1950;
        ELSIF x = 3802 THEN
            tanh_f := 1950;
        ELSIF x = 3803 THEN
            tanh_f := 1951;
        ELSIF x = 3804 THEN
            tanh_f := 1951;
        ELSIF x = 3805 THEN
            tanh_f := 1951;
        ELSIF x = 3806 THEN
            tanh_f := 1951;
        ELSIF x = 3807 THEN
            tanh_f := 1951;
        ELSIF x = 3808 THEN
            tanh_f := 1951;
        ELSIF x = 3809 THEN
            tanh_f := 1951;
        ELSIF x = 3810 THEN
            tanh_f := 1951;
        ELSIF x = 3811 THEN
            tanh_f := 1951;
        ELSIF x = 3812 THEN
            tanh_f := 1952;
        ELSIF x = 3813 THEN
            tanh_f := 1952;
        ELSIF x = 3814 THEN
            tanh_f := 1952;
        ELSIF x = 3815 THEN
            tanh_f := 1952;
        ELSIF x = 3816 THEN
            tanh_f := 1952;
        ELSIF x = 3817 THEN
            tanh_f := 1952;
        ELSIF x = 3818 THEN
            tanh_f := 1952;
        ELSIF x = 3819 THEN
            tanh_f := 1952;
        ELSIF x = 3820 THEN
            tanh_f := 1952;
        ELSIF x = 3821 THEN
            tanh_f := 1952;
        ELSIF x = 3822 THEN
            tanh_f := 1953;
        ELSIF x = 3823 THEN
            tanh_f := 1953;
        ELSIF x = 3824 THEN
            tanh_f := 1953;
        ELSIF x = 3825 THEN
            tanh_f := 1953;
        ELSIF x = 3826 THEN
            tanh_f := 1953;
        ELSIF x = 3827 THEN
            tanh_f := 1953;
        ELSIF x = 3828 THEN
            tanh_f := 1953;
        ELSIF x = 3829 THEN
            tanh_f := 1953;
        ELSIF x = 3830 THEN
            tanh_f := 1953;
        ELSIF x = 3831 THEN
            tanh_f := 1954;
        ELSIF x = 3832 THEN
            tanh_f := 1954;
        ELSIF x = 3833 THEN
            tanh_f := 1954;
        ELSIF x = 3834 THEN
            tanh_f := 1954;
        ELSIF x = 3835 THEN
            tanh_f := 1954;
        ELSIF x = 3836 THEN
            tanh_f := 1954;
        ELSIF x = 3837 THEN
            tanh_f := 1954;
        ELSIF x = 3838 THEN
            tanh_f := 1954;
        ELSIF x = 3839 THEN
            tanh_f := 1954;
        ELSIF x = 3840 THEN
            tanh_f := 1954;
        ELSIF x = 3841 THEN
            tanh_f := 1954;
        ELSIF x = 3842 THEN
            tanh_f := 1954;
        ELSIF x = 3843 THEN
            tanh_f := 1954;
        ELSIF x = 3844 THEN
            tanh_f := 1954;
        ELSIF x = 3845 THEN
            tanh_f := 1954;
        ELSIF x = 3846 THEN
            tanh_f := 1954;
        ELSIF x = 3847 THEN
            tanh_f := 1955;
        ELSIF x = 3848 THEN
            tanh_f := 1955;
        ELSIF x = 3849 THEN
            tanh_f := 1955;
        ELSIF x = 3850 THEN
            tanh_f := 1955;
        ELSIF x = 3851 THEN
            tanh_f := 1955;
        ELSIF x = 3852 THEN
            tanh_f := 1955;
        ELSIF x = 3853 THEN
            tanh_f := 1955;
        ELSIF x = 3854 THEN
            tanh_f := 1955;
        ELSIF x = 3855 THEN
            tanh_f := 1955;
        ELSIF x = 3856 THEN
            tanh_f := 1955;
        ELSIF x = 3857 THEN
            tanh_f := 1955;
        ELSIF x = 3858 THEN
            tanh_f := 1955;
        ELSIF x = 3859 THEN
            tanh_f := 1955;
        ELSIF x = 3860 THEN
            tanh_f := 1956;
        ELSIF x = 3861 THEN
            tanh_f := 1956;
        ELSIF x = 3862 THEN
            tanh_f := 1956;
        ELSIF x = 3863 THEN
            tanh_f := 1956;
        ELSIF x = 3864 THEN
            tanh_f := 1956;
        ELSIF x = 3865 THEN
            tanh_f := 1956;
        ELSIF x = 3866 THEN
            tanh_f := 1956;
        ELSIF x = 3867 THEN
            tanh_f := 1956;
        ELSIF x = 3868 THEN
            tanh_f := 1956;
        ELSIF x = 3869 THEN
            tanh_f := 1956;
        ELSIF x = 3870 THEN
            tanh_f := 1956;
        ELSIF x = 3871 THEN
            tanh_f := 1956;
        ELSIF x = 3872 THEN
            tanh_f := 1956;
        ELSIF x = 3873 THEN
            tanh_f := 1957;
        ELSIF x = 3874 THEN
            tanh_f := 1957;
        ELSIF x = 3875 THEN
            tanh_f := 1957;
        ELSIF x = 3876 THEN
            tanh_f := 1957;
        ELSIF x = 3877 THEN
            tanh_f := 1957;
        ELSIF x = 3878 THEN
            tanh_f := 1957;
        ELSIF x = 3879 THEN
            tanh_f := 1957;
        ELSIF x = 3880 THEN
            tanh_f := 1957;
        ELSIF x = 3881 THEN
            tanh_f := 1957;
        ELSIF x = 3882 THEN
            tanh_f := 1957;
        ELSIF x = 3883 THEN
            tanh_f := 1957;
        ELSIF x = 3884 THEN
            tanh_f := 1957;
        ELSIF x = 3885 THEN
            tanh_f := 1957;
        ELSIF x = 3886 THEN
            tanh_f := 1958;
        ELSIF x = 3887 THEN
            tanh_f := 1958;
        ELSIF x = 3888 THEN
            tanh_f := 1958;
        ELSIF x = 3889 THEN
            tanh_f := 1958;
        ELSIF x = 3890 THEN
            tanh_f := 1958;
        ELSIF x = 3891 THEN
            tanh_f := 1958;
        ELSIF x = 3892 THEN
            tanh_f := 1958;
        ELSIF x = 3893 THEN
            tanh_f := 1958;
        ELSIF x = 3894 THEN
            tanh_f := 1958;
        ELSIF x = 3895 THEN
            tanh_f := 1958;
        ELSIF x = 3896 THEN
            tanh_f := 1958;
        ELSIF x = 3897 THEN
            tanh_f := 1958;
        ELSIF x = 3898 THEN
            tanh_f := 1958;
        ELSIF x = 3899 THEN
            tanh_f := 1958;
        ELSIF x = 3900 THEN
            tanh_f := 1959;
        ELSIF x = 3901 THEN
            tanh_f := 1959;
        ELSIF x = 3902 THEN
            tanh_f := 1959;
        ELSIF x = 3903 THEN
            tanh_f := 1959;
        ELSIF x = 3904 THEN
            tanh_f := 1959;
        ELSIF x = 3905 THEN
            tanh_f := 1959;
        ELSIF x = 3906 THEN
            tanh_f := 1959;
        ELSIF x = 3907 THEN
            tanh_f := 1959;
        ELSIF x = 3908 THEN
            tanh_f := 1959;
        ELSIF x = 3909 THEN
            tanh_f := 1959;
        ELSIF x = 3910 THEN
            tanh_f := 1959;
        ELSIF x = 3911 THEN
            tanh_f := 1959;
        ELSIF x = 3912 THEN
            tanh_f := 1959;
        ELSIF x = 3913 THEN
            tanh_f := 1960;
        ELSIF x = 3914 THEN
            tanh_f := 1960;
        ELSIF x = 3915 THEN
            tanh_f := 1960;
        ELSIF x = 3916 THEN
            tanh_f := 1960;
        ELSIF x = 3917 THEN
            tanh_f := 1960;
        ELSIF x = 3918 THEN
            tanh_f := 1960;
        ELSIF x = 3919 THEN
            tanh_f := 1960;
        ELSIF x = 3920 THEN
            tanh_f := 1960;
        ELSIF x = 3921 THEN
            tanh_f := 1960;
        ELSIF x = 3922 THEN
            tanh_f := 1960;
        ELSIF x = 3923 THEN
            tanh_f := 1960;
        ELSIF x = 3924 THEN
            tanh_f := 1960;
        ELSIF x = 3925 THEN
            tanh_f := 1960;
        ELSIF x = 3926 THEN
            tanh_f := 1961;
        ELSIF x = 3927 THEN
            tanh_f := 1961;
        ELSIF x = 3928 THEN
            tanh_f := 1961;
        ELSIF x = 3929 THEN
            tanh_f := 1961;
        ELSIF x = 3930 THEN
            tanh_f := 1961;
        ELSIF x = 3931 THEN
            tanh_f := 1961;
        ELSIF x = 3932 THEN
            tanh_f := 1961;
        ELSIF x = 3933 THEN
            tanh_f := 1961;
        ELSIF x = 3934 THEN
            tanh_f := 1961;
        ELSIF x = 3935 THEN
            tanh_f := 1961;
        ELSIF x = 3936 THEN
            tanh_f := 1961;
        ELSIF x = 3937 THEN
            tanh_f := 1961;
        ELSIF x = 3938 THEN
            tanh_f := 1961;
        ELSIF x = 3939 THEN
            tanh_f := 1962;
        ELSIF x = 3940 THEN
            tanh_f := 1962;
        ELSIF x = 3941 THEN
            tanh_f := 1962;
        ELSIF x = 3942 THEN
            tanh_f := 1962;
        ELSIF x = 3943 THEN
            tanh_f := 1962;
        ELSIF x = 3944 THEN
            tanh_f := 1962;
        ELSIF x = 3945 THEN
            tanh_f := 1962;
        ELSIF x = 3946 THEN
            tanh_f := 1962;
        ELSIF x = 3947 THEN
            tanh_f := 1962;
        ELSIF x = 3948 THEN
            tanh_f := 1962;
        ELSIF x = 3949 THEN
            tanh_f := 1962;
        ELSIF x = 3950 THEN
            tanh_f := 1962;
        ELSIF x = 3951 THEN
            tanh_f := 1962;
        ELSIF x = 3952 THEN
            tanh_f := 1963;
        ELSIF x = 3953 THEN
            tanh_f := 1963;
        ELSIF x = 3954 THEN
            tanh_f := 1963;
        ELSIF x = 3955 THEN
            tanh_f := 1963;
        ELSIF x = 3956 THEN
            tanh_f := 1963;
        ELSIF x = 3957 THEN
            tanh_f := 1963;
        ELSIF x = 3958 THEN
            tanh_f := 1963;
        ELSIF x = 3959 THEN
            tanh_f := 1963;
        ELSIF x = 3960 THEN
            tanh_f := 1963;
        ELSIF x = 3961 THEN
            tanh_f := 1963;
        ELSIF x = 3962 THEN
            tanh_f := 1963;
        ELSIF x = 3963 THEN
            tanh_f := 1963;
        ELSIF x = 3964 THEN
            tanh_f := 1963;
        ELSIF x = 3965 THEN
            tanh_f := 1964;
        ELSIF x = 3966 THEN
            tanh_f := 1964;
        ELSIF x = 3967 THEN
            tanh_f := 1964;
        ELSIF x = 3968 THEN
            tanh_f := 1964;
        ELSIF x = 3969 THEN
            tanh_f := 1964;
        ELSIF x = 3970 THEN
            tanh_f := 1964;
        ELSIF x = 3971 THEN
            tanh_f := 1964;
        ELSIF x = 3972 THEN
            tanh_f := 1964;
        ELSIF x = 3973 THEN
            tanh_f := 1964;
        ELSIF x = 3974 THEN
            tanh_f := 1964;
        ELSIF x = 3975 THEN
            tanh_f := 1964;
        ELSIF x = 3976 THEN
            tanh_f := 1964;
        ELSIF x = 3977 THEN
            tanh_f := 1964;
        ELSIF x = 3978 THEN
            tanh_f := 1965;
        ELSIF x = 3979 THEN
            tanh_f := 1965;
        ELSIF x = 3980 THEN
            tanh_f := 1965;
        ELSIF x = 3981 THEN
            tanh_f := 1965;
        ELSIF x = 3982 THEN
            tanh_f := 1965;
        ELSIF x = 3983 THEN
            tanh_f := 1965;
        ELSIF x = 3984 THEN
            tanh_f := 1965;
        ELSIF x = 3985 THEN
            tanh_f := 1965;
        ELSIF x = 3986 THEN
            tanh_f := 1965;
        ELSIF x = 3987 THEN
            tanh_f := 1965;
        ELSIF x = 3988 THEN
            tanh_f := 1965;
        ELSIF x = 3989 THEN
            tanh_f := 1965;
        ELSIF x = 3990 THEN
            tanh_f := 1965;
        ELSIF x = 3991 THEN
            tanh_f := 1966;
        ELSIF x = 3992 THEN
            tanh_f := 1966;
        ELSIF x = 3993 THEN
            tanh_f := 1966;
        ELSIF x = 3994 THEN
            tanh_f := 1966;
        ELSIF x = 3995 THEN
            tanh_f := 1966;
        ELSIF x = 3996 THEN
            tanh_f := 1966;
        ELSIF x = 3997 THEN
            tanh_f := 1966;
        ELSIF x = 3998 THEN
            tanh_f := 1966;
        ELSIF x = 3999 THEN
            tanh_f := 1966;
        ELSIF x = 4000 THEN
            tanh_f := 1966;
        ELSIF x = 4001 THEN
            tanh_f := 1966;
        ELSIF x = 4002 THEN
            tanh_f := 1966;
        ELSIF x = 4003 THEN
            tanh_f := 1966;
        ELSIF x = 4004 THEN
            tanh_f := 1966;
        ELSIF x = 4005 THEN
            tanh_f := 1967;
        ELSIF x = 4006 THEN
            tanh_f := 1967;
        ELSIF x = 4007 THEN
            tanh_f := 1967;
        ELSIF x = 4008 THEN
            tanh_f := 1967;
        ELSIF x = 4009 THEN
            tanh_f := 1967;
        ELSIF x = 4010 THEN
            tanh_f := 1967;
        ELSIF x = 4011 THEN
            tanh_f := 1967;
        ELSIF x = 4012 THEN
            tanh_f := 1967;
        ELSIF x = 4013 THEN
            tanh_f := 1967;
        ELSIF x = 4014 THEN
            tanh_f := 1967;
        ELSIF x = 4015 THEN
            tanh_f := 1967;
        ELSIF x = 4016 THEN
            tanh_f := 1967;
        ELSIF x = 4017 THEN
            tanh_f := 1967;
        ELSIF x = 4018 THEN
            tanh_f := 1968;
        ELSIF x = 4019 THEN
            tanh_f := 1968;
        ELSIF x = 4020 THEN
            tanh_f := 1968;
        ELSIF x = 4021 THEN
            tanh_f := 1968;
        ELSIF x = 4022 THEN
            tanh_f := 1968;
        ELSIF x = 4023 THEN
            tanh_f := 1968;
        ELSIF x = 4024 THEN
            tanh_f := 1968;
        ELSIF x = 4025 THEN
            tanh_f := 1968;
        ELSIF x = 4026 THEN
            tanh_f := 1968;
        ELSIF x = 4027 THEN
            tanh_f := 1968;
        ELSIF x = 4028 THEN
            tanh_f := 1968;
        ELSIF x = 4029 THEN
            tanh_f := 1968;
        ELSIF x = 4030 THEN
            tanh_f := 1968;
        ELSIF x = 4031 THEN
            tanh_f := 1969;
        ELSIF x = 4032 THEN
            tanh_f := 1969;
        ELSIF x = 4033 THEN
            tanh_f := 1969;
        ELSIF x = 4034 THEN
            tanh_f := 1969;
        ELSIF x = 4035 THEN
            tanh_f := 1969;
        ELSIF x = 4036 THEN
            tanh_f := 1969;
        ELSIF x = 4037 THEN
            tanh_f := 1969;
        ELSIF x = 4038 THEN
            tanh_f := 1969;
        ELSIF x = 4039 THEN
            tanh_f := 1969;
        ELSIF x = 4040 THEN
            tanh_f := 1969;
        ELSIF x = 4041 THEN
            tanh_f := 1969;
        ELSIF x = 4042 THEN
            tanh_f := 1969;
        ELSIF x = 4043 THEN
            tanh_f := 1969;
        ELSIF x = 4044 THEN
            tanh_f := 1970;
        ELSIF x = 4045 THEN
            tanh_f := 1970;
        ELSIF x = 4046 THEN
            tanh_f := 1970;
        ELSIF x = 4047 THEN
            tanh_f := 1970;
        ELSIF x = 4048 THEN
            tanh_f := 1970;
        ELSIF x = 4049 THEN
            tanh_f := 1970;
        ELSIF x = 4050 THEN
            tanh_f := 1970;
        ELSIF x = 4051 THEN
            tanh_f := 1970;
        ELSIF x = 4052 THEN
            tanh_f := 1970;
        ELSIF x = 4053 THEN
            tanh_f := 1970;
        ELSIF x = 4054 THEN
            tanh_f := 1970;
        ELSIF x = 4055 THEN
            tanh_f := 1970;
        ELSIF x = 4056 THEN
            tanh_f := 1970;
        ELSIF x = 4057 THEN
            tanh_f := 1971;
        ELSIF x = 4058 THEN
            tanh_f := 1971;
        ELSIF x = 4059 THEN
            tanh_f := 1971;
        ELSIF x = 4060 THEN
            tanh_f := 1971;
        ELSIF x = 4061 THEN
            tanh_f := 1971;
        ELSIF x = 4062 THEN
            tanh_f := 1971;
        ELSIF x = 4063 THEN
            tanh_f := 1971;
        ELSIF x = 4064 THEN
            tanh_f := 1971;
        ELSIF x = 4065 THEN
            tanh_f := 1971;
        ELSIF x = 4066 THEN
            tanh_f := 1971;
        ELSIF x = 4067 THEN
            tanh_f := 1971;
        ELSIF x = 4068 THEN
            tanh_f := 1971;
        ELSIF x = 4069 THEN
            tanh_f := 1971;
        ELSIF x = 4070 THEN
            tanh_f := 1972;
        ELSIF x = 4071 THEN
            tanh_f := 1972;
        ELSIF x = 4072 THEN
            tanh_f := 1972;
        ELSIF x = 4073 THEN
            tanh_f := 1972;
        ELSIF x = 4074 THEN
            tanh_f := 1972;
        ELSIF x = 4075 THEN
            tanh_f := 1972;
        ELSIF x = 4076 THEN
            tanh_f := 1972;
        ELSIF x = 4077 THEN
            tanh_f := 1972;
        ELSIF x = 4078 THEN
            tanh_f := 1972;
        ELSIF x = 4079 THEN
            tanh_f := 1972;
        ELSIF x = 4080 THEN
            tanh_f := 1972;
        ELSIF x = 4081 THEN
            tanh_f := 1972;
        ELSIF x = 4082 THEN
            tanh_f := 1972;
        ELSIF x = 4083 THEN
            tanh_f := 1973;
        ELSIF x = 4084 THEN
            tanh_f := 1973;
        ELSIF x = 4085 THEN
            tanh_f := 1973;
        ELSIF x = 4086 THEN
            tanh_f := 1973;
        ELSIF x = 4087 THEN
            tanh_f := 1973;
        ELSIF x = 4088 THEN
            tanh_f := 1973;
        ELSIF x = 4089 THEN
            tanh_f := 1973;
        ELSIF x = 4090 THEN
            tanh_f := 1973;
        ELSIF x = 4091 THEN
            tanh_f := 1973;
        ELSIF x = 4092 THEN
            tanh_f := 1973;
        ELSIF x = 4093 THEN
            tanh_f := 1973;
        ELSIF x = 4094 THEN
            tanh_f := 1973;
        ELSIF x = 4095 THEN
            tanh_f := 1973;
        ELSIF x = 4096 THEN
            tanh_f := 1974;
        ELSIF x = 4097 THEN
            tanh_f := 1974;
        ELSIF x = 4098 THEN
            tanh_f := 1974;
        ELSIF x = 4099 THEN
            tanh_f := 1974;
        ELSIF x = 4100 THEN
            tanh_f := 1974;
        ELSIF x = 4101 THEN
            tanh_f := 1974;
        ELSIF x = 4102 THEN
            tanh_f := 1974;
        ELSIF x = 4103 THEN
            tanh_f := 1974;
        ELSIF x = 4104 THEN
            tanh_f := 1974;
        ELSIF x = 4105 THEN
            tanh_f := 1974;
        ELSIF x = 4106 THEN
            tanh_f := 1974;
        ELSIF x = 4107 THEN
            tanh_f := 1974;
        ELSIF x = 4108 THEN
            tanh_f := 1974;
        ELSIF x = 4109 THEN
            tanh_f := 1974;
        ELSIF x = 4110 THEN
            tanh_f := 1974;
        ELSIF x = 4111 THEN
            tanh_f := 1974;
        ELSIF x = 4112 THEN
            tanh_f := 1975;
        ELSIF x = 4113 THEN
            tanh_f := 1975;
        ELSIF x = 4114 THEN
            tanh_f := 1975;
        ELSIF x = 4115 THEN
            tanh_f := 1975;
        ELSIF x = 4116 THEN
            tanh_f := 1975;
        ELSIF x = 4117 THEN
            tanh_f := 1975;
        ELSIF x = 4118 THEN
            tanh_f := 1975;
        ELSIF x = 4119 THEN
            tanh_f := 1975;
        ELSIF x = 4120 THEN
            tanh_f := 1975;
        ELSIF x = 4121 THEN
            tanh_f := 1975;
        ELSIF x = 4122 THEN
            tanh_f := 1975;
        ELSIF x = 4123 THEN
            tanh_f := 1975;
        ELSIF x = 4124 THEN
            tanh_f := 1975;
        ELSIF x = 4125 THEN
            tanh_f := 1975;
        ELSIF x = 4126 THEN
            tanh_f := 1975;
        ELSIF x = 4127 THEN
            tanh_f := 1976;
        ELSIF x = 4128 THEN
            tanh_f := 1976;
        ELSIF x = 4129 THEN
            tanh_f := 1976;
        ELSIF x = 4130 THEN
            tanh_f := 1976;
        ELSIF x = 4131 THEN
            tanh_f := 1976;
        ELSIF x = 4132 THEN
            tanh_f := 1976;
        ELSIF x = 4133 THEN
            tanh_f := 1976;
        ELSIF x = 4134 THEN
            tanh_f := 1976;
        ELSIF x = 4135 THEN
            tanh_f := 1976;
        ELSIF x = 4136 THEN
            tanh_f := 1976;
        ELSIF x = 4137 THEN
            tanh_f := 1976;
        ELSIF x = 4138 THEN
            tanh_f := 1976;
        ELSIF x = 4139 THEN
            tanh_f := 1976;
        ELSIF x = 4140 THEN
            tanh_f := 1976;
        ELSIF x = 4141 THEN
            tanh_f := 1976;
        ELSIF x = 4142 THEN
            tanh_f := 1977;
        ELSIF x = 4143 THEN
            tanh_f := 1977;
        ELSIF x = 4144 THEN
            tanh_f := 1977;
        ELSIF x = 4145 THEN
            tanh_f := 1977;
        ELSIF x = 4146 THEN
            tanh_f := 1977;
        ELSIF x = 4147 THEN
            tanh_f := 1977;
        ELSIF x = 4148 THEN
            tanh_f := 1977;
        ELSIF x = 4149 THEN
            tanh_f := 1977;
        ELSIF x = 4150 THEN
            tanh_f := 1977;
        ELSIF x = 4151 THEN
            tanh_f := 1977;
        ELSIF x = 4152 THEN
            tanh_f := 1977;
        ELSIF x = 4153 THEN
            tanh_f := 1977;
        ELSIF x = 4154 THEN
            tanh_f := 1977;
        ELSIF x = 4155 THEN
            tanh_f := 1977;
        ELSIF x = 4156 THEN
            tanh_f := 1977;
        ELSIF x = 4157 THEN
            tanh_f := 1978;
        ELSIF x = 4158 THEN
            tanh_f := 1978;
        ELSIF x = 4159 THEN
            tanh_f := 1978;
        ELSIF x = 4160 THEN
            tanh_f := 1978;
        ELSIF x = 4161 THEN
            tanh_f := 1978;
        ELSIF x = 4162 THEN
            tanh_f := 1978;
        ELSIF x = 4163 THEN
            tanh_f := 1978;
        ELSIF x = 4164 THEN
            tanh_f := 1978;
        ELSIF x = 4165 THEN
            tanh_f := 1978;
        ELSIF x = 4166 THEN
            tanh_f := 1978;
        ELSIF x = 4167 THEN
            tanh_f := 1978;
        ELSIF x = 4168 THEN
            tanh_f := 1978;
        ELSIF x = 4169 THEN
            tanh_f := 1978;
        ELSIF x = 4170 THEN
            tanh_f := 1978;
        ELSIF x = 4171 THEN
            tanh_f := 1978;
        ELSIF x = 4172 THEN
            tanh_f := 1979;
        ELSIF x = 4173 THEN
            tanh_f := 1979;
        ELSIF x = 4174 THEN
            tanh_f := 1979;
        ELSIF x = 4175 THEN
            tanh_f := 1979;
        ELSIF x = 4176 THEN
            tanh_f := 1979;
        ELSIF x = 4177 THEN
            tanh_f := 1979;
        ELSIF x = 4178 THEN
            tanh_f := 1979;
        ELSIF x = 4179 THEN
            tanh_f := 1979;
        ELSIF x = 4180 THEN
            tanh_f := 1979;
        ELSIF x = 4181 THEN
            tanh_f := 1979;
        ELSIF x = 4182 THEN
            tanh_f := 1979;
        ELSIF x = 4183 THEN
            tanh_f := 1979;
        ELSIF x = 4184 THEN
            tanh_f := 1979;
        ELSIF x = 4185 THEN
            tanh_f := 1979;
        ELSIF x = 4186 THEN
            tanh_f := 1979;
        ELSIF x = 4187 THEN
            tanh_f := 1980;
        ELSIF x = 4188 THEN
            tanh_f := 1980;
        ELSIF x = 4189 THEN
            tanh_f := 1980;
        ELSIF x = 4190 THEN
            tanh_f := 1980;
        ELSIF x = 4191 THEN
            tanh_f := 1980;
        ELSIF x = 4192 THEN
            tanh_f := 1980;
        ELSIF x = 4193 THEN
            tanh_f := 1980;
        ELSIF x = 4194 THEN
            tanh_f := 1980;
        ELSIF x = 4195 THEN
            tanh_f := 1980;
        ELSIF x = 4196 THEN
            tanh_f := 1980;
        ELSIF x = 4197 THEN
            tanh_f := 1980;
        ELSIF x = 4198 THEN
            tanh_f := 1980;
        ELSIF x = 4199 THEN
            tanh_f := 1980;
        ELSIF x = 4200 THEN
            tanh_f := 1980;
        ELSIF x = 4201 THEN
            tanh_f := 1980;
        ELSIF x = 4202 THEN
            tanh_f := 1981;
        ELSIF x = 4203 THEN
            tanh_f := 1981;
        ELSIF x = 4204 THEN
            tanh_f := 1981;
        ELSIF x = 4205 THEN
            tanh_f := 1981;
        ELSIF x = 4206 THEN
            tanh_f := 1981;
        ELSIF x = 4207 THEN
            tanh_f := 1981;
        ELSIF x = 4208 THEN
            tanh_f := 1981;
        ELSIF x = 4209 THEN
            tanh_f := 1981;
        ELSIF x = 4210 THEN
            tanh_f := 1981;
        ELSIF x = 4211 THEN
            tanh_f := 1981;
        ELSIF x = 4212 THEN
            tanh_f := 1981;
        ELSIF x = 4213 THEN
            tanh_f := 1981;
        ELSIF x = 4214 THEN
            tanh_f := 1981;
        ELSIF x = 4215 THEN
            tanh_f := 1981;
        ELSIF x = 4216 THEN
            tanh_f := 1981;
        ELSIF x = 4217 THEN
            tanh_f := 1982;
        ELSIF x = 4218 THEN
            tanh_f := 1982;
        ELSIF x = 4219 THEN
            tanh_f := 1982;
        ELSIF x = 4220 THEN
            tanh_f := 1982;
        ELSIF x = 4221 THEN
            tanh_f := 1982;
        ELSIF x = 4222 THEN
            tanh_f := 1982;
        ELSIF x = 4223 THEN
            tanh_f := 1982;
        ELSIF x = 4224 THEN
            tanh_f := 1982;
        ELSIF x = 4225 THEN
            tanh_f := 1982;
        ELSIF x = 4226 THEN
            tanh_f := 1982;
        ELSIF x = 4227 THEN
            tanh_f := 1982;
        ELSIF x = 4228 THEN
            tanh_f := 1982;
        ELSIF x = 4229 THEN
            tanh_f := 1982;
        ELSIF x = 4230 THEN
            tanh_f := 1982;
        ELSIF x = 4231 THEN
            tanh_f := 1982;
        ELSIF x = 4232 THEN
            tanh_f := 1983;
        ELSIF x = 4233 THEN
            tanh_f := 1983;
        ELSIF x = 4234 THEN
            tanh_f := 1983;
        ELSIF x = 4235 THEN
            tanh_f := 1983;
        ELSIF x = 4236 THEN
            tanh_f := 1983;
        ELSIF x = 4237 THEN
            tanh_f := 1983;
        ELSIF x = 4238 THEN
            tanh_f := 1983;
        ELSIF x = 4239 THEN
            tanh_f := 1983;
        ELSIF x = 4240 THEN
            tanh_f := 1983;
        ELSIF x = 4241 THEN
            tanh_f := 1983;
        ELSIF x = 4242 THEN
            tanh_f := 1983;
        ELSIF x = 4243 THEN
            tanh_f := 1983;
        ELSIF x = 4244 THEN
            tanh_f := 1983;
        ELSIF x = 4245 THEN
            tanh_f := 1983;
        ELSIF x = 4246 THEN
            tanh_f := 1983;
        ELSIF x = 4247 THEN
            tanh_f := 1984;
        ELSIF x = 4248 THEN
            tanh_f := 1984;
        ELSIF x = 4249 THEN
            tanh_f := 1984;
        ELSIF x = 4250 THEN
            tanh_f := 1984;
        ELSIF x = 4251 THEN
            tanh_f := 1984;
        ELSIF x = 4252 THEN
            tanh_f := 1984;
        ELSIF x = 4253 THEN
            tanh_f := 1984;
        ELSIF x = 4254 THEN
            tanh_f := 1984;
        ELSIF x = 4255 THEN
            tanh_f := 1984;
        ELSIF x = 4256 THEN
            tanh_f := 1984;
        ELSIF x = 4257 THEN
            tanh_f := 1984;
        ELSIF x = 4258 THEN
            tanh_f := 1984;
        ELSIF x = 4259 THEN
            tanh_f := 1984;
        ELSIF x = 4260 THEN
            tanh_f := 1984;
        ELSIF x = 4261 THEN
            tanh_f := 1984;
        ELSIF x = 4262 THEN
            tanh_f := 1985;
        ELSIF x = 4263 THEN
            tanh_f := 1985;
        ELSIF x = 4264 THEN
            tanh_f := 1985;
        ELSIF x = 4265 THEN
            tanh_f := 1985;
        ELSIF x = 4266 THEN
            tanh_f := 1985;
        ELSIF x = 4267 THEN
            tanh_f := 1985;
        ELSIF x = 4268 THEN
            tanh_f := 1985;
        ELSIF x = 4269 THEN
            tanh_f := 1985;
        ELSIF x = 4270 THEN
            tanh_f := 1985;
        ELSIF x = 4271 THEN
            tanh_f := 1985;
        ELSIF x = 4272 THEN
            tanh_f := 1985;
        ELSIF x = 4273 THEN
            tanh_f := 1985;
        ELSIF x = 4274 THEN
            tanh_f := 1985;
        ELSIF x = 4275 THEN
            tanh_f := 1985;
        ELSIF x = 4276 THEN
            tanh_f := 1985;
        ELSIF x = 4277 THEN
            tanh_f := 1986;
        ELSIF x = 4278 THEN
            tanh_f := 1986;
        ELSIF x = 4279 THEN
            tanh_f := 1986;
        ELSIF x = 4280 THEN
            tanh_f := 1986;
        ELSIF x = 4281 THEN
            tanh_f := 1986;
        ELSIF x = 4282 THEN
            tanh_f := 1986;
        ELSIF x = 4283 THEN
            tanh_f := 1986;
        ELSIF x = 4284 THEN
            tanh_f := 1986;
        ELSIF x = 4285 THEN
            tanh_f := 1986;
        ELSIF x = 4286 THEN
            tanh_f := 1986;
        ELSIF x = 4287 THEN
            tanh_f := 1986;
        ELSIF x = 4288 THEN
            tanh_f := 1986;
        ELSIF x = 4289 THEN
            tanh_f := 1986;
        ELSIF x = 4290 THEN
            tanh_f := 1986;
        ELSIF x = 4291 THEN
            tanh_f := 1986;
        ELSIF x = 4292 THEN
            tanh_f := 1987;
        ELSIF x = 4293 THEN
            tanh_f := 1987;
        ELSIF x = 4294 THEN
            tanh_f := 1987;
        ELSIF x = 4295 THEN
            tanh_f := 1987;
        ELSIF x = 4296 THEN
            tanh_f := 1987;
        ELSIF x = 4297 THEN
            tanh_f := 1987;
        ELSIF x = 4298 THEN
            tanh_f := 1987;
        ELSIF x = 4299 THEN
            tanh_f := 1987;
        ELSIF x = 4300 THEN
            tanh_f := 1987;
        ELSIF x = 4301 THEN
            tanh_f := 1987;
        ELSIF x = 4302 THEN
            tanh_f := 1987;
        ELSIF x = 4303 THEN
            tanh_f := 1987;
        ELSIF x = 4304 THEN
            tanh_f := 1987;
        ELSIF x = 4305 THEN
            tanh_f := 1987;
        ELSIF x = 4306 THEN
            tanh_f := 1987;
        ELSIF x = 4307 THEN
            tanh_f := 1988;
        ELSIF x = 4308 THEN
            tanh_f := 1988;
        ELSIF x = 4309 THEN
            tanh_f := 1988;
        ELSIF x = 4310 THEN
            tanh_f := 1988;
        ELSIF x = 4311 THEN
            tanh_f := 1988;
        ELSIF x = 4312 THEN
            tanh_f := 1988;
        ELSIF x = 4313 THEN
            tanh_f := 1988;
        ELSIF x = 4314 THEN
            tanh_f := 1988;
        ELSIF x = 4315 THEN
            tanh_f := 1988;
        ELSIF x = 4316 THEN
            tanh_f := 1988;
        ELSIF x = 4317 THEN
            tanh_f := 1988;
        ELSIF x = 4318 THEN
            tanh_f := 1988;
        ELSIF x = 4319 THEN
            tanh_f := 1988;
        ELSIF x = 4320 THEN
            tanh_f := 1988;
        ELSIF x = 4321 THEN
            tanh_f := 1988;
        ELSIF x = 4322 THEN
            tanh_f := 1989;
        ELSIF x = 4323 THEN
            tanh_f := 1989;
        ELSIF x = 4324 THEN
            tanh_f := 1989;
        ELSIF x = 4325 THEN
            tanh_f := 1989;
        ELSIF x = 4326 THEN
            tanh_f := 1989;
        ELSIF x = 4327 THEN
            tanh_f := 1989;
        ELSIF x = 4328 THEN
            tanh_f := 1989;
        ELSIF x = 4329 THEN
            tanh_f := 1989;
        ELSIF x = 4330 THEN
            tanh_f := 1989;
        ELSIF x = 4331 THEN
            tanh_f := 1989;
        ELSIF x = 4332 THEN
            tanh_f := 1989;
        ELSIF x = 4333 THEN
            tanh_f := 1989;
        ELSIF x = 4334 THEN
            tanh_f := 1989;
        ELSIF x = 4335 THEN
            tanh_f := 1989;
        ELSIF x = 4336 THEN
            tanh_f := 1989;
        ELSIF x = 4337 THEN
            tanh_f := 1990;
        ELSIF x = 4338 THEN
            tanh_f := 1990;
        ELSIF x = 4339 THEN
            tanh_f := 1990;
        ELSIF x = 4340 THEN
            tanh_f := 1990;
        ELSIF x = 4341 THEN
            tanh_f := 1990;
        ELSIF x = 4342 THEN
            tanh_f := 1990;
        ELSIF x = 4343 THEN
            tanh_f := 1990;
        ELSIF x = 4344 THEN
            tanh_f := 1990;
        ELSIF x = 4345 THEN
            tanh_f := 1990;
        ELSIF x = 4346 THEN
            tanh_f := 1990;
        ELSIF x = 4347 THEN
            tanh_f := 1990;
        ELSIF x = 4348 THEN
            tanh_f := 1990;
        ELSIF x = 4349 THEN
            tanh_f := 1990;
        ELSIF x = 4350 THEN
            tanh_f := 1990;
        ELSIF x = 4351 THEN
            tanh_f := 1990;
        ELSIF x = 4352 THEN
            tanh_f := 1990;
        ELSIF x = 4353 THEN
            tanh_f := 1990;
        ELSIF x = 4354 THEN
            tanh_f := 1990;
        ELSIF x = 4355 THEN
            tanh_f := 1990;
        ELSIF x = 4356 THEN
            tanh_f := 1990;
        ELSIF x = 4357 THEN
            tanh_f := 1990;
        ELSIF x = 4358 THEN
            tanh_f := 1990;
        ELSIF x = 4359 THEN
            tanh_f := 1990;
        ELSIF x = 4360 THEN
            tanh_f := 1990;
        ELSIF x = 4361 THEN
            tanh_f := 1990;
        ELSIF x = 4362 THEN
            tanh_f := 1990;
        ELSIF x = 4363 THEN
            tanh_f := 1991;
        ELSIF x = 4364 THEN
            tanh_f := 1991;
        ELSIF x = 4365 THEN
            tanh_f := 1991;
        ELSIF x = 4366 THEN
            tanh_f := 1991;
        ELSIF x = 4367 THEN
            tanh_f := 1991;
        ELSIF x = 4368 THEN
            tanh_f := 1991;
        ELSIF x = 4369 THEN
            tanh_f := 1991;
        ELSIF x = 4370 THEN
            tanh_f := 1991;
        ELSIF x = 4371 THEN
            tanh_f := 1991;
        ELSIF x = 4372 THEN
            tanh_f := 1991;
        ELSIF x = 4373 THEN
            tanh_f := 1991;
        ELSIF x = 4374 THEN
            tanh_f := 1991;
        ELSIF x = 4375 THEN
            tanh_f := 1991;
        ELSIF x = 4376 THEN
            tanh_f := 1991;
        ELSIF x = 4377 THEN
            tanh_f := 1991;
        ELSIF x = 4378 THEN
            tanh_f := 1991;
        ELSIF x = 4379 THEN
            tanh_f := 1991;
        ELSIF x = 4380 THEN
            tanh_f := 1991;
        ELSIF x = 4381 THEN
            tanh_f := 1991;
        ELSIF x = 4382 THEN
            tanh_f := 1991;
        ELSIF x = 4383 THEN
            tanh_f := 1992;
        ELSIF x = 4384 THEN
            tanh_f := 1992;
        ELSIF x = 4385 THEN
            tanh_f := 1992;
        ELSIF x = 4386 THEN
            tanh_f := 1992;
        ELSIF x = 4387 THEN
            tanh_f := 1992;
        ELSIF x = 4388 THEN
            tanh_f := 1992;
        ELSIF x = 4389 THEN
            tanh_f := 1992;
        ELSIF x = 4390 THEN
            tanh_f := 1992;
        ELSIF x = 4391 THEN
            tanh_f := 1992;
        ELSIF x = 4392 THEN
            tanh_f := 1992;
        ELSIF x = 4393 THEN
            tanh_f := 1992;
        ELSIF x = 4394 THEN
            tanh_f := 1992;
        ELSIF x = 4395 THEN
            tanh_f := 1992;
        ELSIF x = 4396 THEN
            tanh_f := 1992;
        ELSIF x = 4397 THEN
            tanh_f := 1992;
        ELSIF x = 4398 THEN
            tanh_f := 1992;
        ELSIF x = 4399 THEN
            tanh_f := 1992;
        ELSIF x = 4400 THEN
            tanh_f := 1992;
        ELSIF x = 4401 THEN
            tanh_f := 1992;
        ELSIF x = 4402 THEN
            tanh_f := 1992;
        ELSIF x = 4403 THEN
            tanh_f := 1992;
        ELSIF x = 4404 THEN
            tanh_f := 1993;
        ELSIF x = 4405 THEN
            tanh_f := 1993;
        ELSIF x = 4406 THEN
            tanh_f := 1993;
        ELSIF x = 4407 THEN
            tanh_f := 1993;
        ELSIF x = 4408 THEN
            tanh_f := 1993;
        ELSIF x = 4409 THEN
            tanh_f := 1993;
        ELSIF x = 4410 THEN
            tanh_f := 1993;
        ELSIF x = 4411 THEN
            tanh_f := 1993;
        ELSIF x = 4412 THEN
            tanh_f := 1993;
        ELSIF x = 4413 THEN
            tanh_f := 1993;
        ELSIF x = 4414 THEN
            tanh_f := 1993;
        ELSIF x = 4415 THEN
            tanh_f := 1993;
        ELSIF x = 4416 THEN
            tanh_f := 1993;
        ELSIF x = 4417 THEN
            tanh_f := 1993;
        ELSIF x = 4418 THEN
            tanh_f := 1993;
        ELSIF x = 4419 THEN
            tanh_f := 1993;
        ELSIF x = 4420 THEN
            tanh_f := 1993;
        ELSIF x = 4421 THEN
            tanh_f := 1993;
        ELSIF x = 4422 THEN
            tanh_f := 1993;
        ELSIF x = 4423 THEN
            tanh_f := 1993;
        ELSIF x = 4424 THEN
            tanh_f := 1994;
        ELSIF x = 4425 THEN
            tanh_f := 1994;
        ELSIF x = 4426 THEN
            tanh_f := 1994;
        ELSIF x = 4427 THEN
            tanh_f := 1994;
        ELSIF x = 4428 THEN
            tanh_f := 1994;
        ELSIF x = 4429 THEN
            tanh_f := 1994;
        ELSIF x = 4430 THEN
            tanh_f := 1994;
        ELSIF x = 4431 THEN
            tanh_f := 1994;
        ELSIF x = 4432 THEN
            tanh_f := 1994;
        ELSIF x = 4433 THEN
            tanh_f := 1994;
        ELSIF x = 4434 THEN
            tanh_f := 1994;
        ELSIF x = 4435 THEN
            tanh_f := 1994;
        ELSIF x = 4436 THEN
            tanh_f := 1994;
        ELSIF x = 4437 THEN
            tanh_f := 1994;
        ELSIF x = 4438 THEN
            tanh_f := 1994;
        ELSIF x = 4439 THEN
            tanh_f := 1994;
        ELSIF x = 4440 THEN
            tanh_f := 1994;
        ELSIF x = 4441 THEN
            tanh_f := 1994;
        ELSIF x = 4442 THEN
            tanh_f := 1994;
        ELSIF x = 4443 THEN
            tanh_f := 1994;
        ELSIF x = 4444 THEN
            tanh_f := 1994;
        ELSIF x = 4445 THEN
            tanh_f := 1995;
        ELSIF x = 4446 THEN
            tanh_f := 1995;
        ELSIF x = 4447 THEN
            tanh_f := 1995;
        ELSIF x = 4448 THEN
            tanh_f := 1995;
        ELSIF x = 4449 THEN
            tanh_f := 1995;
        ELSIF x = 4450 THEN
            tanh_f := 1995;
        ELSIF x = 4451 THEN
            tanh_f := 1995;
        ELSIF x = 4452 THEN
            tanh_f := 1995;
        ELSIF x = 4453 THEN
            tanh_f := 1995;
        ELSIF x = 4454 THEN
            tanh_f := 1995;
        ELSIF x = 4455 THEN
            tanh_f := 1995;
        ELSIF x = 4456 THEN
            tanh_f := 1995;
        ELSIF x = 4457 THEN
            tanh_f := 1995;
        ELSIF x = 4458 THEN
            tanh_f := 1995;
        ELSIF x = 4459 THEN
            tanh_f := 1995;
        ELSIF x = 4460 THEN
            tanh_f := 1995;
        ELSIF x = 4461 THEN
            tanh_f := 1995;
        ELSIF x = 4462 THEN
            tanh_f := 1995;
        ELSIF x = 4463 THEN
            tanh_f := 1995;
        ELSIF x = 4464 THEN
            tanh_f := 1995;
        ELSIF x = 4465 THEN
            tanh_f := 1996;
        ELSIF x = 4466 THEN
            tanh_f := 1996;
        ELSIF x = 4467 THEN
            tanh_f := 1996;
        ELSIF x = 4468 THEN
            tanh_f := 1996;
        ELSIF x = 4469 THEN
            tanh_f := 1996;
        ELSIF x = 4470 THEN
            tanh_f := 1996;
        ELSIF x = 4471 THEN
            tanh_f := 1996;
        ELSIF x = 4472 THEN
            tanh_f := 1996;
        ELSIF x = 4473 THEN
            tanh_f := 1996;
        ELSIF x = 4474 THEN
            tanh_f := 1996;
        ELSIF x = 4475 THEN
            tanh_f := 1996;
        ELSIF x = 4476 THEN
            tanh_f := 1996;
        ELSIF x = 4477 THEN
            tanh_f := 1996;
        ELSIF x = 4478 THEN
            tanh_f := 1996;
        ELSIF x = 4479 THEN
            tanh_f := 1996;
        ELSIF x = 4480 THEN
            tanh_f := 1996;
        ELSIF x = 4481 THEN
            tanh_f := 1996;
        ELSIF x = 4482 THEN
            tanh_f := 1996;
        ELSIF x = 4483 THEN
            tanh_f := 1996;
        ELSIF x = 4484 THEN
            tanh_f := 1996;
        ELSIF x = 4485 THEN
            tanh_f := 1996;
        ELSIF x = 4486 THEN
            tanh_f := 1997;
        ELSIF x = 4487 THEN
            tanh_f := 1997;
        ELSIF x = 4488 THEN
            tanh_f := 1997;
        ELSIF x = 4489 THEN
            tanh_f := 1997;
        ELSIF x = 4490 THEN
            tanh_f := 1997;
        ELSIF x = 4491 THEN
            tanh_f := 1997;
        ELSIF x = 4492 THEN
            tanh_f := 1997;
        ELSIF x = 4493 THEN
            tanh_f := 1997;
        ELSIF x = 4494 THEN
            tanh_f := 1997;
        ELSIF x = 4495 THEN
            tanh_f := 1997;
        ELSIF x = 4496 THEN
            tanh_f := 1997;
        ELSIF x = 4497 THEN
            tanh_f := 1997;
        ELSIF x = 4498 THEN
            tanh_f := 1997;
        ELSIF x = 4499 THEN
            tanh_f := 1997;
        ELSIF x = 4500 THEN
            tanh_f := 1997;
        ELSIF x = 4501 THEN
            tanh_f := 1997;
        ELSIF x = 4502 THEN
            tanh_f := 1997;
        ELSIF x = 4503 THEN
            tanh_f := 1997;
        ELSIF x = 4504 THEN
            tanh_f := 1997;
        ELSIF x = 4505 THEN
            tanh_f := 1997;
        ELSIF x = 4506 THEN
            tanh_f := 1998;
        ELSIF x = 4507 THEN
            tanh_f := 1998;
        ELSIF x = 4508 THEN
            tanh_f := 1998;
        ELSIF x = 4509 THEN
            tanh_f := 1998;
        ELSIF x = 4510 THEN
            tanh_f := 1998;
        ELSIF x = 4511 THEN
            tanh_f := 1998;
        ELSIF x = 4512 THEN
            tanh_f := 1998;
        ELSIF x = 4513 THEN
            tanh_f := 1998;
        ELSIF x = 4514 THEN
            tanh_f := 1998;
        ELSIF x = 4515 THEN
            tanh_f := 1998;
        ELSIF x = 4516 THEN
            tanh_f := 1998;
        ELSIF x = 4517 THEN
            tanh_f := 1998;
        ELSIF x = 4518 THEN
            tanh_f := 1998;
        ELSIF x = 4519 THEN
            tanh_f := 1998;
        ELSIF x = 4520 THEN
            tanh_f := 1998;
        ELSIF x = 4521 THEN
            tanh_f := 1998;
        ELSIF x = 4522 THEN
            tanh_f := 1998;
        ELSIF x = 4523 THEN
            tanh_f := 1998;
        ELSIF x = 4524 THEN
            tanh_f := 1998;
        ELSIF x = 4525 THEN
            tanh_f := 1998;
        ELSIF x = 4526 THEN
            tanh_f := 1998;
        ELSIF x = 4527 THEN
            tanh_f := 1999;
        ELSIF x = 4528 THEN
            tanh_f := 1999;
        ELSIF x = 4529 THEN
            tanh_f := 1999;
        ELSIF x = 4530 THEN
            tanh_f := 1999;
        ELSIF x = 4531 THEN
            tanh_f := 1999;
        ELSIF x = 4532 THEN
            tanh_f := 1999;
        ELSIF x = 4533 THEN
            tanh_f := 1999;
        ELSIF x = 4534 THEN
            tanh_f := 1999;
        ELSIF x = 4535 THEN
            tanh_f := 1999;
        ELSIF x = 4536 THEN
            tanh_f := 1999;
        ELSIF x = 4537 THEN
            tanh_f := 1999;
        ELSIF x = 4538 THEN
            tanh_f := 1999;
        ELSIF x = 4539 THEN
            tanh_f := 1999;
        ELSIF x = 4540 THEN
            tanh_f := 1999;
        ELSIF x = 4541 THEN
            tanh_f := 1999;
        ELSIF x = 4542 THEN
            tanh_f := 1999;
        ELSIF x = 4543 THEN
            tanh_f := 1999;
        ELSIF x = 4544 THEN
            tanh_f := 1999;
        ELSIF x = 4545 THEN
            tanh_f := 1999;
        ELSIF x = 4546 THEN
            tanh_f := 1999;
        ELSIF x = 4547 THEN
            tanh_f := 2000;
        ELSIF x = 4548 THEN
            tanh_f := 2000;
        ELSIF x = 4549 THEN
            tanh_f := 2000;
        ELSIF x = 4550 THEN
            tanh_f := 2000;
        ELSIF x = 4551 THEN
            tanh_f := 2000;
        ELSIF x = 4552 THEN
            tanh_f := 2000;
        ELSIF x = 4553 THEN
            tanh_f := 2000;
        ELSIF x = 4554 THEN
            tanh_f := 2000;
        ELSIF x = 4555 THEN
            tanh_f := 2000;
        ELSIF x = 4556 THEN
            tanh_f := 2000;
        ELSIF x = 4557 THEN
            tanh_f := 2000;
        ELSIF x = 4558 THEN
            tanh_f := 2000;
        ELSIF x = 4559 THEN
            tanh_f := 2000;
        ELSIF x = 4560 THEN
            tanh_f := 2000;
        ELSIF x = 4561 THEN
            tanh_f := 2000;
        ELSIF x = 4562 THEN
            tanh_f := 2000;
        ELSIF x = 4563 THEN
            tanh_f := 2000;
        ELSIF x = 4564 THEN
            tanh_f := 2000;
        ELSIF x = 4565 THEN
            tanh_f := 2000;
        ELSIF x = 4566 THEN
            tanh_f := 2000;
        ELSIF x = 4567 THEN
            tanh_f := 2000;
        ELSIF x = 4568 THEN
            tanh_f := 2001;
        ELSIF x = 4569 THEN
            tanh_f := 2001;
        ELSIF x = 4570 THEN
            tanh_f := 2001;
        ELSIF x = 4571 THEN
            tanh_f := 2001;
        ELSIF x = 4572 THEN
            tanh_f := 2001;
        ELSIF x = 4573 THEN
            tanh_f := 2001;
        ELSIF x = 4574 THEN
            tanh_f := 2001;
        ELSIF x = 4575 THEN
            tanh_f := 2001;
        ELSIF x = 4576 THEN
            tanh_f := 2001;
        ELSIF x = 4577 THEN
            tanh_f := 2001;
        ELSIF x = 4578 THEN
            tanh_f := 2001;
        ELSIF x = 4579 THEN
            tanh_f := 2001;
        ELSIF x = 4580 THEN
            tanh_f := 2001;
        ELSIF x = 4581 THEN
            tanh_f := 2001;
        ELSIF x = 4582 THEN
            tanh_f := 2001;
        ELSIF x = 4583 THEN
            tanh_f := 2001;
        ELSIF x = 4584 THEN
            tanh_f := 2001;
        ELSIF x = 4585 THEN
            tanh_f := 2001;
        ELSIF x = 4586 THEN
            tanh_f := 2001;
        ELSIF x = 4587 THEN
            tanh_f := 2001;
        ELSIF x = 4588 THEN
            tanh_f := 2002;
        ELSIF x = 4589 THEN
            tanh_f := 2002;
        ELSIF x = 4590 THEN
            tanh_f := 2002;
        ELSIF x = 4591 THEN
            tanh_f := 2002;
        ELSIF x = 4592 THEN
            tanh_f := 2002;
        ELSIF x = 4593 THEN
            tanh_f := 2002;
        ELSIF x = 4594 THEN
            tanh_f := 2002;
        ELSIF x = 4595 THEN
            tanh_f := 2002;
        ELSIF x = 4596 THEN
            tanh_f := 2002;
        ELSIF x = 4597 THEN
            tanh_f := 2002;
        ELSIF x = 4598 THEN
            tanh_f := 2002;
        ELSIF x = 4599 THEN
            tanh_f := 2002;
        ELSIF x = 4600 THEN
            tanh_f := 2002;
        ELSIF x = 4601 THEN
            tanh_f := 2002;
        ELSIF x = 4602 THEN
            tanh_f := 2002;
        ELSIF x = 4603 THEN
            tanh_f := 2002;
        ELSIF x = 4604 THEN
            tanh_f := 2002;
        ELSIF x = 4605 THEN
            tanh_f := 2002;
        ELSIF x = 4606 THEN
            tanh_f := 2002;
        ELSIF x = 4607 THEN
            tanh_f := 2002;
        ELSIF x = 4608 THEN
            tanh_f := 2003;
        ELSIF x = 4609 THEN
            tanh_f := 2003;
        ELSIF x = 4610 THEN
            tanh_f := 2003;
        ELSIF x = 4611 THEN
            tanh_f := 2003;
        ELSIF x = 4612 THEN
            tanh_f := 2003;
        ELSIF x = 4613 THEN
            tanh_f := 2003;
        ELSIF x = 4614 THEN
            tanh_f := 2003;
        ELSIF x = 4615 THEN
            tanh_f := 2003;
        ELSIF x = 4616 THEN
            tanh_f := 2003;
        ELSIF x = 4617 THEN
            tanh_f := 2003;
        ELSIF x = 4618 THEN
            tanh_f := 2003;
        ELSIF x = 4619 THEN
            tanh_f := 2003;
        ELSIF x = 4620 THEN
            tanh_f := 2003;
        ELSIF x = 4621 THEN
            tanh_f := 2003;
        ELSIF x = 4622 THEN
            tanh_f := 2003;
        ELSIF x = 4623 THEN
            tanh_f := 2003;
        ELSIF x = 4624 THEN
            tanh_f := 2003;
        ELSIF x = 4625 THEN
            tanh_f := 2003;
        ELSIF x = 4626 THEN
            tanh_f := 2003;
        ELSIF x = 4627 THEN
            tanh_f := 2003;
        ELSIF x = 4628 THEN
            tanh_f := 2003;
        ELSIF x = 4629 THEN
            tanh_f := 2003;
        ELSIF x = 4630 THEN
            tanh_f := 2003;
        ELSIF x = 4631 THEN
            tanh_f := 2003;
        ELSIF x = 4632 THEN
            tanh_f := 2003;
        ELSIF x = 4633 THEN
            tanh_f := 2004;
        ELSIF x = 4634 THEN
            tanh_f := 2004;
        ELSIF x = 4635 THEN
            tanh_f := 2004;
        ELSIF x = 4636 THEN
            tanh_f := 2004;
        ELSIF x = 4637 THEN
            tanh_f := 2004;
        ELSIF x = 4638 THEN
            tanh_f := 2004;
        ELSIF x = 4639 THEN
            tanh_f := 2004;
        ELSIF x = 4640 THEN
            tanh_f := 2004;
        ELSIF x = 4641 THEN
            tanh_f := 2004;
        ELSIF x = 4642 THEN
            tanh_f := 2004;
        ELSIF x = 4643 THEN
            tanh_f := 2004;
        ELSIF x = 4644 THEN
            tanh_f := 2004;
        ELSIF x = 4645 THEN
            tanh_f := 2004;
        ELSIF x = 4646 THEN
            tanh_f := 2004;
        ELSIF x = 4647 THEN
            tanh_f := 2004;
        ELSIF x = 4648 THEN
            tanh_f := 2004;
        ELSIF x = 4649 THEN
            tanh_f := 2004;
        ELSIF x = 4650 THEN
            tanh_f := 2004;
        ELSIF x = 4651 THEN
            tanh_f := 2004;
        ELSIF x = 4652 THEN
            tanh_f := 2004;
        ELSIF x = 4653 THEN
            tanh_f := 2004;
        ELSIF x = 4654 THEN
            tanh_f := 2004;
        ELSIF x = 4655 THEN
            tanh_f := 2004;
        ELSIF x = 4656 THEN
            tanh_f := 2004;
        ELSIF x = 4657 THEN
            tanh_f := 2005;
        ELSIF x = 4658 THEN
            tanh_f := 2005;
        ELSIF x = 4659 THEN
            tanh_f := 2005;
        ELSIF x = 4660 THEN
            tanh_f := 2005;
        ELSIF x = 4661 THEN
            tanh_f := 2005;
        ELSIF x = 4662 THEN
            tanh_f := 2005;
        ELSIF x = 4663 THEN
            tanh_f := 2005;
        ELSIF x = 4664 THEN
            tanh_f := 2005;
        ELSIF x = 4665 THEN
            tanh_f := 2005;
        ELSIF x = 4666 THEN
            tanh_f := 2005;
        ELSIF x = 4667 THEN
            tanh_f := 2005;
        ELSIF x = 4668 THEN
            tanh_f := 2005;
        ELSIF x = 4669 THEN
            tanh_f := 2005;
        ELSIF x = 4670 THEN
            tanh_f := 2005;
        ELSIF x = 4671 THEN
            tanh_f := 2005;
        ELSIF x = 4672 THEN
            tanh_f := 2005;
        ELSIF x = 4673 THEN
            tanh_f := 2005;
        ELSIF x = 4674 THEN
            tanh_f := 2005;
        ELSIF x = 4675 THEN
            tanh_f := 2005;
        ELSIF x = 4676 THEN
            tanh_f := 2005;
        ELSIF x = 4677 THEN
            tanh_f := 2005;
        ELSIF x = 4678 THEN
            tanh_f := 2005;
        ELSIF x = 4679 THEN
            tanh_f := 2005;
        ELSIF x = 4680 THEN
            tanh_f := 2005;
        ELSIF x = 4681 THEN
            tanh_f := 2005;
        ELSIF x = 4682 THEN
            tanh_f := 2006;
        ELSIF x = 4683 THEN
            tanh_f := 2006;
        ELSIF x = 4684 THEN
            tanh_f := 2006;
        ELSIF x = 4685 THEN
            tanh_f := 2006;
        ELSIF x = 4686 THEN
            tanh_f := 2006;
        ELSIF x = 4687 THEN
            tanh_f := 2006;
        ELSIF x = 4688 THEN
            tanh_f := 2006;
        ELSIF x = 4689 THEN
            tanh_f := 2006;
        ELSIF x = 4690 THEN
            tanh_f := 2006;
        ELSIF x = 4691 THEN
            tanh_f := 2006;
        ELSIF x = 4692 THEN
            tanh_f := 2006;
        ELSIF x = 4693 THEN
            tanh_f := 2006;
        ELSIF x = 4694 THEN
            tanh_f := 2006;
        ELSIF x = 4695 THEN
            tanh_f := 2006;
        ELSIF x = 4696 THEN
            tanh_f := 2006;
        ELSIF x = 4697 THEN
            tanh_f := 2006;
        ELSIF x = 4698 THEN
            tanh_f := 2006;
        ELSIF x = 4699 THEN
            tanh_f := 2006;
        ELSIF x = 4700 THEN
            tanh_f := 2006;
        ELSIF x = 4701 THEN
            tanh_f := 2006;
        ELSIF x = 4702 THEN
            tanh_f := 2006;
        ELSIF x = 4703 THEN
            tanh_f := 2006;
        ELSIF x = 4704 THEN
            tanh_f := 2006;
        ELSIF x = 4705 THEN
            tanh_f := 2006;
        ELSIF x = 4706 THEN
            tanh_f := 2007;
        ELSIF x = 4707 THEN
            tanh_f := 2007;
        ELSIF x = 4708 THEN
            tanh_f := 2007;
        ELSIF x = 4709 THEN
            tanh_f := 2007;
        ELSIF x = 4710 THEN
            tanh_f := 2007;
        ELSIF x = 4711 THEN
            tanh_f := 2007;
        ELSIF x = 4712 THEN
            tanh_f := 2007;
        ELSIF x = 4713 THEN
            tanh_f := 2007;
        ELSIF x = 4714 THEN
            tanh_f := 2007;
        ELSIF x = 4715 THEN
            tanh_f := 2007;
        ELSIF x = 4716 THEN
            tanh_f := 2007;
        ELSIF x = 4717 THEN
            tanh_f := 2007;
        ELSIF x = 4718 THEN
            tanh_f := 2007;
        ELSIF x = 4719 THEN
            tanh_f := 2007;
        ELSIF x = 4720 THEN
            tanh_f := 2007;
        ELSIF x = 4721 THEN
            tanh_f := 2007;
        ELSIF x = 4722 THEN
            tanh_f := 2007;
        ELSIF x = 4723 THEN
            tanh_f := 2007;
        ELSIF x = 4724 THEN
            tanh_f := 2007;
        ELSIF x = 4725 THEN
            tanh_f := 2007;
        ELSIF x = 4726 THEN
            tanh_f := 2007;
        ELSIF x = 4727 THEN
            tanh_f := 2007;
        ELSIF x = 4728 THEN
            tanh_f := 2007;
        ELSIF x = 4729 THEN
            tanh_f := 2007;
        ELSIF x = 4730 THEN
            tanh_f := 2008;
        ELSIF x = 4731 THEN
            tanh_f := 2008;
        ELSIF x = 4732 THEN
            tanh_f := 2008;
        ELSIF x = 4733 THEN
            tanh_f := 2008;
        ELSIF x = 4734 THEN
            tanh_f := 2008;
        ELSIF x = 4735 THEN
            tanh_f := 2008;
        ELSIF x = 4736 THEN
            tanh_f := 2008;
        ELSIF x = 4737 THEN
            tanh_f := 2008;
        ELSIF x = 4738 THEN
            tanh_f := 2008;
        ELSIF x = 4739 THEN
            tanh_f := 2008;
        ELSIF x = 4740 THEN
            tanh_f := 2008;
        ELSIF x = 4741 THEN
            tanh_f := 2008;
        ELSIF x = 4742 THEN
            tanh_f := 2008;
        ELSIF x = 4743 THEN
            tanh_f := 2008;
        ELSIF x = 4744 THEN
            tanh_f := 2008;
        ELSIF x = 4745 THEN
            tanh_f := 2008;
        ELSIF x = 4746 THEN
            tanh_f := 2008;
        ELSIF x = 4747 THEN
            tanh_f := 2008;
        ELSIF x = 4748 THEN
            tanh_f := 2008;
        ELSIF x = 4749 THEN
            tanh_f := 2008;
        ELSIF x = 4750 THEN
            tanh_f := 2008;
        ELSIF x = 4751 THEN
            tanh_f := 2008;
        ELSIF x = 4752 THEN
            tanh_f := 2008;
        ELSIF x = 4753 THEN
            tanh_f := 2008;
        ELSIF x = 4754 THEN
            tanh_f := 2008;
        ELSIF x = 4755 THEN
            tanh_f := 2009;
        ELSIF x = 4756 THEN
            tanh_f := 2009;
        ELSIF x = 4757 THEN
            tanh_f := 2009;
        ELSIF x = 4758 THEN
            tanh_f := 2009;
        ELSIF x = 4759 THEN
            tanh_f := 2009;
        ELSIF x = 4760 THEN
            tanh_f := 2009;
        ELSIF x = 4761 THEN
            tanh_f := 2009;
        ELSIF x = 4762 THEN
            tanh_f := 2009;
        ELSIF x = 4763 THEN
            tanh_f := 2009;
        ELSIF x = 4764 THEN
            tanh_f := 2009;
        ELSIF x = 4765 THEN
            tanh_f := 2009;
        ELSIF x = 4766 THEN
            tanh_f := 2009;
        ELSIF x = 4767 THEN
            tanh_f := 2009;
        ELSIF x = 4768 THEN
            tanh_f := 2009;
        ELSIF x = 4769 THEN
            tanh_f := 2009;
        ELSIF x = 4770 THEN
            tanh_f := 2009;
        ELSIF x = 4771 THEN
            tanh_f := 2009;
        ELSIF x = 4772 THEN
            tanh_f := 2009;
        ELSIF x = 4773 THEN
            tanh_f := 2009;
        ELSIF x = 4774 THEN
            tanh_f := 2009;
        ELSIF x = 4775 THEN
            tanh_f := 2009;
        ELSIF x = 4776 THEN
            tanh_f := 2009;
        ELSIF x = 4777 THEN
            tanh_f := 2009;
        ELSIF x = 4778 THEN
            tanh_f := 2009;
        ELSIF x = 4779 THEN
            tanh_f := 2010;
        ELSIF x = 4780 THEN
            tanh_f := 2010;
        ELSIF x = 4781 THEN
            tanh_f := 2010;
        ELSIF x = 4782 THEN
            tanh_f := 2010;
        ELSIF x = 4783 THEN
            tanh_f := 2010;
        ELSIF x = 4784 THEN
            tanh_f := 2010;
        ELSIF x = 4785 THEN
            tanh_f := 2010;
        ELSIF x = 4786 THEN
            tanh_f := 2010;
        ELSIF x = 4787 THEN
            tanh_f := 2010;
        ELSIF x = 4788 THEN
            tanh_f := 2010;
        ELSIF x = 4789 THEN
            tanh_f := 2010;
        ELSIF x = 4790 THEN
            tanh_f := 2010;
        ELSIF x = 4791 THEN
            tanh_f := 2010;
        ELSIF x = 4792 THEN
            tanh_f := 2010;
        ELSIF x = 4793 THEN
            tanh_f := 2010;
        ELSIF x = 4794 THEN
            tanh_f := 2010;
        ELSIF x = 4795 THEN
            tanh_f := 2010;
        ELSIF x = 4796 THEN
            tanh_f := 2010;
        ELSIF x = 4797 THEN
            tanh_f := 2010;
        ELSIF x = 4798 THEN
            tanh_f := 2010;
        ELSIF x = 4799 THEN
            tanh_f := 2010;
        ELSIF x = 4800 THEN
            tanh_f := 2010;
        ELSIF x = 4801 THEN
            tanh_f := 2010;
        ELSIF x = 4802 THEN
            tanh_f := 2010;
        ELSIF x = 4803 THEN
            tanh_f := 2010;
        ELSIF x = 4804 THEN
            tanh_f := 2011;
        ELSIF x = 4805 THEN
            tanh_f := 2011;
        ELSIF x = 4806 THEN
            tanh_f := 2011;
        ELSIF x = 4807 THEN
            tanh_f := 2011;
        ELSIF x = 4808 THEN
            tanh_f := 2011;
        ELSIF x = 4809 THEN
            tanh_f := 2011;
        ELSIF x = 4810 THEN
            tanh_f := 2011;
        ELSIF x = 4811 THEN
            tanh_f := 2011;
        ELSIF x = 4812 THEN
            tanh_f := 2011;
        ELSIF x = 4813 THEN
            tanh_f := 2011;
        ELSIF x = 4814 THEN
            tanh_f := 2011;
        ELSIF x = 4815 THEN
            tanh_f := 2011;
        ELSIF x = 4816 THEN
            tanh_f := 2011;
        ELSIF x = 4817 THEN
            tanh_f := 2011;
        ELSIF x = 4818 THEN
            tanh_f := 2011;
        ELSIF x = 4819 THEN
            tanh_f := 2011;
        ELSIF x = 4820 THEN
            tanh_f := 2011;
        ELSIF x = 4821 THEN
            tanh_f := 2011;
        ELSIF x = 4822 THEN
            tanh_f := 2011;
        ELSIF x = 4823 THEN
            tanh_f := 2011;
        ELSIF x = 4824 THEN
            tanh_f := 2011;
        ELSIF x = 4825 THEN
            tanh_f := 2011;
        ELSIF x = 4826 THEN
            tanh_f := 2011;
        ELSIF x = 4827 THEN
            tanh_f := 2011;
        ELSIF x = 4828 THEN
            tanh_f := 2012;
        ELSIF x = 4829 THEN
            tanh_f := 2012;
        ELSIF x = 4830 THEN
            tanh_f := 2012;
        ELSIF x = 4831 THEN
            tanh_f := 2012;
        ELSIF x = 4832 THEN
            tanh_f := 2012;
        ELSIF x = 4833 THEN
            tanh_f := 2012;
        ELSIF x = 4834 THEN
            tanh_f := 2012;
        ELSIF x = 4835 THEN
            tanh_f := 2012;
        ELSIF x = 4836 THEN
            tanh_f := 2012;
        ELSIF x = 4837 THEN
            tanh_f := 2012;
        ELSIF x = 4838 THEN
            tanh_f := 2012;
        ELSIF x = 4839 THEN
            tanh_f := 2012;
        ELSIF x = 4840 THEN
            tanh_f := 2012;
        ELSIF x = 4841 THEN
            tanh_f := 2012;
        ELSIF x = 4842 THEN
            tanh_f := 2012;
        ELSIF x = 4843 THEN
            tanh_f := 2012;
        ELSIF x = 4844 THEN
            tanh_f := 2012;
        ELSIF x = 4845 THEN
            tanh_f := 2012;
        ELSIF x = 4846 THEN
            tanh_f := 2012;
        ELSIF x = 4847 THEN
            tanh_f := 2012;
        ELSIF x = 4848 THEN
            tanh_f := 2012;
        ELSIF x = 4849 THEN
            tanh_f := 2012;
        ELSIF x = 4850 THEN
            tanh_f := 2012;
        ELSIF x = 4851 THEN
            tanh_f := 2012;
        ELSIF x = 4852 THEN
            tanh_f := 2013;
        ELSIF x = 4853 THEN
            tanh_f := 2013;
        ELSIF x = 4854 THEN
            tanh_f := 2013;
        ELSIF x = 4855 THEN
            tanh_f := 2013;
        ELSIF x = 4856 THEN
            tanh_f := 2013;
        ELSIF x = 4857 THEN
            tanh_f := 2013;
        ELSIF x = 4858 THEN
            tanh_f := 2013;
        ELSIF x = 4859 THEN
            tanh_f := 2013;
        ELSIF x = 4860 THEN
            tanh_f := 2013;
        ELSIF x = 4861 THEN
            tanh_f := 2013;
        ELSIF x = 4862 THEN
            tanh_f := 2013;
        ELSIF x = 4863 THEN
            tanh_f := 2013;
        ELSIF x = 4864 THEN
            tanh_f := 2013;
        ELSIF x = 4865 THEN
            tanh_f := 2013;
        ELSIF x = 4866 THEN
            tanh_f := 2013;
        ELSIF x = 4867 THEN
            tanh_f := 2013;
        ELSIF x = 4868 THEN
            tanh_f := 2013;
        ELSIF x = 4869 THEN
            tanh_f := 2013;
        ELSIF x = 4870 THEN
            tanh_f := 2013;
        ELSIF x = 4871 THEN
            tanh_f := 2013;
        ELSIF x = 4872 THEN
            tanh_f := 2013;
        ELSIF x = 4873 THEN
            tanh_f := 2013;
        ELSIF x = 4874 THEN
            tanh_f := 2013;
        ELSIF x = 4875 THEN
            tanh_f := 2013;
        ELSIF x = 4876 THEN
            tanh_f := 2013;
        ELSIF x = 4877 THEN
            tanh_f := 2013;
        ELSIF x = 4878 THEN
            tanh_f := 2013;
        ELSIF x = 4879 THEN
            tanh_f := 2013;
        ELSIF x = 4880 THEN
            tanh_f := 2013;
        ELSIF x = 4881 THEN
            tanh_f := 2013;
        ELSIF x = 4882 THEN
            tanh_f := 2013;
        ELSIF x = 4883 THEN
            tanh_f := 2013;
        ELSIF x = 4884 THEN
            tanh_f := 2014;
        ELSIF x = 4885 THEN
            tanh_f := 2014;
        ELSIF x = 4886 THEN
            tanh_f := 2014;
        ELSIF x = 4887 THEN
            tanh_f := 2014;
        ELSIF x = 4888 THEN
            tanh_f := 2014;
        ELSIF x = 4889 THEN
            tanh_f := 2014;
        ELSIF x = 4890 THEN
            tanh_f := 2014;
        ELSIF x = 4891 THEN
            tanh_f := 2014;
        ELSIF x = 4892 THEN
            tanh_f := 2014;
        ELSIF x = 4893 THEN
            tanh_f := 2014;
        ELSIF x = 4894 THEN
            tanh_f := 2014;
        ELSIF x = 4895 THEN
            tanh_f := 2014;
        ELSIF x = 4896 THEN
            tanh_f := 2014;
        ELSIF x = 4897 THEN
            tanh_f := 2014;
        ELSIF x = 4898 THEN
            tanh_f := 2014;
        ELSIF x = 4899 THEN
            tanh_f := 2014;
        ELSIF x = 4900 THEN
            tanh_f := 2014;
        ELSIF x = 4901 THEN
            tanh_f := 2014;
        ELSIF x = 4902 THEN
            tanh_f := 2014;
        ELSIF x = 4903 THEN
            tanh_f := 2014;
        ELSIF x = 4904 THEN
            tanh_f := 2014;
        ELSIF x = 4905 THEN
            tanh_f := 2014;
        ELSIF x = 4906 THEN
            tanh_f := 2014;
        ELSIF x = 4907 THEN
            tanh_f := 2014;
        ELSIF x = 4908 THEN
            tanh_f := 2014;
        ELSIF x = 4909 THEN
            tanh_f := 2014;
        ELSIF x = 4910 THEN
            tanh_f := 2014;
        ELSIF x = 4911 THEN
            tanh_f := 2014;
        ELSIF x = 4912 THEN
            tanh_f := 2014;
        ELSIF x = 4913 THEN
            tanh_f := 2014;
        ELSIF x = 4914 THEN
            tanh_f := 2014;
        ELSIF x = 4915 THEN
            tanh_f := 2014;
        ELSIF x = 4916 THEN
            tanh_f := 2014;
        ELSIF x = 4917 THEN
            tanh_f := 2014;
        ELSIF x = 4918 THEN
            tanh_f := 2014;
        ELSIF x = 4919 THEN
            tanh_f := 2014;
        ELSIF x = 4920 THEN
            tanh_f := 2014;
        ELSIF x = 4921 THEN
            tanh_f := 2014;
        ELSIF x = 4922 THEN
            tanh_f := 2014;
        ELSIF x = 4923 THEN
            tanh_f := 2014;
        ELSIF x = 4924 THEN
            tanh_f := 2015;
        ELSIF x = 4925 THEN
            tanh_f := 2015;
        ELSIF x = 4926 THEN
            tanh_f := 2015;
        ELSIF x = 4927 THEN
            tanh_f := 2015;
        ELSIF x = 4928 THEN
            tanh_f := 2015;
        ELSIF x = 4929 THEN
            tanh_f := 2015;
        ELSIF x = 4930 THEN
            tanh_f := 2015;
        ELSIF x = 4931 THEN
            tanh_f := 2015;
        ELSIF x = 4932 THEN
            tanh_f := 2015;
        ELSIF x = 4933 THEN
            tanh_f := 2015;
        ELSIF x = 4934 THEN
            tanh_f := 2015;
        ELSIF x = 4935 THEN
            tanh_f := 2015;
        ELSIF x = 4936 THEN
            tanh_f := 2015;
        ELSIF x = 4937 THEN
            tanh_f := 2015;
        ELSIF x = 4938 THEN
            tanh_f := 2015;
        ELSIF x = 4939 THEN
            tanh_f := 2015;
        ELSIF x = 4940 THEN
            tanh_f := 2015;
        ELSIF x = 4941 THEN
            tanh_f := 2015;
        ELSIF x = 4942 THEN
            tanh_f := 2015;
        ELSIF x = 4943 THEN
            tanh_f := 2015;
        ELSIF x = 4944 THEN
            tanh_f := 2015;
        ELSIF x = 4945 THEN
            tanh_f := 2015;
        ELSIF x = 4946 THEN
            tanh_f := 2015;
        ELSIF x = 4947 THEN
            tanh_f := 2015;
        ELSIF x = 4948 THEN
            tanh_f := 2015;
        ELSIF x = 4949 THEN
            tanh_f := 2015;
        ELSIF x = 4950 THEN
            tanh_f := 2015;
        ELSIF x = 4951 THEN
            tanh_f := 2015;
        ELSIF x = 4952 THEN
            tanh_f := 2015;
        ELSIF x = 4953 THEN
            tanh_f := 2015;
        ELSIF x = 4954 THEN
            tanh_f := 2015;
        ELSIF x = 4955 THEN
            tanh_f := 2015;
        ELSIF x = 4956 THEN
            tanh_f := 2015;
        ELSIF x = 4957 THEN
            tanh_f := 2015;
        ELSIF x = 4958 THEN
            tanh_f := 2015;
        ELSIF x = 4959 THEN
            tanh_f := 2015;
        ELSIF x = 4960 THEN
            tanh_f := 2015;
        ELSIF x = 4961 THEN
            tanh_f := 2015;
        ELSIF x = 4962 THEN
            tanh_f := 2015;
        ELSIF x = 4963 THEN
            tanh_f := 2016;
        ELSIF x = 4964 THEN
            tanh_f := 2016;
        ELSIF x = 4965 THEN
            tanh_f := 2016;
        ELSIF x = 4966 THEN
            tanh_f := 2016;
        ELSIF x = 4967 THEN
            tanh_f := 2016;
        ELSIF x = 4968 THEN
            tanh_f := 2016;
        ELSIF x = 4969 THEN
            tanh_f := 2016;
        ELSIF x = 4970 THEN
            tanh_f := 2016;
        ELSIF x = 4971 THEN
            tanh_f := 2016;
        ELSIF x = 4972 THEN
            tanh_f := 2016;
        ELSIF x = 4973 THEN
            tanh_f := 2016;
        ELSIF x = 4974 THEN
            tanh_f := 2016;
        ELSIF x = 4975 THEN
            tanh_f := 2016;
        ELSIF x = 4976 THEN
            tanh_f := 2016;
        ELSIF x = 4977 THEN
            tanh_f := 2016;
        ELSIF x = 4978 THEN
            tanh_f := 2016;
        ELSIF x = 4979 THEN
            tanh_f := 2016;
        ELSIF x = 4980 THEN
            tanh_f := 2016;
        ELSIF x = 4981 THEN
            tanh_f := 2016;
        ELSIF x = 4982 THEN
            tanh_f := 2016;
        ELSIF x = 4983 THEN
            tanh_f := 2016;
        ELSIF x = 4984 THEN
            tanh_f := 2016;
        ELSIF x = 4985 THEN
            tanh_f := 2016;
        ELSIF x = 4986 THEN
            tanh_f := 2016;
        ELSIF x = 4987 THEN
            tanh_f := 2016;
        ELSIF x = 4988 THEN
            tanh_f := 2016;
        ELSIF x = 4989 THEN
            tanh_f := 2016;
        ELSIF x = 4990 THEN
            tanh_f := 2016;
        ELSIF x = 4991 THEN
            tanh_f := 2016;
        ELSIF x = 4992 THEN
            tanh_f := 2016;
        ELSIF x = 4993 THEN
            tanh_f := 2016;
        ELSIF x = 4994 THEN
            tanh_f := 2016;
        ELSIF x = 4995 THEN
            tanh_f := 2016;
        ELSIF x = 4996 THEN
            tanh_f := 2016;
        ELSIF x = 4997 THEN
            tanh_f := 2016;
        ELSIF x = 4998 THEN
            tanh_f := 2016;
        ELSIF x = 4999 THEN
            tanh_f := 2016;
        ELSIF x = 5000 THEN
            tanh_f := 2016;
        ELSIF x = 5001 THEN
            tanh_f := 2016;
        ELSIF x = 5002 THEN
            tanh_f := 2017;
        ELSIF x = 5003 THEN
            tanh_f := 2017;
        ELSIF x = 5004 THEN
            tanh_f := 2017;
        ELSIF x = 5005 THEN
            tanh_f := 2017;
        ELSIF x = 5006 THEN
            tanh_f := 2017;
        ELSIF x = 5007 THEN
            tanh_f := 2017;
        ELSIF x = 5008 THEN
            tanh_f := 2017;
        ELSIF x = 5009 THEN
            tanh_f := 2017;
        ELSIF x = 5010 THEN
            tanh_f := 2017;
        ELSIF x = 5011 THEN
            tanh_f := 2017;
        ELSIF x = 5012 THEN
            tanh_f := 2017;
        ELSIF x = 5013 THEN
            tanh_f := 2017;
        ELSIF x = 5014 THEN
            tanh_f := 2017;
        ELSIF x = 5015 THEN
            tanh_f := 2017;
        ELSIF x = 5016 THEN
            tanh_f := 2017;
        ELSIF x = 5017 THEN
            tanh_f := 2017;
        ELSIF x = 5018 THEN
            tanh_f := 2017;
        ELSIF x = 5019 THEN
            tanh_f := 2017;
        ELSIF x = 5020 THEN
            tanh_f := 2017;
        ELSIF x = 5021 THEN
            tanh_f := 2017;
        ELSIF x = 5022 THEN
            tanh_f := 2017;
        ELSIF x = 5023 THEN
            tanh_f := 2017;
        ELSIF x = 5024 THEN
            tanh_f := 2017;
        ELSIF x = 5025 THEN
            tanh_f := 2017;
        ELSIF x = 5026 THEN
            tanh_f := 2017;
        ELSIF x = 5027 THEN
            tanh_f := 2017;
        ELSIF x = 5028 THEN
            tanh_f := 2017;
        ELSIF x = 5029 THEN
            tanh_f := 2017;
        ELSIF x = 5030 THEN
            tanh_f := 2017;
        ELSIF x = 5031 THEN
            tanh_f := 2017;
        ELSIF x = 5032 THEN
            tanh_f := 2017;
        ELSIF x = 5033 THEN
            tanh_f := 2017;
        ELSIF x = 5034 THEN
            tanh_f := 2017;
        ELSIF x = 5035 THEN
            tanh_f := 2017;
        ELSIF x = 5036 THEN
            tanh_f := 2017;
        ELSIF x = 5037 THEN
            tanh_f := 2017;
        ELSIF x = 5038 THEN
            tanh_f := 2017;
        ELSIF x = 5039 THEN
            tanh_f := 2017;
        ELSIF x = 5040 THEN
            tanh_f := 2017;
        ELSIF x = 5041 THEN
            tanh_f := 2017;
        ELSIF x = 5042 THEN
            tanh_f := 2018;
        ELSIF x = 5043 THEN
            tanh_f := 2018;
        ELSIF x = 5044 THEN
            tanh_f := 2018;
        ELSIF x = 5045 THEN
            tanh_f := 2018;
        ELSIF x = 5046 THEN
            tanh_f := 2018;
        ELSIF x = 5047 THEN
            tanh_f := 2018;
        ELSIF x = 5048 THEN
            tanh_f := 2018;
        ELSIF x = 5049 THEN
            tanh_f := 2018;
        ELSIF x = 5050 THEN
            tanh_f := 2018;
        ELSIF x = 5051 THEN
            tanh_f := 2018;
        ELSIF x = 5052 THEN
            tanh_f := 2018;
        ELSIF x = 5053 THEN
            tanh_f := 2018;
        ELSIF x = 5054 THEN
            tanh_f := 2018;
        ELSIF x = 5055 THEN
            tanh_f := 2018;
        ELSIF x = 5056 THEN
            tanh_f := 2018;
        ELSIF x = 5057 THEN
            tanh_f := 2018;
        ELSIF x = 5058 THEN
            tanh_f := 2018;
        ELSIF x = 5059 THEN
            tanh_f := 2018;
        ELSIF x = 5060 THEN
            tanh_f := 2018;
        ELSIF x = 5061 THEN
            tanh_f := 2018;
        ELSIF x = 5062 THEN
            tanh_f := 2018;
        ELSIF x = 5063 THEN
            tanh_f := 2018;
        ELSIF x = 5064 THEN
            tanh_f := 2018;
        ELSIF x = 5065 THEN
            tanh_f := 2018;
        ELSIF x = 5066 THEN
            tanh_f := 2018;
        ELSIF x = 5067 THEN
            tanh_f := 2018;
        ELSIF x = 5068 THEN
            tanh_f := 2018;
        ELSIF x = 5069 THEN
            tanh_f := 2018;
        ELSIF x = 5070 THEN
            tanh_f := 2018;
        ELSIF x = 5071 THEN
            tanh_f := 2018;
        ELSIF x = 5072 THEN
            tanh_f := 2018;
        ELSIF x = 5073 THEN
            tanh_f := 2018;
        ELSIF x = 5074 THEN
            tanh_f := 2018;
        ELSIF x = 5075 THEN
            tanh_f := 2018;
        ELSIF x = 5076 THEN
            tanh_f := 2018;
        ELSIF x = 5077 THEN
            tanh_f := 2018;
        ELSIF x = 5078 THEN
            tanh_f := 2018;
        ELSIF x = 5079 THEN
            tanh_f := 2018;
        ELSIF x = 5080 THEN
            tanh_f := 2018;
        ELSIF x = 5081 THEN
            tanh_f := 2019;
        ELSIF x = 5082 THEN
            tanh_f := 2019;
        ELSIF x = 5083 THEN
            tanh_f := 2019;
        ELSIF x = 5084 THEN
            tanh_f := 2019;
        ELSIF x = 5085 THEN
            tanh_f := 2019;
        ELSIF x = 5086 THEN
            tanh_f := 2019;
        ELSIF x = 5087 THEN
            tanh_f := 2019;
        ELSIF x = 5088 THEN
            tanh_f := 2019;
        ELSIF x = 5089 THEN
            tanh_f := 2019;
        ELSIF x = 5090 THEN
            tanh_f := 2019;
        ELSIF x = 5091 THEN
            tanh_f := 2019;
        ELSIF x = 5092 THEN
            tanh_f := 2019;
        ELSIF x = 5093 THEN
            tanh_f := 2019;
        ELSIF x = 5094 THEN
            tanh_f := 2019;
        ELSIF x = 5095 THEN
            tanh_f := 2019;
        ELSIF x = 5096 THEN
            tanh_f := 2019;
        ELSIF x = 5097 THEN
            tanh_f := 2019;
        ELSIF x = 5098 THEN
            tanh_f := 2019;
        ELSIF x = 5099 THEN
            tanh_f := 2019;
        ELSIF x = 5100 THEN
            tanh_f := 2019;
        ELSIF x = 5101 THEN
            tanh_f := 2019;
        ELSIF x = 5102 THEN
            tanh_f := 2019;
        ELSIF x = 5103 THEN
            tanh_f := 2019;
        ELSIF x = 5104 THEN
            tanh_f := 2019;
        ELSIF x = 5105 THEN
            tanh_f := 2019;
        ELSIF x = 5106 THEN
            tanh_f := 2019;
        ELSIF x = 5107 THEN
            tanh_f := 2019;
        ELSIF x = 5108 THEN
            tanh_f := 2019;
        ELSIF x = 5109 THEN
            tanh_f := 2019;
        ELSIF x = 5110 THEN
            tanh_f := 2019;
        ELSIF x = 5111 THEN
            tanh_f := 2019;
        ELSIF x = 5112 THEN
            tanh_f := 2019;
        ELSIF x = 5113 THEN
            tanh_f := 2019;
        ELSIF x = 5114 THEN
            tanh_f := 2019;
        ELSIF x = 5115 THEN
            tanh_f := 2019;
        ELSIF x = 5116 THEN
            tanh_f := 2019;
        ELSIF x = 5117 THEN
            tanh_f := 2019;
        ELSIF x = 5118 THEN
            tanh_f := 2019;
        ELSIF x = 5119 THEN
            tanh_f := 2019;
        ELSIF x = 5120 THEN
            tanh_f := 2020;
        ELSIF x = 5121 THEN
            tanh_f := 2020;
        ELSIF x = 5122 THEN
            tanh_f := 2020;
        ELSIF x = 5123 THEN
            tanh_f := 2020;
        ELSIF x = 5124 THEN
            tanh_f := 2020;
        ELSIF x = 5125 THEN
            tanh_f := 2020;
        ELSIF x = 5126 THEN
            tanh_f := 2020;
        ELSIF x = 5127 THEN
            tanh_f := 2020;
        ELSIF x = 5128 THEN
            tanh_f := 2020;
        ELSIF x = 5129 THEN
            tanh_f := 2020;
        ELSIF x = 5130 THEN
            tanh_f := 2020;
        ELSIF x = 5131 THEN
            tanh_f := 2020;
        ELSIF x = 5132 THEN
            tanh_f := 2020;
        ELSIF x = 5133 THEN
            tanh_f := 2020;
        ELSIF x = 5134 THEN
            tanh_f := 2020;
        ELSIF x = 5135 THEN
            tanh_f := 2020;
        ELSIF x = 5136 THEN
            tanh_f := 2020;
        ELSIF x = 5137 THEN
            tanh_f := 2020;
        ELSIF x = 5138 THEN
            tanh_f := 2020;
        ELSIF x = 5139 THEN
            tanh_f := 2020;
        ELSIF x = 5140 THEN
            tanh_f := 2020;
        ELSIF x = 5141 THEN
            tanh_f := 2020;
        ELSIF x = 5142 THEN
            tanh_f := 2020;
        ELSIF x = 5143 THEN
            tanh_f := 2020;
        ELSIF x = 5144 THEN
            tanh_f := 2020;
        ELSIF x = 5145 THEN
            tanh_f := 2020;
        ELSIF x = 5146 THEN
            tanh_f := 2020;
        ELSIF x = 5147 THEN
            tanh_f := 2020;
        ELSIF x = 5148 THEN
            tanh_f := 2020;
        ELSIF x = 5149 THEN
            tanh_f := 2020;
        ELSIF x = 5150 THEN
            tanh_f := 2020;
        ELSIF x = 5151 THEN
            tanh_f := 2020;
        ELSIF x = 5152 THEN
            tanh_f := 2020;
        ELSIF x = 5153 THEN
            tanh_f := 2020;
        ELSIF x = 5154 THEN
            tanh_f := 2020;
        ELSIF x = 5155 THEN
            tanh_f := 2020;
        ELSIF x = 5156 THEN
            tanh_f := 2020;
        ELSIF x = 5157 THEN
            tanh_f := 2021;
        ELSIF x = 5158 THEN
            tanh_f := 2021;
        ELSIF x = 5159 THEN
            tanh_f := 2021;
        ELSIF x = 5160 THEN
            tanh_f := 2021;
        ELSIF x = 5161 THEN
            tanh_f := 2021;
        ELSIF x = 5162 THEN
            tanh_f := 2021;
        ELSIF x = 5163 THEN
            tanh_f := 2021;
        ELSIF x = 5164 THEN
            tanh_f := 2021;
        ELSIF x = 5165 THEN
            tanh_f := 2021;
        ELSIF x = 5166 THEN
            tanh_f := 2021;
        ELSIF x = 5167 THEN
            tanh_f := 2021;
        ELSIF x = 5168 THEN
            tanh_f := 2021;
        ELSIF x = 5169 THEN
            tanh_f := 2021;
        ELSIF x = 5170 THEN
            tanh_f := 2021;
        ELSIF x = 5171 THEN
            tanh_f := 2021;
        ELSIF x = 5172 THEN
            tanh_f := 2021;
        ELSIF x = 5173 THEN
            tanh_f := 2021;
        ELSIF x = 5174 THEN
            tanh_f := 2021;
        ELSIF x = 5175 THEN
            tanh_f := 2021;
        ELSIF x = 5176 THEN
            tanh_f := 2021;
        ELSIF x = 5177 THEN
            tanh_f := 2021;
        ELSIF x = 5178 THEN
            tanh_f := 2021;
        ELSIF x = 5179 THEN
            tanh_f := 2021;
        ELSIF x = 5180 THEN
            tanh_f := 2021;
        ELSIF x = 5181 THEN
            tanh_f := 2021;
        ELSIF x = 5182 THEN
            tanh_f := 2021;
        ELSIF x = 5183 THEN
            tanh_f := 2021;
        ELSIF x = 5184 THEN
            tanh_f := 2021;
        ELSIF x = 5185 THEN
            tanh_f := 2021;
        ELSIF x = 5186 THEN
            tanh_f := 2021;
        ELSIF x = 5187 THEN
            tanh_f := 2021;
        ELSIF x = 5188 THEN
            tanh_f := 2021;
        ELSIF x = 5189 THEN
            tanh_f := 2021;
        ELSIF x = 5190 THEN
            tanh_f := 2021;
        ELSIF x = 5191 THEN
            tanh_f := 2021;
        ELSIF x = 5192 THEN
            tanh_f := 2021;
        ELSIF x = 5193 THEN
            tanh_f := 2021;
        ELSIF x = 5194 THEN
            tanh_f := 2022;
        ELSIF x = 5195 THEN
            tanh_f := 2022;
        ELSIF x = 5196 THEN
            tanh_f := 2022;
        ELSIF x = 5197 THEN
            tanh_f := 2022;
        ELSIF x = 5198 THEN
            tanh_f := 2022;
        ELSIF x = 5199 THEN
            tanh_f := 2022;
        ELSIF x = 5200 THEN
            tanh_f := 2022;
        ELSIF x = 5201 THEN
            tanh_f := 2022;
        ELSIF x = 5202 THEN
            tanh_f := 2022;
        ELSIF x = 5203 THEN
            tanh_f := 2022;
        ELSIF x = 5204 THEN
            tanh_f := 2022;
        ELSIF x = 5205 THEN
            tanh_f := 2022;
        ELSIF x = 5206 THEN
            tanh_f := 2022;
        ELSIF x = 5207 THEN
            tanh_f := 2022;
        ELSIF x = 5208 THEN
            tanh_f := 2022;
        ELSIF x = 5209 THEN
            tanh_f := 2022;
        ELSIF x = 5210 THEN
            tanh_f := 2022;
        ELSIF x = 5211 THEN
            tanh_f := 2022;
        ELSIF x = 5212 THEN
            tanh_f := 2022;
        ELSIF x = 5213 THEN
            tanh_f := 2022;
        ELSIF x = 5214 THEN
            tanh_f := 2022;
        ELSIF x = 5215 THEN
            tanh_f := 2022;
        ELSIF x = 5216 THEN
            tanh_f := 2022;
        ELSIF x = 5217 THEN
            tanh_f := 2022;
        ELSIF x = 5218 THEN
            tanh_f := 2022;
        ELSIF x = 5219 THEN
            tanh_f := 2022;
        ELSIF x = 5220 THEN
            tanh_f := 2022;
        ELSIF x = 5221 THEN
            tanh_f := 2022;
        ELSIF x = 5222 THEN
            tanh_f := 2022;
        ELSIF x = 5223 THEN
            tanh_f := 2022;
        ELSIF x = 5224 THEN
            tanh_f := 2022;
        ELSIF x = 5225 THEN
            tanh_f := 2022;
        ELSIF x = 5226 THEN
            tanh_f := 2022;
        ELSIF x = 5227 THEN
            tanh_f := 2022;
        ELSIF x = 5228 THEN
            tanh_f := 2022;
        ELSIF x = 5229 THEN
            tanh_f := 2022;
        ELSIF x = 5230 THEN
            tanh_f := 2023;
        ELSIF x = 5231 THEN
            tanh_f := 2023;
        ELSIF x = 5232 THEN
            tanh_f := 2023;
        ELSIF x = 5233 THEN
            tanh_f := 2023;
        ELSIF x = 5234 THEN
            tanh_f := 2023;
        ELSIF x = 5235 THEN
            tanh_f := 2023;
        ELSIF x = 5236 THEN
            tanh_f := 2023;
        ELSIF x = 5237 THEN
            tanh_f := 2023;
        ELSIF x = 5238 THEN
            tanh_f := 2023;
        ELSIF x = 5239 THEN
            tanh_f := 2023;
        ELSIF x = 5240 THEN
            tanh_f := 2023;
        ELSIF x = 5241 THEN
            tanh_f := 2023;
        ELSIF x = 5242 THEN
            tanh_f := 2023;
        ELSIF x = 5243 THEN
            tanh_f := 2023;
        ELSIF x = 5244 THEN
            tanh_f := 2023;
        ELSIF x = 5245 THEN
            tanh_f := 2023;
        ELSIF x = 5246 THEN
            tanh_f := 2023;
        ELSIF x = 5247 THEN
            tanh_f := 2023;
        ELSIF x = 5248 THEN
            tanh_f := 2023;
        ELSIF x = 5249 THEN
            tanh_f := 2023;
        ELSIF x = 5250 THEN
            tanh_f := 2023;
        ELSIF x = 5251 THEN
            tanh_f := 2023;
        ELSIF x = 5252 THEN
            tanh_f := 2023;
        ELSIF x = 5253 THEN
            tanh_f := 2023;
        ELSIF x = 5254 THEN
            tanh_f := 2023;
        ELSIF x = 5255 THEN
            tanh_f := 2023;
        ELSIF x = 5256 THEN
            tanh_f := 2023;
        ELSIF x = 5257 THEN
            tanh_f := 2023;
        ELSIF x = 5258 THEN
            tanh_f := 2023;
        ELSIF x = 5259 THEN
            tanh_f := 2023;
        ELSIF x = 5260 THEN
            tanh_f := 2023;
        ELSIF x = 5261 THEN
            tanh_f := 2023;
        ELSIF x = 5262 THEN
            tanh_f := 2023;
        ELSIF x = 5263 THEN
            tanh_f := 2023;
        ELSIF x = 5264 THEN
            tanh_f := 2023;
        ELSIF x = 5265 THEN
            tanh_f := 2023;
        ELSIF x = 5266 THEN
            tanh_f := 2023;
        ELSIF x = 5267 THEN
            tanh_f := 2024;
        ELSIF x = 5268 THEN
            tanh_f := 2024;
        ELSIF x = 5269 THEN
            tanh_f := 2024;
        ELSIF x = 5270 THEN
            tanh_f := 2024;
        ELSIF x = 5271 THEN
            tanh_f := 2024;
        ELSIF x = 5272 THEN
            tanh_f := 2024;
        ELSIF x = 5273 THEN
            tanh_f := 2024;
        ELSIF x = 5274 THEN
            tanh_f := 2024;
        ELSIF x = 5275 THEN
            tanh_f := 2024;
        ELSIF x = 5276 THEN
            tanh_f := 2024;
        ELSIF x = 5277 THEN
            tanh_f := 2024;
        ELSIF x = 5278 THEN
            tanh_f := 2024;
        ELSIF x = 5279 THEN
            tanh_f := 2024;
        ELSIF x = 5280 THEN
            tanh_f := 2024;
        ELSIF x = 5281 THEN
            tanh_f := 2024;
        ELSIF x = 5282 THEN
            tanh_f := 2024;
        ELSIF x = 5283 THEN
            tanh_f := 2024;
        ELSIF x = 5284 THEN
            tanh_f := 2024;
        ELSIF x = 5285 THEN
            tanh_f := 2024;
        ELSIF x = 5286 THEN
            tanh_f := 2024;
        ELSIF x = 5287 THEN
            tanh_f := 2024;
        ELSIF x = 5288 THEN
            tanh_f := 2024;
        ELSIF x = 5289 THEN
            tanh_f := 2024;
        ELSIF x = 5290 THEN
            tanh_f := 2024;
        ELSIF x = 5291 THEN
            tanh_f := 2024;
        ELSIF x = 5292 THEN
            tanh_f := 2024;
        ELSIF x = 5293 THEN
            tanh_f := 2024;
        ELSIF x = 5294 THEN
            tanh_f := 2024;
        ELSIF x = 5295 THEN
            tanh_f := 2024;
        ELSIF x = 5296 THEN
            tanh_f := 2024;
        ELSIF x = 5297 THEN
            tanh_f := 2024;
        ELSIF x = 5298 THEN
            tanh_f := 2024;
        ELSIF x = 5299 THEN
            tanh_f := 2024;
        ELSIF x = 5300 THEN
            tanh_f := 2024;
        ELSIF x = 5301 THEN
            tanh_f := 2024;
        ELSIF x = 5302 THEN
            tanh_f := 2024;
        ELSIF x = 5303 THEN
            tanh_f := 2025;
        ELSIF x = 5304 THEN
            tanh_f := 2025;
        ELSIF x = 5305 THEN
            tanh_f := 2025;
        ELSIF x = 5306 THEN
            tanh_f := 2025;
        ELSIF x = 5307 THEN
            tanh_f := 2025;
        ELSIF x = 5308 THEN
            tanh_f := 2025;
        ELSIF x = 5309 THEN
            tanh_f := 2025;
        ELSIF x = 5310 THEN
            tanh_f := 2025;
        ELSIF x = 5311 THEN
            tanh_f := 2025;
        ELSIF x = 5312 THEN
            tanh_f := 2025;
        ELSIF x = 5313 THEN
            tanh_f := 2025;
        ELSIF x = 5314 THEN
            tanh_f := 2025;
        ELSIF x = 5315 THEN
            tanh_f := 2025;
        ELSIF x = 5316 THEN
            tanh_f := 2025;
        ELSIF x = 5317 THEN
            tanh_f := 2025;
        ELSIF x = 5318 THEN
            tanh_f := 2025;
        ELSIF x = 5319 THEN
            tanh_f := 2025;
        ELSIF x = 5320 THEN
            tanh_f := 2025;
        ELSIF x = 5321 THEN
            tanh_f := 2025;
        ELSIF x = 5322 THEN
            tanh_f := 2025;
        ELSIF x = 5323 THEN
            tanh_f := 2025;
        ELSIF x = 5324 THEN
            tanh_f := 2025;
        ELSIF x = 5325 THEN
            tanh_f := 2025;
        ELSIF x = 5326 THEN
            tanh_f := 2025;
        ELSIF x = 5327 THEN
            tanh_f := 2025;
        ELSIF x = 5328 THEN
            tanh_f := 2025;
        ELSIF x = 5329 THEN
            tanh_f := 2025;
        ELSIF x = 5330 THEN
            tanh_f := 2025;
        ELSIF x = 5331 THEN
            tanh_f := 2025;
        ELSIF x = 5332 THEN
            tanh_f := 2025;
        ELSIF x = 5333 THEN
            tanh_f := 2025;
        ELSIF x = 5334 THEN
            tanh_f := 2025;
        ELSIF x = 5335 THEN
            tanh_f := 2025;
        ELSIF x = 5336 THEN
            tanh_f := 2025;
        ELSIF x = 5337 THEN
            tanh_f := 2025;
        ELSIF x = 5338 THEN
            tanh_f := 2025;
        ELSIF x = 5339 THEN
            tanh_f := 2025;
        ELSIF x = 5340 THEN
            tanh_f := 2026;
        ELSIF x = 5341 THEN
            tanh_f := 2026;
        ELSIF x = 5342 THEN
            tanh_f := 2026;
        ELSIF x = 5343 THEN
            tanh_f := 2026;
        ELSIF x = 5344 THEN
            tanh_f := 2026;
        ELSIF x = 5345 THEN
            tanh_f := 2026;
        ELSIF x = 5346 THEN
            tanh_f := 2026;
        ELSIF x = 5347 THEN
            tanh_f := 2026;
        ELSIF x = 5348 THEN
            tanh_f := 2026;
        ELSIF x = 5349 THEN
            tanh_f := 2026;
        ELSIF x = 5350 THEN
            tanh_f := 2026;
        ELSIF x = 5351 THEN
            tanh_f := 2026;
        ELSIF x = 5352 THEN
            tanh_f := 2026;
        ELSIF x = 5353 THEN
            tanh_f := 2026;
        ELSIF x = 5354 THEN
            tanh_f := 2026;
        ELSIF x = 5355 THEN
            tanh_f := 2026;
        ELSIF x = 5356 THEN
            tanh_f := 2026;
        ELSIF x = 5357 THEN
            tanh_f := 2026;
        ELSIF x = 5358 THEN
            tanh_f := 2026;
        ELSIF x = 5359 THEN
            tanh_f := 2026;
        ELSIF x = 5360 THEN
            tanh_f := 2026;
        ELSIF x = 5361 THEN
            tanh_f := 2026;
        ELSIF x = 5362 THEN
            tanh_f := 2026;
        ELSIF x = 5363 THEN
            tanh_f := 2026;
        ELSIF x = 5364 THEN
            tanh_f := 2026;
        ELSIF x = 5365 THEN
            tanh_f := 2026;
        ELSIF x = 5366 THEN
            tanh_f := 2026;
        ELSIF x = 5367 THEN
            tanh_f := 2026;
        ELSIF x = 5368 THEN
            tanh_f := 2026;
        ELSIF x = 5369 THEN
            tanh_f := 2026;
        ELSIF x = 5370 THEN
            tanh_f := 2026;
        ELSIF x = 5371 THEN
            tanh_f := 2026;
        ELSIF x = 5372 THEN
            tanh_f := 2026;
        ELSIF x = 5373 THEN
            tanh_f := 2026;
        ELSIF x = 5374 THEN
            tanh_f := 2026;
        ELSIF x = 5375 THEN
            tanh_f := 2026;
        ELSIF x = 5376 THEN
            tanh_f := 2026;
        ELSIF x = 5377 THEN
            tanh_f := 2026;
        ELSIF x = 5378 THEN
            tanh_f := 2026;
        ELSIF x = 5379 THEN
            tanh_f := 2026;
        ELSIF x = 5380 THEN
            tanh_f := 2026;
        ELSIF x = 5381 THEN
            tanh_f := 2026;
        ELSIF x = 5382 THEN
            tanh_f := 2026;
        ELSIF x = 5383 THEN
            tanh_f := 2026;
        ELSIF x = 5384 THEN
            tanh_f := 2026;
        ELSIF x = 5385 THEN
            tanh_f := 2026;
        ELSIF x = 5386 THEN
            tanh_f := 2026;
        ELSIF x = 5387 THEN
            tanh_f := 2026;
        ELSIF x = 5388 THEN
            tanh_f := 2026;
        ELSIF x = 5389 THEN
            tanh_f := 2026;
        ELSIF x = 5390 THEN
            tanh_f := 2026;
        ELSIF x = 5391 THEN
            tanh_f := 2026;
        ELSIF x = 5392 THEN
            tanh_f := 2026;
        ELSIF x = 5393 THEN
            tanh_f := 2026;
        ELSIF x = 5394 THEN
            tanh_f := 2026;
        ELSIF x = 5395 THEN
            tanh_f := 2026;
        ELSIF x = 5396 THEN
            tanh_f := 2026;
        ELSIF x = 5397 THEN
            tanh_f := 2026;
        ELSIF x = 5398 THEN
            tanh_f := 2026;
        ELSIF x = 5399 THEN
            tanh_f := 2026;
        ELSIF x = 5400 THEN
            tanh_f := 2026;
        ELSIF x = 5401 THEN
            tanh_f := 2026;
        ELSIF x = 5402 THEN
            tanh_f := 2026;
        ELSIF x = 5403 THEN
            tanh_f := 2026;
        ELSIF x = 5404 THEN
            tanh_f := 2026;
        ELSIF x = 5405 THEN
            tanh_f := 2026;
        ELSIF x = 5406 THEN
            tanh_f := 2026;
        ELSIF x = 5407 THEN
            tanh_f := 2026;
        ELSIF x = 5408 THEN
            tanh_f := 2026;
        ELSIF x = 5409 THEN
            tanh_f := 2026;
        ELSIF x = 5410 THEN
            tanh_f := 2026;
        ELSIF x = 5411 THEN
            tanh_f := 2026;
        ELSIF x = 5412 THEN
            tanh_f := 2026;
        ELSIF x = 5413 THEN
            tanh_f := 2026;
        ELSIF x = 5414 THEN
            tanh_f := 2026;
        ELSIF x = 5415 THEN
            tanh_f := 2026;
        ELSIF x = 5416 THEN
            tanh_f := 2026;
        ELSIF x = 5417 THEN
            tanh_f := 2026;
        ELSIF x = 5418 THEN
            tanh_f := 2026;
        ELSIF x = 5419 THEN
            tanh_f := 2027;
        ELSIF x = 5420 THEN
            tanh_f := 2027;
        ELSIF x = 5421 THEN
            tanh_f := 2027;
        ELSIF x = 5422 THEN
            tanh_f := 2027;
        ELSIF x = 5423 THEN
            tanh_f := 2027;
        ELSIF x = 5424 THEN
            tanh_f := 2027;
        ELSIF x = 5425 THEN
            tanh_f := 2027;
        ELSIF x = 5426 THEN
            tanh_f := 2027;
        ELSIF x = 5427 THEN
            tanh_f := 2027;
        ELSIF x = 5428 THEN
            tanh_f := 2027;
        ELSIF x = 5429 THEN
            tanh_f := 2027;
        ELSIF x = 5430 THEN
            tanh_f := 2027;
        ELSIF x = 5431 THEN
            tanh_f := 2027;
        ELSIF x = 5432 THEN
            tanh_f := 2027;
        ELSIF x = 5433 THEN
            tanh_f := 2027;
        ELSIF x = 5434 THEN
            tanh_f := 2027;
        ELSIF x = 5435 THEN
            tanh_f := 2027;
        ELSIF x = 5436 THEN
            tanh_f := 2027;
        ELSIF x = 5437 THEN
            tanh_f := 2027;
        ELSIF x = 5438 THEN
            tanh_f := 2027;
        ELSIF x = 5439 THEN
            tanh_f := 2027;
        ELSIF x = 5440 THEN
            tanh_f := 2027;
        ELSIF x = 5441 THEN
            tanh_f := 2027;
        ELSIF x = 5442 THEN
            tanh_f := 2027;
        ELSIF x = 5443 THEN
            tanh_f := 2027;
        ELSIF x = 5444 THEN
            tanh_f := 2027;
        ELSIF x = 5445 THEN
            tanh_f := 2027;
        ELSIF x = 5446 THEN
            tanh_f := 2027;
        ELSIF x = 5447 THEN
            tanh_f := 2027;
        ELSIF x = 5448 THEN
            tanh_f := 2027;
        ELSIF x = 5449 THEN
            tanh_f := 2027;
        ELSIF x = 5450 THEN
            tanh_f := 2027;
        ELSIF x = 5451 THEN
            tanh_f := 2027;
        ELSIF x = 5452 THEN
            tanh_f := 2027;
        ELSIF x = 5453 THEN
            tanh_f := 2027;
        ELSIF x = 5454 THEN
            tanh_f := 2027;
        ELSIF x = 5455 THEN
            tanh_f := 2027;
        ELSIF x = 5456 THEN
            tanh_f := 2027;
        ELSIF x = 5457 THEN
            tanh_f := 2027;
        ELSIF x = 5458 THEN
            tanh_f := 2027;
        ELSIF x = 5459 THEN
            tanh_f := 2027;
        ELSIF x = 5460 THEN
            tanh_f := 2027;
        ELSIF x = 5461 THEN
            tanh_f := 2027;
        ELSIF x = 5462 THEN
            tanh_f := 2028;
        ELSIF x = 5463 THEN
            tanh_f := 2028;
        ELSIF x = 5464 THEN
            tanh_f := 2028;
        ELSIF x = 5465 THEN
            tanh_f := 2028;
        ELSIF x = 5466 THEN
            tanh_f := 2028;
        ELSIF x = 5467 THEN
            tanh_f := 2028;
        ELSIF x = 5468 THEN
            tanh_f := 2028;
        ELSIF x = 5469 THEN
            tanh_f := 2028;
        ELSIF x = 5470 THEN
            tanh_f := 2028;
        ELSIF x = 5471 THEN
            tanh_f := 2028;
        ELSIF x = 5472 THEN
            tanh_f := 2028;
        ELSIF x = 5473 THEN
            tanh_f := 2028;
        ELSIF x = 5474 THEN
            tanh_f := 2028;
        ELSIF x = 5475 THEN
            tanh_f := 2028;
        ELSIF x = 5476 THEN
            tanh_f := 2028;
        ELSIF x = 5477 THEN
            tanh_f := 2028;
        ELSIF x = 5478 THEN
            tanh_f := 2028;
        ELSIF x = 5479 THEN
            tanh_f := 2028;
        ELSIF x = 5480 THEN
            tanh_f := 2028;
        ELSIF x = 5481 THEN
            tanh_f := 2028;
        ELSIF x = 5482 THEN
            tanh_f := 2028;
        ELSIF x = 5483 THEN
            tanh_f := 2028;
        ELSIF x = 5484 THEN
            tanh_f := 2028;
        ELSIF x = 5485 THEN
            tanh_f := 2028;
        ELSIF x = 5486 THEN
            tanh_f := 2028;
        ELSIF x = 5487 THEN
            tanh_f := 2028;
        ELSIF x = 5488 THEN
            tanh_f := 2028;
        ELSIF x = 5489 THEN
            tanh_f := 2028;
        ELSIF x = 5490 THEN
            tanh_f := 2028;
        ELSIF x = 5491 THEN
            tanh_f := 2028;
        ELSIF x = 5492 THEN
            tanh_f := 2028;
        ELSIF x = 5493 THEN
            tanh_f := 2028;
        ELSIF x = 5494 THEN
            tanh_f := 2028;
        ELSIF x = 5495 THEN
            tanh_f := 2028;
        ELSIF x = 5496 THEN
            tanh_f := 2028;
        ELSIF x = 5497 THEN
            tanh_f := 2028;
        ELSIF x = 5498 THEN
            tanh_f := 2028;
        ELSIF x = 5499 THEN
            tanh_f := 2028;
        ELSIF x = 5500 THEN
            tanh_f := 2028;
        ELSIF x = 5501 THEN
            tanh_f := 2028;
        ELSIF x = 5502 THEN
            tanh_f := 2028;
        ELSIF x = 5503 THEN
            tanh_f := 2028;
        ELSIF x = 5504 THEN
            tanh_f := 2029;
        ELSIF x = 5505 THEN
            tanh_f := 2029;
        ELSIF x = 5506 THEN
            tanh_f := 2029;
        ELSIF x = 5507 THEN
            tanh_f := 2029;
        ELSIF x = 5508 THEN
            tanh_f := 2029;
        ELSIF x = 5509 THEN
            tanh_f := 2029;
        ELSIF x = 5510 THEN
            tanh_f := 2029;
        ELSIF x = 5511 THEN
            tanh_f := 2029;
        ELSIF x = 5512 THEN
            tanh_f := 2029;
        ELSIF x = 5513 THEN
            tanh_f := 2029;
        ELSIF x = 5514 THEN
            tanh_f := 2029;
        ELSIF x = 5515 THEN
            tanh_f := 2029;
        ELSIF x = 5516 THEN
            tanh_f := 2029;
        ELSIF x = 5517 THEN
            tanh_f := 2029;
        ELSIF x = 5518 THEN
            tanh_f := 2029;
        ELSIF x = 5519 THEN
            tanh_f := 2029;
        ELSIF x = 5520 THEN
            tanh_f := 2029;
        ELSIF x = 5521 THEN
            tanh_f := 2029;
        ELSIF x = 5522 THEN
            tanh_f := 2029;
        ELSIF x = 5523 THEN
            tanh_f := 2029;
        ELSIF x = 5524 THEN
            tanh_f := 2029;
        ELSIF x = 5525 THEN
            tanh_f := 2029;
        ELSIF x = 5526 THEN
            tanh_f := 2029;
        ELSIF x = 5527 THEN
            tanh_f := 2029;
        ELSIF x = 5528 THEN
            tanh_f := 2029;
        ELSIF x = 5529 THEN
            tanh_f := 2029;
        ELSIF x = 5530 THEN
            tanh_f := 2029;
        ELSIF x = 5531 THEN
            tanh_f := 2029;
        ELSIF x = 5532 THEN
            tanh_f := 2029;
        ELSIF x = 5533 THEN
            tanh_f := 2029;
        ELSIF x = 5534 THEN
            tanh_f := 2029;
        ELSIF x = 5535 THEN
            tanh_f := 2029;
        ELSIF x = 5536 THEN
            tanh_f := 2029;
        ELSIF x = 5537 THEN
            tanh_f := 2029;
        ELSIF x = 5538 THEN
            tanh_f := 2029;
        ELSIF x = 5539 THEN
            tanh_f := 2029;
        ELSIF x = 5540 THEN
            tanh_f := 2029;
        ELSIF x = 5541 THEN
            tanh_f := 2029;
        ELSIF x = 5542 THEN
            tanh_f := 2029;
        ELSIF x = 5543 THEN
            tanh_f := 2029;
        ELSIF x = 5544 THEN
            tanh_f := 2029;
        ELSIF x = 5545 THEN
            tanh_f := 2029;
        ELSIF x = 5546 THEN
            tanh_f := 2029;
        ELSIF x = 5547 THEN
            tanh_f := 2030;
        ELSIF x = 5548 THEN
            tanh_f := 2030;
        ELSIF x = 5549 THEN
            tanh_f := 2030;
        ELSIF x = 5550 THEN
            tanh_f := 2030;
        ELSIF x = 5551 THEN
            tanh_f := 2030;
        ELSIF x = 5552 THEN
            tanh_f := 2030;
        ELSIF x = 5553 THEN
            tanh_f := 2030;
        ELSIF x = 5554 THEN
            tanh_f := 2030;
        ELSIF x = 5555 THEN
            tanh_f := 2030;
        ELSIF x = 5556 THEN
            tanh_f := 2030;
        ELSIF x = 5557 THEN
            tanh_f := 2030;
        ELSIF x = 5558 THEN
            tanh_f := 2030;
        ELSIF x = 5559 THEN
            tanh_f := 2030;
        ELSIF x = 5560 THEN
            tanh_f := 2030;
        ELSIF x = 5561 THEN
            tanh_f := 2030;
        ELSIF x = 5562 THEN
            tanh_f := 2030;
        ELSIF x = 5563 THEN
            tanh_f := 2030;
        ELSIF x = 5564 THEN
            tanh_f := 2030;
        ELSIF x = 5565 THEN
            tanh_f := 2030;
        ELSIF x = 5566 THEN
            tanh_f := 2030;
        ELSIF x = 5567 THEN
            tanh_f := 2030;
        ELSIF x = 5568 THEN
            tanh_f := 2030;
        ELSIF x = 5569 THEN
            tanh_f := 2030;
        ELSIF x = 5570 THEN
            tanh_f := 2030;
        ELSIF x = 5571 THEN
            tanh_f := 2030;
        ELSIF x = 5572 THEN
            tanh_f := 2030;
        ELSIF x = 5573 THEN
            tanh_f := 2030;
        ELSIF x = 5574 THEN
            tanh_f := 2030;
        ELSIF x = 5575 THEN
            tanh_f := 2030;
        ELSIF x = 5576 THEN
            tanh_f := 2030;
        ELSIF x = 5577 THEN
            tanh_f := 2030;
        ELSIF x = 5578 THEN
            tanh_f := 2030;
        ELSIF x = 5579 THEN
            tanh_f := 2030;
        ELSIF x = 5580 THEN
            tanh_f := 2030;
        ELSIF x = 5581 THEN
            tanh_f := 2030;
        ELSIF x = 5582 THEN
            tanh_f := 2030;
        ELSIF x = 5583 THEN
            tanh_f := 2030;
        ELSIF x = 5584 THEN
            tanh_f := 2030;
        ELSIF x = 5585 THEN
            tanh_f := 2030;
        ELSIF x = 5586 THEN
            tanh_f := 2030;
        ELSIF x = 5587 THEN
            tanh_f := 2030;
        ELSIF x = 5588 THEN
            tanh_f := 2030;
        ELSIF x = 5589 THEN
            tanh_f := 2030;
        ELSIF x = 5590 THEN
            tanh_f := 2031;
        ELSIF x = 5591 THEN
            tanh_f := 2031;
        ELSIF x = 5592 THEN
            tanh_f := 2031;
        ELSIF x = 5593 THEN
            tanh_f := 2031;
        ELSIF x = 5594 THEN
            tanh_f := 2031;
        ELSIF x = 5595 THEN
            tanh_f := 2031;
        ELSIF x = 5596 THEN
            tanh_f := 2031;
        ELSIF x = 5597 THEN
            tanh_f := 2031;
        ELSIF x = 5598 THEN
            tanh_f := 2031;
        ELSIF x = 5599 THEN
            tanh_f := 2031;
        ELSIF x = 5600 THEN
            tanh_f := 2031;
        ELSIF x = 5601 THEN
            tanh_f := 2031;
        ELSIF x = 5602 THEN
            tanh_f := 2031;
        ELSIF x = 5603 THEN
            tanh_f := 2031;
        ELSIF x = 5604 THEN
            tanh_f := 2031;
        ELSIF x = 5605 THEN
            tanh_f := 2031;
        ELSIF x = 5606 THEN
            tanh_f := 2031;
        ELSIF x = 5607 THEN
            tanh_f := 2031;
        ELSIF x = 5608 THEN
            tanh_f := 2031;
        ELSIF x = 5609 THEN
            tanh_f := 2031;
        ELSIF x = 5610 THEN
            tanh_f := 2031;
        ELSIF x = 5611 THEN
            tanh_f := 2031;
        ELSIF x = 5612 THEN
            tanh_f := 2031;
        ELSIF x = 5613 THEN
            tanh_f := 2031;
        ELSIF x = 5614 THEN
            tanh_f := 2031;
        ELSIF x = 5615 THEN
            tanh_f := 2031;
        ELSIF x = 5616 THEN
            tanh_f := 2031;
        ELSIF x = 5617 THEN
            tanh_f := 2031;
        ELSIF x = 5618 THEN
            tanh_f := 2031;
        ELSIF x = 5619 THEN
            tanh_f := 2031;
        ELSIF x = 5620 THEN
            tanh_f := 2031;
        ELSIF x = 5621 THEN
            tanh_f := 2031;
        ELSIF x = 5622 THEN
            tanh_f := 2031;
        ELSIF x = 5623 THEN
            tanh_f := 2031;
        ELSIF x = 5624 THEN
            tanh_f := 2031;
        ELSIF x = 5625 THEN
            tanh_f := 2031;
        ELSIF x = 5626 THEN
            tanh_f := 2031;
        ELSIF x = 5627 THEN
            tanh_f := 2031;
        ELSIF x = 5628 THEN
            tanh_f := 2031;
        ELSIF x = 5629 THEN
            tanh_f := 2031;
        ELSIF x = 5630 THEN
            tanh_f := 2031;
        ELSIF x = 5631 THEN
            tanh_f := 2031;
        ELSIF x = 5632 THEN
            tanh_f := 2031;
        ELSIF x = 5633 THEN
            tanh_f := 2031;
        ELSIF x = 5634 THEN
            tanh_f := 2031;
        ELSIF x = 5635 THEN
            tanh_f := 2031;
        ELSIF x = 5636 THEN
            tanh_f := 2031;
        ELSIF x = 5637 THEN
            tanh_f := 2031;
        ELSIF x = 5638 THEN
            tanh_f := 2031;
        ELSIF x = 5639 THEN
            tanh_f := 2031;
        ELSIF x = 5640 THEN
            tanh_f := 2031;
        ELSIF x = 5641 THEN
            tanh_f := 2031;
        ELSIF x = 5642 THEN
            tanh_f := 2031;
        ELSIF x = 5643 THEN
            tanh_f := 2031;
        ELSIF x = 5644 THEN
            tanh_f := 2031;
        ELSIF x = 5645 THEN
            tanh_f := 2031;
        ELSIF x = 5646 THEN
            tanh_f := 2031;
        ELSIF x = 5647 THEN
            tanh_f := 2031;
        ELSIF x = 5648 THEN
            tanh_f := 2031;
        ELSIF x = 5649 THEN
            tanh_f := 2031;
        ELSIF x = 5650 THEN
            tanh_f := 2031;
        ELSIF x = 5651 THEN
            tanh_f := 2031;
        ELSIF x = 5652 THEN
            tanh_f := 2031;
        ELSIF x = 5653 THEN
            tanh_f := 2031;
        ELSIF x = 5654 THEN
            tanh_f := 2031;
        ELSIF x = 5655 THEN
            tanh_f := 2031;
        ELSIF x = 5656 THEN
            tanh_f := 2031;
        ELSIF x = 5657 THEN
            tanh_f := 2031;
        ELSIF x = 5658 THEN
            tanh_f := 2031;
        ELSIF x = 5659 THEN
            tanh_f := 2031;
        ELSIF x = 5660 THEN
            tanh_f := 2031;
        ELSIF x = 5661 THEN
            tanh_f := 2031;
        ELSIF x = 5662 THEN
            tanh_f := 2031;
        ELSIF x = 5663 THEN
            tanh_f := 2031;
        ELSIF x = 5664 THEN
            tanh_f := 2031;
        ELSIF x = 5665 THEN
            tanh_f := 2031;
        ELSIF x = 5666 THEN
            tanh_f := 2031;
        ELSIF x = 5667 THEN
            tanh_f := 2031;
        ELSIF x = 5668 THEN
            tanh_f := 2031;
        ELSIF x = 5669 THEN
            tanh_f := 2031;
        ELSIF x = 5670 THEN
            tanh_f := 2031;
        ELSIF x = 5671 THEN
            tanh_f := 2031;
        ELSIF x = 5672 THEN
            tanh_f := 2031;
        ELSIF x = 5673 THEN
            tanh_f := 2031;
        ELSIF x = 5674 THEN
            tanh_f := 2031;
        ELSIF x = 5675 THEN
            tanh_f := 2031;
        ELSIF x = 5676 THEN
            tanh_f := 2031;
        ELSIF x = 5677 THEN
            tanh_f := 2031;
        ELSIF x = 5678 THEN
            tanh_f := 2031;
        ELSIF x = 5679 THEN
            tanh_f := 2031;
        ELSIF x = 5680 THEN
            tanh_f := 2031;
        ELSIF x = 5681 THEN
            tanh_f := 2031;
        ELSIF x = 5682 THEN
            tanh_f := 2031;
        ELSIF x = 5683 THEN
            tanh_f := 2031;
        ELSIF x = 5684 THEN
            tanh_f := 2031;
        ELSIF x = 5685 THEN
            tanh_f := 2031;
        ELSIF x = 5686 THEN
            tanh_f := 2031;
        ELSIF x = 5687 THEN
            tanh_f := 2031;
        ELSIF x = 5688 THEN
            tanh_f := 2031;
        ELSIF x = 5689 THEN
            tanh_f := 2032;
        ELSIF x = 5690 THEN
            tanh_f := 2032;
        ELSIF x = 5691 THEN
            tanh_f := 2032;
        ELSIF x = 5692 THEN
            tanh_f := 2032;
        ELSIF x = 5693 THEN
            tanh_f := 2032;
        ELSIF x = 5694 THEN
            tanh_f := 2032;
        ELSIF x = 5695 THEN
            tanh_f := 2032;
        ELSIF x = 5696 THEN
            tanh_f := 2032;
        ELSIF x = 5697 THEN
            tanh_f := 2032;
        ELSIF x = 5698 THEN
            tanh_f := 2032;
        ELSIF x = 5699 THEN
            tanh_f := 2032;
        ELSIF x = 5700 THEN
            tanh_f := 2032;
        ELSIF x = 5701 THEN
            tanh_f := 2032;
        ELSIF x = 5702 THEN
            tanh_f := 2032;
        ELSIF x = 5703 THEN
            tanh_f := 2032;
        ELSIF x = 5704 THEN
            tanh_f := 2032;
        ELSIF x = 5705 THEN
            tanh_f := 2032;
        ELSIF x = 5706 THEN
            tanh_f := 2032;
        ELSIF x = 5707 THEN
            tanh_f := 2032;
        ELSIF x = 5708 THEN
            tanh_f := 2032;
        ELSIF x = 5709 THEN
            tanh_f := 2032;
        ELSIF x = 5710 THEN
            tanh_f := 2032;
        ELSIF x = 5711 THEN
            tanh_f := 2032;
        ELSIF x = 5712 THEN
            tanh_f := 2032;
        ELSIF x = 5713 THEN
            tanh_f := 2032;
        ELSIF x = 5714 THEN
            tanh_f := 2032;
        ELSIF x = 5715 THEN
            tanh_f := 2032;
        ELSIF x = 5716 THEN
            tanh_f := 2032;
        ELSIF x = 5717 THEN
            tanh_f := 2032;
        ELSIF x = 5718 THEN
            tanh_f := 2032;
        ELSIF x = 5719 THEN
            tanh_f := 2032;
        ELSIF x = 5720 THEN
            tanh_f := 2032;
        ELSIF x = 5721 THEN
            tanh_f := 2032;
        ELSIF x = 5722 THEN
            tanh_f := 2032;
        ELSIF x = 5723 THEN
            tanh_f := 2032;
        ELSIF x = 5724 THEN
            tanh_f := 2032;
        ELSIF x = 5725 THEN
            tanh_f := 2032;
        ELSIF x = 5726 THEN
            tanh_f := 2032;
        ELSIF x = 5727 THEN
            tanh_f := 2032;
        ELSIF x = 5728 THEN
            tanh_f := 2032;
        ELSIF x = 5729 THEN
            tanh_f := 2032;
        ELSIF x = 5730 THEN
            tanh_f := 2032;
        ELSIF x = 5731 THEN
            tanh_f := 2032;
        ELSIF x = 5732 THEN
            tanh_f := 2032;
        ELSIF x = 5733 THEN
            tanh_f := 2032;
        ELSIF x = 5734 THEN
            tanh_f := 2032;
        ELSIF x = 5735 THEN
            tanh_f := 2032;
        ELSIF x = 5736 THEN
            tanh_f := 2032;
        ELSIF x = 5737 THEN
            tanh_f := 2032;
        ELSIF x = 5738 THEN
            tanh_f := 2032;
        ELSIF x = 5739 THEN
            tanh_f := 2032;
        ELSIF x = 5740 THEN
            tanh_f := 2032;
        ELSIF x = 5741 THEN
            tanh_f := 2032;
        ELSIF x = 5742 THEN
            tanh_f := 2032;
        ELSIF x = 5743 THEN
            tanh_f := 2032;
        ELSIF x = 5744 THEN
            tanh_f := 2032;
        ELSIF x = 5745 THEN
            tanh_f := 2032;
        ELSIF x = 5746 THEN
            tanh_f := 2033;
        ELSIF x = 5747 THEN
            tanh_f := 2033;
        ELSIF x = 5748 THEN
            tanh_f := 2033;
        ELSIF x = 5749 THEN
            tanh_f := 2033;
        ELSIF x = 5750 THEN
            tanh_f := 2033;
        ELSIF x = 5751 THEN
            tanh_f := 2033;
        ELSIF x = 5752 THEN
            tanh_f := 2033;
        ELSIF x = 5753 THEN
            tanh_f := 2033;
        ELSIF x = 5754 THEN
            tanh_f := 2033;
        ELSIF x = 5755 THEN
            tanh_f := 2033;
        ELSIF x = 5756 THEN
            tanh_f := 2033;
        ELSIF x = 5757 THEN
            tanh_f := 2033;
        ELSIF x = 5758 THEN
            tanh_f := 2033;
        ELSIF x = 5759 THEN
            tanh_f := 2033;
        ELSIF x = 5760 THEN
            tanh_f := 2033;
        ELSIF x = 5761 THEN
            tanh_f := 2033;
        ELSIF x = 5762 THEN
            tanh_f := 2033;
        ELSIF x = 5763 THEN
            tanh_f := 2033;
        ELSIF x = 5764 THEN
            tanh_f := 2033;
        ELSIF x = 5765 THEN
            tanh_f := 2033;
        ELSIF x = 5766 THEN
            tanh_f := 2033;
        ELSIF x = 5767 THEN
            tanh_f := 2033;
        ELSIF x = 5768 THEN
            tanh_f := 2033;
        ELSIF x = 5769 THEN
            tanh_f := 2033;
        ELSIF x = 5770 THEN
            tanh_f := 2033;
        ELSIF x = 5771 THEN
            tanh_f := 2033;
        ELSIF x = 5772 THEN
            tanh_f := 2033;
        ELSIF x = 5773 THEN
            tanh_f := 2033;
        ELSIF x = 5774 THEN
            tanh_f := 2033;
        ELSIF x = 5775 THEN
            tanh_f := 2033;
        ELSIF x = 5776 THEN
            tanh_f := 2033;
        ELSIF x = 5777 THEN
            tanh_f := 2033;
        ELSIF x = 5778 THEN
            tanh_f := 2033;
        ELSIF x = 5779 THEN
            tanh_f := 2033;
        ELSIF x = 5780 THEN
            tanh_f := 2033;
        ELSIF x = 5781 THEN
            tanh_f := 2033;
        ELSIF x = 5782 THEN
            tanh_f := 2033;
        ELSIF x = 5783 THEN
            tanh_f := 2033;
        ELSIF x = 5784 THEN
            tanh_f := 2033;
        ELSIF x = 5785 THEN
            tanh_f := 2033;
        ELSIF x = 5786 THEN
            tanh_f := 2033;
        ELSIF x = 5787 THEN
            tanh_f := 2033;
        ELSIF x = 5788 THEN
            tanh_f := 2033;
        ELSIF x = 5789 THEN
            tanh_f := 2033;
        ELSIF x = 5790 THEN
            tanh_f := 2033;
        ELSIF x = 5791 THEN
            tanh_f := 2033;
        ELSIF x = 5792 THEN
            tanh_f := 2033;
        ELSIF x = 5793 THEN
            tanh_f := 2033;
        ELSIF x = 5794 THEN
            tanh_f := 2033;
        ELSIF x = 5795 THEN
            tanh_f := 2033;
        ELSIF x = 5796 THEN
            tanh_f := 2033;
        ELSIF x = 5797 THEN
            tanh_f := 2033;
        ELSIF x = 5798 THEN
            tanh_f := 2033;
        ELSIF x = 5799 THEN
            tanh_f := 2033;
        ELSIF x = 5800 THEN
            tanh_f := 2033;
        ELSIF x = 5801 THEN
            tanh_f := 2033;
        ELSIF x = 5802 THEN
            tanh_f := 2033;
        ELSIF x = 5803 THEN
            tanh_f := 2034;
        ELSIF x = 5804 THEN
            tanh_f := 2034;
        ELSIF x = 5805 THEN
            tanh_f := 2034;
        ELSIF x = 5806 THEN
            tanh_f := 2034;
        ELSIF x = 5807 THEN
            tanh_f := 2034;
        ELSIF x = 5808 THEN
            tanh_f := 2034;
        ELSIF x = 5809 THEN
            tanh_f := 2034;
        ELSIF x = 5810 THEN
            tanh_f := 2034;
        ELSIF x = 5811 THEN
            tanh_f := 2034;
        ELSIF x = 5812 THEN
            tanh_f := 2034;
        ELSIF x = 5813 THEN
            tanh_f := 2034;
        ELSIF x = 5814 THEN
            tanh_f := 2034;
        ELSIF x = 5815 THEN
            tanh_f := 2034;
        ELSIF x = 5816 THEN
            tanh_f := 2034;
        ELSIF x = 5817 THEN
            tanh_f := 2034;
        ELSIF x = 5818 THEN
            tanh_f := 2034;
        ELSIF x = 5819 THEN
            tanh_f := 2034;
        ELSIF x = 5820 THEN
            tanh_f := 2034;
        ELSIF x = 5821 THEN
            tanh_f := 2034;
        ELSIF x = 5822 THEN
            tanh_f := 2034;
        ELSIF x = 5823 THEN
            tanh_f := 2034;
        ELSIF x = 5824 THEN
            tanh_f := 2034;
        ELSIF x = 5825 THEN
            tanh_f := 2034;
        ELSIF x = 5826 THEN
            tanh_f := 2034;
        ELSIF x = 5827 THEN
            tanh_f := 2034;
        ELSIF x = 5828 THEN
            tanh_f := 2034;
        ELSIF x = 5829 THEN
            tanh_f := 2034;
        ELSIF x = 5830 THEN
            tanh_f := 2034;
        ELSIF x = 5831 THEN
            tanh_f := 2034;
        ELSIF x = 5832 THEN
            tanh_f := 2034;
        ELSIF x = 5833 THEN
            tanh_f := 2034;
        ELSIF x = 5834 THEN
            tanh_f := 2034;
        ELSIF x = 5835 THEN
            tanh_f := 2034;
        ELSIF x = 5836 THEN
            tanh_f := 2034;
        ELSIF x = 5837 THEN
            tanh_f := 2034;
        ELSIF x = 5838 THEN
            tanh_f := 2034;
        ELSIF x = 5839 THEN
            tanh_f := 2034;
        ELSIF x = 5840 THEN
            tanh_f := 2034;
        ELSIF x = 5841 THEN
            tanh_f := 2034;
        ELSIF x = 5842 THEN
            tanh_f := 2034;
        ELSIF x = 5843 THEN
            tanh_f := 2034;
        ELSIF x = 5844 THEN
            tanh_f := 2034;
        ELSIF x = 5845 THEN
            tanh_f := 2034;
        ELSIF x = 5846 THEN
            tanh_f := 2034;
        ELSIF x = 5847 THEN
            tanh_f := 2034;
        ELSIF x = 5848 THEN
            tanh_f := 2034;
        ELSIF x = 5849 THEN
            tanh_f := 2034;
        ELSIF x = 5850 THEN
            tanh_f := 2034;
        ELSIF x = 5851 THEN
            tanh_f := 2034;
        ELSIF x = 5852 THEN
            tanh_f := 2034;
        ELSIF x = 5853 THEN
            tanh_f := 2034;
        ELSIF x = 5854 THEN
            tanh_f := 2034;
        ELSIF x = 5855 THEN
            tanh_f := 2034;
        ELSIF x = 5856 THEN
            tanh_f := 2034;
        ELSIF x = 5857 THEN
            tanh_f := 2034;
        ELSIF x = 5858 THEN
            tanh_f := 2034;
        ELSIF x = 5859 THEN
            tanh_f := 2034;
        ELSIF x = 5860 THEN
            tanh_f := 2035;
        ELSIF x = 5861 THEN
            tanh_f := 2035;
        ELSIF x = 5862 THEN
            tanh_f := 2035;
        ELSIF x = 5863 THEN
            tanh_f := 2035;
        ELSIF x = 5864 THEN
            tanh_f := 2035;
        ELSIF x = 5865 THEN
            tanh_f := 2035;
        ELSIF x = 5866 THEN
            tanh_f := 2035;
        ELSIF x = 5867 THEN
            tanh_f := 2035;
        ELSIF x = 5868 THEN
            tanh_f := 2035;
        ELSIF x = 5869 THEN
            tanh_f := 2035;
        ELSIF x = 5870 THEN
            tanh_f := 2035;
        ELSIF x = 5871 THEN
            tanh_f := 2035;
        ELSIF x = 5872 THEN
            tanh_f := 2035;
        ELSIF x = 5873 THEN
            tanh_f := 2035;
        ELSIF x = 5874 THEN
            tanh_f := 2035;
        ELSIF x = 5875 THEN
            tanh_f := 2035;
        ELSIF x = 5876 THEN
            tanh_f := 2035;
        ELSIF x = 5877 THEN
            tanh_f := 2035;
        ELSIF x = 5878 THEN
            tanh_f := 2035;
        ELSIF x = 5879 THEN
            tanh_f := 2035;
        ELSIF x = 5880 THEN
            tanh_f := 2035;
        ELSIF x = 5881 THEN
            tanh_f := 2035;
        ELSIF x = 5882 THEN
            tanh_f := 2035;
        ELSIF x = 5883 THEN
            tanh_f := 2035;
        ELSIF x = 5884 THEN
            tanh_f := 2035;
        ELSIF x = 5885 THEN
            tanh_f := 2035;
        ELSIF x = 5886 THEN
            tanh_f := 2035;
        ELSIF x = 5887 THEN
            tanh_f := 2035;
        ELSIF x = 5888 THEN
            tanh_f := 2036;
        ELSIF x = 5889 THEN
            tanh_f := 2036;
        ELSIF x = 5890 THEN
            tanh_f := 2036;
        ELSIF x = 5891 THEN
            tanh_f := 2036;
        ELSIF x = 5892 THEN
            tanh_f := 2036;
        ELSIF x = 5893 THEN
            tanh_f := 2036;
        ELSIF x = 5894 THEN
            tanh_f := 2036;
        ELSIF x = 5895 THEN
            tanh_f := 2036;
        ELSIF x = 5896 THEN
            tanh_f := 2036;
        ELSIF x = 5897 THEN
            tanh_f := 2036;
        ELSIF x = 5898 THEN
            tanh_f := 2036;
        ELSIF x = 5899 THEN
            tanh_f := 2036;
        ELSIF x = 5900 THEN
            tanh_f := 2036;
        ELSIF x = 5901 THEN
            tanh_f := 2036;
        ELSIF x = 5902 THEN
            tanh_f := 2036;
        ELSIF x = 5903 THEN
            tanh_f := 2036;
        ELSIF x = 5904 THEN
            tanh_f := 2036;
        ELSIF x = 5905 THEN
            tanh_f := 2036;
        ELSIF x = 5906 THEN
            tanh_f := 2036;
        ELSIF x = 5907 THEN
            tanh_f := 2036;
        ELSIF x = 5908 THEN
            tanh_f := 2036;
        ELSIF x = 5909 THEN
            tanh_f := 2036;
        ELSIF x = 5910 THEN
            tanh_f := 2036;
        ELSIF x = 5911 THEN
            tanh_f := 2036;
        ELSIF x = 5912 THEN
            tanh_f := 2036;
        ELSIF x = 5913 THEN
            tanh_f := 2036;
        ELSIF x = 5914 THEN
            tanh_f := 2036;
        ELSIF x = 5915 THEN
            tanh_f := 2036;
        ELSIF x = 5916 THEN
            tanh_f := 2036;
        ELSIF x = 5917 THEN
            tanh_f := 2036;
        ELSIF x = 5918 THEN
            tanh_f := 2036;
        ELSIF x = 5919 THEN
            tanh_f := 2036;
        ELSIF x = 5920 THEN
            tanh_f := 2036;
        ELSIF x = 5921 THEN
            tanh_f := 2036;
        ELSIF x = 5922 THEN
            tanh_f := 2036;
        ELSIF x = 5923 THEN
            tanh_f := 2036;
        ELSIF x = 5924 THEN
            tanh_f := 2036;
        ELSIF x = 5925 THEN
            tanh_f := 2036;
        ELSIF x = 5926 THEN
            tanh_f := 2036;
        ELSIF x = 5927 THEN
            tanh_f := 2036;
        ELSIF x = 5928 THEN
            tanh_f := 2036;
        ELSIF x = 5929 THEN
            tanh_f := 2036;
        ELSIF x = 5930 THEN
            tanh_f := 2036;
        ELSIF x = 5931 THEN
            tanh_f := 2036;
        ELSIF x = 5932 THEN
            tanh_f := 2036;
        ELSIF x = 5933 THEN
            tanh_f := 2036;
        ELSIF x = 5934 THEN
            tanh_f := 2036;
        ELSIF x = 5935 THEN
            tanh_f := 2036;
        ELSIF x = 5936 THEN
            tanh_f := 2036;
        ELSIF x = 5937 THEN
            tanh_f := 2036;
        ELSIF x = 5938 THEN
            tanh_f := 2036;
        ELSIF x = 5939 THEN
            tanh_f := 2036;
        ELSIF x = 5940 THEN
            tanh_f := 2036;
        ELSIF x = 5941 THEN
            tanh_f := 2036;
        ELSIF x = 5942 THEN
            tanh_f := 2036;
        ELSIF x = 5943 THEN
            tanh_f := 2036;
        ELSIF x = 5944 THEN
            tanh_f := 2036;
        ELSIF x = 5945 THEN
            tanh_f := 2036;
        ELSIF x = 5946 THEN
            tanh_f := 2036;
        ELSIF x = 5947 THEN
            tanh_f := 2036;
        ELSIF x = 5948 THEN
            tanh_f := 2036;
        ELSIF x = 5949 THEN
            tanh_f := 2036;
        ELSIF x = 5950 THEN
            tanh_f := 2036;
        ELSIF x = 5951 THEN
            tanh_f := 2036;
        ELSIF x = 5952 THEN
            tanh_f := 2036;
        ELSIF x = 5953 THEN
            tanh_f := 2036;
        ELSIF x = 5954 THEN
            tanh_f := 2036;
        ELSIF x = 5955 THEN
            tanh_f := 2036;
        ELSIF x = 5956 THEN
            tanh_f := 2036;
        ELSIF x = 5957 THEN
            tanh_f := 2036;
        ELSIF x = 5958 THEN
            tanh_f := 2036;
        ELSIF x = 5959 THEN
            tanh_f := 2036;
        ELSIF x = 5960 THEN
            tanh_f := 2036;
        ELSIF x = 5961 THEN
            tanh_f := 2036;
        ELSIF x = 5962 THEN
            tanh_f := 2036;
        ELSIF x = 5963 THEN
            tanh_f := 2036;
        ELSIF x = 5964 THEN
            tanh_f := 2036;
        ELSIF x = 5965 THEN
            tanh_f := 2036;
        ELSIF x = 5966 THEN
            tanh_f := 2036;
        ELSIF x = 5967 THEN
            tanh_f := 2036;
        ELSIF x = 5968 THEN
            tanh_f := 2036;
        ELSIF x = 5969 THEN
            tanh_f := 2036;
        ELSIF x = 5970 THEN
            tanh_f := 2036;
        ELSIF x = 5971 THEN
            tanh_f := 2036;
        ELSIF x = 5972 THEN
            tanh_f := 2036;
        ELSIF x = 5973 THEN
            tanh_f := 2036;
        ELSIF x = 5974 THEN
            tanh_f := 2036;
        ELSIF x = 5975 THEN
            tanh_f := 2036;
        ELSIF x = 5976 THEN
            tanh_f := 2036;
        ELSIF x = 5977 THEN
            tanh_f := 2036;
        ELSIF x = 5978 THEN
            tanh_f := 2036;
        ELSIF x = 5979 THEN
            tanh_f := 2036;
        ELSIF x = 5980 THEN
            tanh_f := 2036;
        ELSIF x = 5981 THEN
            tanh_f := 2036;
        ELSIF x = 5982 THEN
            tanh_f := 2036;
        ELSIF x = 5983 THEN
            tanh_f := 2036;
        ELSIF x = 5984 THEN
            tanh_f := 2036;
        ELSIF x = 5985 THEN
            tanh_f := 2036;
        ELSIF x = 5986 THEN
            tanh_f := 2036;
        ELSIF x = 5987 THEN
            tanh_f := 2036;
        ELSIF x = 5988 THEN
            tanh_f := 2036;
        ELSIF x = 5989 THEN
            tanh_f := 2036;
        ELSIF x = 5990 THEN
            tanh_f := 2036;
        ELSIF x = 5991 THEN
            tanh_f := 2036;
        ELSIF x = 5992 THEN
            tanh_f := 2036;
        ELSIF x = 5993 THEN
            tanh_f := 2036;
        ELSIF x = 5994 THEN
            tanh_f := 2036;
        ELSIF x = 5995 THEN
            tanh_f := 2036;
        ELSIF x = 5996 THEN
            tanh_f := 2036;
        ELSIF x = 5997 THEN
            tanh_f := 2036;
        ELSIF x = 5998 THEN
            tanh_f := 2036;
        ELSIF x = 5999 THEN
            tanh_f := 2036;
        ELSIF x = 6000 THEN
            tanh_f := 2036;
        ELSIF x = 6001 THEN
            tanh_f := 2036;
        ELSIF x = 6002 THEN
            tanh_f := 2036;
        ELSIF x = 6003 THEN
            tanh_f := 2036;
        ELSIF x = 6004 THEN
            tanh_f := 2036;
        ELSIF x = 6005 THEN
            tanh_f := 2036;
        ELSIF x = 6006 THEN
            tanh_f := 2036;
        ELSIF x = 6007 THEN
            tanh_f := 2036;
        ELSIF x = 6008 THEN
            tanh_f := 2036;
        ELSIF x = 6009 THEN
            tanh_f := 2036;
        ELSIF x = 6010 THEN
            tanh_f := 2036;
        ELSIF x = 6011 THEN
            tanh_f := 2036;
        ELSIF x = 6012 THEN
            tanh_f := 2036;
        ELSIF x = 6013 THEN
            tanh_f := 2036;
        ELSIF x = 6014 THEN
            tanh_f := 2036;
        ELSIF x = 6015 THEN
            tanh_f := 2036;
        ELSIF x = 6016 THEN
            tanh_f := 2036;
        ELSIF x = 6017 THEN
            tanh_f := 2036;
        ELSIF x = 6018 THEN
            tanh_f := 2036;
        ELSIF x = 6019 THEN
            tanh_f := 2036;
        ELSIF x = 6020 THEN
            tanh_f := 2036;
        ELSIF x = 6021 THEN
            tanh_f := 2036;
        ELSIF x = 6022 THEN
            tanh_f := 2036;
        ELSIF x = 6023 THEN
            tanh_f := 2036;
        ELSIF x = 6024 THEN
            tanh_f := 2036;
        ELSIF x = 6025 THEN
            tanh_f := 2036;
        ELSIF x = 6026 THEN
            tanh_f := 2036;
        ELSIF x = 6027 THEN
            tanh_f := 2036;
        ELSIF x = 6028 THEN
            tanh_f := 2036;
        ELSIF x = 6029 THEN
            tanh_f := 2036;
        ELSIF x = 6030 THEN
            tanh_f := 2036;
        ELSIF x = 6031 THEN
            tanh_f := 2036;
        ELSIF x = 6032 THEN
            tanh_f := 2036;
        ELSIF x = 6033 THEN
            tanh_f := 2036;
        ELSIF x = 6034 THEN
            tanh_f := 2036;
        ELSIF x = 6035 THEN
            tanh_f := 2036;
        ELSIF x = 6036 THEN
            tanh_f := 2036;
        ELSIF x = 6037 THEN
            tanh_f := 2036;
        ELSIF x = 6038 THEN
            tanh_f := 2036;
        ELSIF x = 6039 THEN
            tanh_f := 2036;
        ELSIF x = 6040 THEN
            tanh_f := 2036;
        ELSIF x = 6041 THEN
            tanh_f := 2036;
        ELSIF x = 6042 THEN
            tanh_f := 2036;
        ELSIF x = 6043 THEN
            tanh_f := 2036;
        ELSIF x = 6044 THEN
            tanh_f := 2036;
        ELSIF x = 6045 THEN
            tanh_f := 2036;
        ELSIF x = 6046 THEN
            tanh_f := 2036;
        ELSIF x = 6047 THEN
            tanh_f := 2036;
        ELSIF x = 6048 THEN
            tanh_f := 2036;
        ELSIF x = 6049 THEN
            tanh_f := 2036;
        ELSIF x = 6050 THEN
            tanh_f := 2036;
        ELSIF x = 6051 THEN
            tanh_f := 2036;
        ELSIF x = 6052 THEN
            tanh_f := 2036;
        ELSIF x = 6053 THEN
            tanh_f := 2036;
        ELSIF x = 6054 THEN
            tanh_f := 2036;
        ELSIF x = 6055 THEN
            tanh_f := 2036;
        ELSIF x = 6056 THEN
            tanh_f := 2036;
        ELSIF x = 6057 THEN
            tanh_f := 2036;
        ELSIF x = 6058 THEN
            tanh_f := 2036;
        ELSIF x = 6059 THEN
            tanh_f := 2036;
        ELSIF x = 6060 THEN
            tanh_f := 2036;
        ELSIF x = 6061 THEN
            tanh_f := 2036;
        ELSIF x = 6062 THEN
            tanh_f := 2036;
        ELSIF x = 6063 THEN
            tanh_f := 2036;
        ELSIF x = 6064 THEN
            tanh_f := 2036;
        ELSIF x = 6065 THEN
            tanh_f := 2036;
        ELSIF x = 6066 THEN
            tanh_f := 2036;
        ELSIF x = 6067 THEN
            tanh_f := 2036;
        ELSIF x = 6068 THEN
            tanh_f := 2036;
        ELSIF x = 6069 THEN
            tanh_f := 2036;
        ELSIF x = 6070 THEN
            tanh_f := 2036;
        ELSIF x = 6071 THEN
            tanh_f := 2036;
        ELSIF x = 6072 THEN
            tanh_f := 2036;
        ELSIF x = 6073 THEN
            tanh_f := 2036;
        ELSIF x = 6074 THEN
            tanh_f := 2036;
        ELSIF x = 6075 THEN
            tanh_f := 2036;
        ELSIF x = 6076 THEN
            tanh_f := 2036;
        ELSIF x = 6077 THEN
            tanh_f := 2036;
        ELSIF x = 6078 THEN
            tanh_f := 2036;
        ELSIF x = 6079 THEN
            tanh_f := 2036;
        ELSIF x = 6080 THEN
            tanh_f := 2036;
        ELSIF x = 6081 THEN
            tanh_f := 2036;
        ELSIF x = 6082 THEN
            tanh_f := 2036;
        ELSIF x = 6083 THEN
            tanh_f := 2036;
        ELSIF x = 6084 THEN
            tanh_f := 2036;
        ELSIF x = 6085 THEN
            tanh_f := 2036;
        ELSIF x = 6086 THEN
            tanh_f := 2036;
        ELSIF x = 6087 THEN
            tanh_f := 2036;
        ELSIF x = 6088 THEN
            tanh_f := 2036;
        ELSIF x = 6089 THEN
            tanh_f := 2036;
        ELSIF x = 6090 THEN
            tanh_f := 2036;
        ELSIF x = 6091 THEN
            tanh_f := 2036;
        ELSIF x = 6092 THEN
            tanh_f := 2036;
        ELSIF x = 6093 THEN
            tanh_f := 2036;
        ELSIF x = 6094 THEN
            tanh_f := 2036;
        ELSIF x = 6095 THEN
            tanh_f := 2036;
        ELSIF x = 6096 THEN
            tanh_f := 2036;
        ELSIF x = 6097 THEN
            tanh_f := 2036;
        ELSIF x = 6098 THEN
            tanh_f := 2036;
        ELSIF x = 6099 THEN
            tanh_f := 2036;
        ELSIF x = 6100 THEN
            tanh_f := 2036;
        ELSIF x = 6101 THEN
            tanh_f := 2036;
        ELSIF x = 6102 THEN
            tanh_f := 2036;
        ELSIF x = 6103 THEN
            tanh_f := 2036;
        ELSIF x = 6104 THEN
            tanh_f := 2036;
        ELSIF x = 6105 THEN
            tanh_f := 2036;
        ELSIF x = 6106 THEN
            tanh_f := 2036;
        ELSIF x = 6107 THEN
            tanh_f := 2036;
        ELSIF x = 6108 THEN
            tanh_f := 2036;
        ELSIF x = 6109 THEN
            tanh_f := 2036;
        ELSIF x = 6110 THEN
            tanh_f := 2036;
        ELSIF x = 6111 THEN
            tanh_f := 2036;
        ELSIF x = 6112 THEN
            tanh_f := 2036;
        ELSIF x = 6113 THEN
            tanh_f := 2036;
        ELSIF x = 6114 THEN
            tanh_f := 2036;
        ELSIF x = 6115 THEN
            tanh_f := 2036;
        ELSIF x = 6116 THEN
            tanh_f := 2036;
        ELSIF x = 6117 THEN
            tanh_f := 2036;
        ELSIF x = 6118 THEN
            tanh_f := 2036;
        ELSIF x = 6119 THEN
            tanh_f := 2036;
        ELSIF x = 6120 THEN
            tanh_f := 2036;
        ELSIF x = 6121 THEN
            tanh_f := 2036;
        ELSIF x = 6122 THEN
            tanh_f := 2036;
        ELSIF x = 6123 THEN
            tanh_f := 2036;
        ELSIF x = 6124 THEN
            tanh_f := 2036;
        ELSIF x = 6125 THEN
            tanh_f := 2036;
        ELSIF x = 6126 THEN
            tanh_f := 2036;
        ELSIF x = 6127 THEN
            tanh_f := 2036;
        ELSIF x = 6128 THEN
            tanh_f := 2036;
        ELSIF x = 6129 THEN
            tanh_f := 2036;
        ELSIF x = 6130 THEN
            tanh_f := 2036;
        ELSIF x = 6131 THEN
            tanh_f := 2036;
        ELSIF x = 6132 THEN
            tanh_f := 2036;
        ELSIF x = 6133 THEN
            tanh_f := 2036;
        ELSIF x = 6134 THEN
            tanh_f := 2036;
        ELSIF x = 6135 THEN
            tanh_f := 2036;
        ELSIF x = 6136 THEN
            tanh_f := 2036;
        ELSIF x = 6137 THEN
            tanh_f := 2036;
        ELSIF x = 6138 THEN
            tanh_f := 2036;
        ELSIF x = 6139 THEN
            tanh_f := 2036;
        ELSIF x = 6140 THEN
            tanh_f := 2036;
        ELSIF x = 6141 THEN
            tanh_f := 2036;
        ELSIF x = 6142 THEN
            tanh_f := 2036;
        ELSIF x = 6143 THEN
            tanh_f := 2036;
        ELSIF x = 6144 THEN
            tanh_f := 2040;
        ELSIF x = 6145 THEN
            tanh_f := 2040;
        ELSIF x = 6146 THEN
            tanh_f := 2040;
        ELSIF x = 6147 THEN
            tanh_f := 2040;
        ELSIF x = 6148 THEN
            tanh_f := 2040;
        ELSIF x = 6149 THEN
            tanh_f := 2040;
        ELSIF x = 6150 THEN
            tanh_f := 2040;
        ELSIF x = 6151 THEN
            tanh_f := 2040;
        ELSIF x = 6152 THEN
            tanh_f := 2040;
        ELSIF x = 6153 THEN
            tanh_f := 2040;
        ELSIF x = 6154 THEN
            tanh_f := 2040;
        ELSIF x = 6155 THEN
            tanh_f := 2040;
        ELSIF x = 6156 THEN
            tanh_f := 2040;
        ELSIF x = 6157 THEN
            tanh_f := 2040;
        ELSIF x = 6158 THEN
            tanh_f := 2040;
        ELSIF x = 6159 THEN
            tanh_f := 2040;
        ELSIF x = 6160 THEN
            tanh_f := 2040;
        ELSIF x = 6161 THEN
            tanh_f := 2040;
        ELSIF x = 6162 THEN
            tanh_f := 2040;
        ELSIF x = 6163 THEN
            tanh_f := 2040;
        ELSIF x = 6164 THEN
            tanh_f := 2040;
        ELSIF x = 6165 THEN
            tanh_f := 2040;
        ELSIF x = 6166 THEN
            tanh_f := 2040;
        ELSIF x = 6167 THEN
            tanh_f := 2040;
        ELSIF x = 6168 THEN
            tanh_f := 2040;
        ELSIF x = 6169 THEN
            tanh_f := 2040;
        ELSIF x = 6170 THEN
            tanh_f := 2040;
        ELSIF x = 6171 THEN
            tanh_f := 2040;
        ELSIF x = 6172 THEN
            tanh_f := 2040;
        ELSIF x = 6173 THEN
            tanh_f := 2040;
        ELSIF x = 6174 THEN
            tanh_f := 2040;
        ELSIF x = 6175 THEN
            tanh_f := 2040;
        ELSIF x = 6176 THEN
            tanh_f := 2040;
        ELSIF x = 6177 THEN
            tanh_f := 2040;
        ELSIF x = 6178 THEN
            tanh_f := 2040;
        ELSIF x = 6179 THEN
            tanh_f := 2040;
        ELSIF x = 6180 THEN
            tanh_f := 2040;
        ELSIF x = 6181 THEN
            tanh_f := 2040;
        ELSIF x = 6182 THEN
            tanh_f := 2040;
        ELSIF x = 6183 THEN
            tanh_f := 2040;
        ELSIF x = 6184 THEN
            tanh_f := 2040;
        ELSIF x = 6185 THEN
            tanh_f := 2040;
        ELSIF x = 6186 THEN
            tanh_f := 2040;
        ELSIF x = 6187 THEN
            tanh_f := 2040;
        ELSIF x = 6188 THEN
            tanh_f := 2040;
        ELSIF x = 6189 THEN
            tanh_f := 2040;
        ELSIF x = 6190 THEN
            tanh_f := 2040;
        ELSIF x = 6191 THEN
            tanh_f := 2040;
        ELSIF x = 6192 THEN
            tanh_f := 2040;
        ELSIF x = 6193 THEN
            tanh_f := 2040;
        ELSIF x = 6194 THEN
            tanh_f := 2040;
        ELSIF x = 6195 THEN
            tanh_f := 2040;
        ELSIF x = 6196 THEN
            tanh_f := 2040;
        ELSIF x = 6197 THEN
            tanh_f := 2040;
        ELSIF x = 6198 THEN
            tanh_f := 2040;
        ELSIF x = 6199 THEN
            tanh_f := 2040;
        ELSIF x = 6200 THEN
            tanh_f := 2040;
        ELSIF x = 6201 THEN
            tanh_f := 2040;
        ELSIF x = 6202 THEN
            tanh_f := 2040;
        ELSIF x = 6203 THEN
            tanh_f := 2040;
        ELSIF x = 6204 THEN
            tanh_f := 2040;
        ELSIF x = 6205 THEN
            tanh_f := 2040;
        ELSIF x = 6206 THEN
            tanh_f := 2040;
        ELSIF x = 6207 THEN
            tanh_f := 2040;
        ELSIF x = 6208 THEN
            tanh_f := 2040;
        ELSIF x = 6209 THEN
            tanh_f := 2040;
        ELSIF x = 6210 THEN
            tanh_f := 2040;
        ELSIF x = 6211 THEN
            tanh_f := 2040;
        ELSIF x = 6212 THEN
            tanh_f := 2040;
        ELSIF x = 6213 THEN
            tanh_f := 2040;
        ELSIF x = 6214 THEN
            tanh_f := 2040;
        ELSIF x = 6215 THEN
            tanh_f := 2040;
        ELSIF x = 6216 THEN
            tanh_f := 2040;
        ELSIF x = 6217 THEN
            tanh_f := 2040;
        ELSIF x = 6218 THEN
            tanh_f := 2040;
        ELSIF x = 6219 THEN
            tanh_f := 2040;
        ELSIF x = 6220 THEN
            tanh_f := 2040;
        ELSIF x = 6221 THEN
            tanh_f := 2040;
        ELSIF x = 6222 THEN
            tanh_f := 2040;
        ELSIF x = 6223 THEN
            tanh_f := 2040;
        ELSIF x = 6224 THEN
            tanh_f := 2040;
        ELSIF x = 6225 THEN
            tanh_f := 2040;
        ELSIF x = 6226 THEN
            tanh_f := 2040;
        ELSIF x = 6227 THEN
            tanh_f := 2040;
        ELSIF x = 6228 THEN
            tanh_f := 2040;
        ELSIF x = 6229 THEN
            tanh_f := 2040;
        ELSIF x = 6230 THEN
            tanh_f := 2040;
        ELSIF x = 6231 THEN
            tanh_f := 2040;
        ELSIF x = 6232 THEN
            tanh_f := 2040;
        ELSIF x = 6233 THEN
            tanh_f := 2040;
        ELSIF x = 6234 THEN
            tanh_f := 2040;
        ELSIF x = 6235 THEN
            tanh_f := 2040;
        ELSIF x = 6236 THEN
            tanh_f := 2040;
        ELSIF x = 6237 THEN
            tanh_f := 2040;
        ELSIF x = 6238 THEN
            tanh_f := 2040;
        ELSIF x = 6239 THEN
            tanh_f := 2040;
        ELSIF x = 6240 THEN
            tanh_f := 2040;
        ELSIF x = 6241 THEN
            tanh_f := 2040;
        ELSIF x = 6242 THEN
            tanh_f := 2040;
        ELSIF x = 6243 THEN
            tanh_f := 2040;
        ELSIF x = 6244 THEN
            tanh_f := 2040;
        ELSIF x = 6245 THEN
            tanh_f := 2040;
        ELSIF x = 6246 THEN
            tanh_f := 2040;
        ELSIF x = 6247 THEN
            tanh_f := 2040;
        ELSIF x = 6248 THEN
            tanh_f := 2040;
        ELSIF x = 6249 THEN
            tanh_f := 2040;
        ELSIF x = 6250 THEN
            tanh_f := 2040;
        ELSIF x = 6251 THEN
            tanh_f := 2040;
        ELSIF x = 6252 THEN
            tanh_f := 2040;
        ELSIF x = 6253 THEN
            tanh_f := 2040;
        ELSIF x = 6254 THEN
            tanh_f := 2040;
        ELSIF x = 6255 THEN
            tanh_f := 2040;
        ELSIF x = 6256 THEN
            tanh_f := 2040;
        ELSIF x = 6257 THEN
            tanh_f := 2040;
        ELSIF x = 6258 THEN
            tanh_f := 2040;
        ELSIF x = 6259 THEN
            tanh_f := 2040;
        ELSIF x = 6260 THEN
            tanh_f := 2040;
        ELSIF x = 6261 THEN
            tanh_f := 2040;
        ELSIF x = 6262 THEN
            tanh_f := 2040;
        ELSIF x = 6263 THEN
            tanh_f := 2040;
        ELSIF x = 6264 THEN
            tanh_f := 2040;
        ELSIF x = 6265 THEN
            tanh_f := 2040;
        ELSIF x = 6266 THEN
            tanh_f := 2040;
        ELSIF x = 6267 THEN
            tanh_f := 2040;
        ELSIF x = 6268 THEN
            tanh_f := 2040;
        ELSIF x = 6269 THEN
            tanh_f := 2040;
        ELSIF x = 6270 THEN
            tanh_f := 2040;
        ELSIF x = 6271 THEN
            tanh_f := 2040;
        ELSIF x = 6272 THEN
            tanh_f := 2040;
        ELSIF x = 6273 THEN
            tanh_f := 2040;
        ELSIF x = 6274 THEN
            tanh_f := 2040;
        ELSIF x = 6275 THEN
            tanh_f := 2040;
        ELSIF x = 6276 THEN
            tanh_f := 2040;
        ELSIF x = 6277 THEN
            tanh_f := 2040;
        ELSIF x = 6278 THEN
            tanh_f := 2040;
        ELSIF x = 6279 THEN
            tanh_f := 2040;
        ELSIF x = 6280 THEN
            tanh_f := 2040;
        ELSIF x = 6281 THEN
            tanh_f := 2040;
        ELSIF x = 6282 THEN
            tanh_f := 2040;
        ELSIF x = 6283 THEN
            tanh_f := 2040;
        ELSIF x = 6284 THEN
            tanh_f := 2040;
        ELSIF x = 6285 THEN
            tanh_f := 2040;
        ELSIF x = 6286 THEN
            tanh_f := 2040;
        ELSIF x = 6287 THEN
            tanh_f := 2040;
        ELSIF x = 6288 THEN
            tanh_f := 2040;
        ELSIF x = 6289 THEN
            tanh_f := 2040;
        ELSIF x = 6290 THEN
            tanh_f := 2040;
        ELSIF x = 6291 THEN
            tanh_f := 2040;
        ELSIF x = 6292 THEN
            tanh_f := 2040;
        ELSIF x = 6293 THEN
            tanh_f := 2040;
        ELSIF x = 6294 THEN
            tanh_f := 2040;
        ELSIF x = 6295 THEN
            tanh_f := 2040;
        ELSIF x = 6296 THEN
            tanh_f := 2040;
        ELSIF x = 6297 THEN
            tanh_f := 2040;
        ELSIF x = 6298 THEN
            tanh_f := 2040;
        ELSIF x = 6299 THEN
            tanh_f := 2040;
        ELSIF x = 6300 THEN
            tanh_f := 2040;
        ELSIF x = 6301 THEN
            tanh_f := 2040;
        ELSIF x = 6302 THEN
            tanh_f := 2040;
        ELSIF x = 6303 THEN
            tanh_f := 2040;
        ELSIF x = 6304 THEN
            tanh_f := 2040;
        ELSIF x = 6305 THEN
            tanh_f := 2040;
        ELSIF x = 6306 THEN
            tanh_f := 2040;
        ELSIF x = 6307 THEN
            tanh_f := 2040;
        ELSIF x = 6308 THEN
            tanh_f := 2040;
        ELSIF x = 6309 THEN
            tanh_f := 2040;
        ELSIF x = 6310 THEN
            tanh_f := 2040;
        ELSIF x = 6311 THEN
            tanh_f := 2040;
        ELSIF x = 6312 THEN
            tanh_f := 2040;
        ELSIF x = 6313 THEN
            tanh_f := 2040;
        ELSIF x = 6314 THEN
            tanh_f := 2040;
        ELSIF x = 6315 THEN
            tanh_f := 2040;
        ELSIF x = 6316 THEN
            tanh_f := 2040;
        ELSIF x = 6317 THEN
            tanh_f := 2040;
        ELSIF x = 6318 THEN
            tanh_f := 2040;
        ELSIF x = 6319 THEN
            tanh_f := 2040;
        ELSIF x = 6320 THEN
            tanh_f := 2040;
        ELSIF x = 6321 THEN
            tanh_f := 2040;
        ELSIF x = 6322 THEN
            tanh_f := 2040;
        ELSIF x = 6323 THEN
            tanh_f := 2040;
        ELSIF x = 6324 THEN
            tanh_f := 2040;
        ELSIF x = 6325 THEN
            tanh_f := 2040;
        ELSIF x = 6326 THEN
            tanh_f := 2040;
        ELSIF x = 6327 THEN
            tanh_f := 2040;
        ELSIF x = 6328 THEN
            tanh_f := 2040;
        ELSIF x = 6329 THEN
            tanh_f := 2040;
        ELSIF x = 6330 THEN
            tanh_f := 2040;
        ELSIF x = 6331 THEN
            tanh_f := 2040;
        ELSIF x = 6332 THEN
            tanh_f := 2040;
        ELSIF x = 6333 THEN
            tanh_f := 2040;
        ELSIF x = 6334 THEN
            tanh_f := 2040;
        ELSIF x = 6335 THEN
            tanh_f := 2040;
        ELSIF x = 6336 THEN
            tanh_f := 2040;
        ELSIF x = 6337 THEN
            tanh_f := 2040;
        ELSIF x = 6338 THEN
            tanh_f := 2040;
        ELSIF x = 6339 THEN
            tanh_f := 2040;
        ELSIF x = 6340 THEN
            tanh_f := 2040;
        ELSIF x = 6341 THEN
            tanh_f := 2040;
        ELSIF x = 6342 THEN
            tanh_f := 2040;
        ELSIF x = 6343 THEN
            tanh_f := 2040;
        ELSIF x = 6344 THEN
            tanh_f := 2040;
        ELSIF x = 6345 THEN
            tanh_f := 2040;
        ELSIF x = 6346 THEN
            tanh_f := 2040;
        ELSIF x = 6347 THEN
            tanh_f := 2040;
        ELSIF x = 6348 THEN
            tanh_f := 2040;
        ELSIF x = 6349 THEN
            tanh_f := 2040;
        ELSIF x = 6350 THEN
            tanh_f := 2040;
        ELSIF x = 6351 THEN
            tanh_f := 2040;
        ELSIF x = 6352 THEN
            tanh_f := 2040;
        ELSIF x = 6353 THEN
            tanh_f := 2040;
        ELSIF x = 6354 THEN
            tanh_f := 2040;
        ELSIF x = 6355 THEN
            tanh_f := 2040;
        ELSIF x = 6356 THEN
            tanh_f := 2040;
        ELSIF x = 6357 THEN
            tanh_f := 2040;
        ELSIF x = 6358 THEN
            tanh_f := 2040;
        ELSIF x = 6359 THEN
            tanh_f := 2040;
        ELSIF x = 6360 THEN
            tanh_f := 2040;
        ELSIF x = 6361 THEN
            tanh_f := 2040;
        ELSIF x = 6362 THEN
            tanh_f := 2040;
        ELSIF x = 6363 THEN
            tanh_f := 2040;
        ELSIF x = 6364 THEN
            tanh_f := 2040;
        ELSIF x = 6365 THEN
            tanh_f := 2040;
        ELSIF x = 6366 THEN
            tanh_f := 2040;
        ELSIF x = 6367 THEN
            tanh_f := 2040;
        ELSIF x = 6368 THEN
            tanh_f := 2040;
        ELSIF x = 6369 THEN
            tanh_f := 2040;
        ELSIF x = 6370 THEN
            tanh_f := 2040;
        ELSIF x = 6371 THEN
            tanh_f := 2040;
        ELSIF x = 6372 THEN
            tanh_f := 2040;
        ELSIF x = 6373 THEN
            tanh_f := 2040;
        ELSIF x = 6374 THEN
            tanh_f := 2040;
        ELSIF x = 6375 THEN
            tanh_f := 2040;
        ELSIF x = 6376 THEN
            tanh_f := 2040;
        ELSIF x = 6377 THEN
            tanh_f := 2040;
        ELSIF x = 6378 THEN
            tanh_f := 2040;
        ELSIF x = 6379 THEN
            tanh_f := 2040;
        ELSIF x = 6380 THEN
            tanh_f := 2040;
        ELSIF x = 6381 THEN
            tanh_f := 2040;
        ELSIF x = 6382 THEN
            tanh_f := 2040;
        ELSIF x = 6383 THEN
            tanh_f := 2040;
        ELSIF x = 6384 THEN
            tanh_f := 2040;
        ELSIF x = 6385 THEN
            tanh_f := 2040;
        ELSIF x = 6386 THEN
            tanh_f := 2040;
        ELSIF x = 6387 THEN
            tanh_f := 2040;
        ELSIF x = 6388 THEN
            tanh_f := 2040;
        ELSIF x = 6389 THEN
            tanh_f := 2040;
        ELSIF x = 6390 THEN
            tanh_f := 2040;
        ELSIF x = 6391 THEN
            tanh_f := 2040;
        ELSIF x = 6392 THEN
            tanh_f := 2040;
        ELSIF x = 6393 THEN
            tanh_f := 2040;
        ELSIF x = 6394 THEN
            tanh_f := 2040;
        ELSIF x = 6395 THEN
            tanh_f := 2040;
        ELSIF x = 6396 THEN
            tanh_f := 2040;
        ELSIF x = 6397 THEN
            tanh_f := 2040;
        ELSIF x = 6398 THEN
            tanh_f := 2040;
        ELSIF x = 6399 THEN
            tanh_f := 2040;
        ELSIF x = 6400 THEN
            tanh_f := 2042;
        ELSIF x = 6401 THEN
            tanh_f := 2042;
        ELSIF x = 6402 THEN
            tanh_f := 2042;
        ELSIF x = 6403 THEN
            tanh_f := 2042;
        ELSIF x = 6404 THEN
            tanh_f := 2042;
        ELSIF x = 6405 THEN
            tanh_f := 2042;
        ELSIF x = 6406 THEN
            tanh_f := 2042;
        ELSIF x = 6407 THEN
            tanh_f := 2042;
        ELSIF x = 6408 THEN
            tanh_f := 2042;
        ELSIF x = 6409 THEN
            tanh_f := 2042;
        ELSIF x = 6410 THEN
            tanh_f := 2042;
        ELSIF x = 6411 THEN
            tanh_f := 2042;
        ELSIF x = 6412 THEN
            tanh_f := 2042;
        ELSIF x = 6413 THEN
            tanh_f := 2042;
        ELSIF x = 6414 THEN
            tanh_f := 2042;
        ELSIF x = 6415 THEN
            tanh_f := 2042;
        ELSIF x = 6416 THEN
            tanh_f := 2042;
        ELSIF x = 6417 THEN
            tanh_f := 2042;
        ELSIF x = 6418 THEN
            tanh_f := 2042;
        ELSIF x = 6419 THEN
            tanh_f := 2042;
        ELSIF x = 6420 THEN
            tanh_f := 2042;
        ELSIF x = 6421 THEN
            tanh_f := 2042;
        ELSIF x = 6422 THEN
            tanh_f := 2042;
        ELSIF x = 6423 THEN
            tanh_f := 2042;
        ELSIF x = 6424 THEN
            tanh_f := 2042;
        ELSIF x = 6425 THEN
            tanh_f := 2042;
        ELSIF x = 6426 THEN
            tanh_f := 2042;
        ELSIF x = 6427 THEN
            tanh_f := 2042;
        ELSIF x = 6428 THEN
            tanh_f := 2042;
        ELSIF x = 6429 THEN
            tanh_f := 2042;
        ELSIF x = 6430 THEN
            tanh_f := 2042;
        ELSIF x = 6431 THEN
            tanh_f := 2042;
        ELSIF x = 6432 THEN
            tanh_f := 2042;
        ELSIF x = 6433 THEN
            tanh_f := 2042;
        ELSIF x = 6434 THEN
            tanh_f := 2042;
        ELSIF x = 6435 THEN
            tanh_f := 2042;
        ELSIF x = 6436 THEN
            tanh_f := 2042;
        ELSIF x = 6437 THEN
            tanh_f := 2042;
        ELSIF x = 6438 THEN
            tanh_f := 2042;
        ELSIF x = 6439 THEN
            tanh_f := 2042;
        ELSIF x = 6440 THEN
            tanh_f := 2042;
        ELSIF x = 6441 THEN
            tanh_f := 2042;
        ELSIF x = 6442 THEN
            tanh_f := 2042;
        ELSIF x = 6443 THEN
            tanh_f := 2042;
        ELSIF x = 6444 THEN
            tanh_f := 2042;
        ELSIF x = 6445 THEN
            tanh_f := 2042;
        ELSIF x = 6446 THEN
            tanh_f := 2042;
        ELSIF x = 6447 THEN
            tanh_f := 2042;
        ELSIF x = 6448 THEN
            tanh_f := 2042;
        ELSIF x = 6449 THEN
            tanh_f := 2042;
        ELSIF x = 6450 THEN
            tanh_f := 2042;
        ELSIF x = 6451 THEN
            tanh_f := 2042;
        ELSIF x = 6452 THEN
            tanh_f := 2042;
        ELSIF x = 6453 THEN
            tanh_f := 2042;
        ELSIF x = 6454 THEN
            tanh_f := 2042;
        ELSIF x = 6455 THEN
            tanh_f := 2042;
        ELSIF x = 6456 THEN
            tanh_f := 2042;
        ELSIF x = 6457 THEN
            tanh_f := 2042;
        ELSIF x = 6458 THEN
            tanh_f := 2042;
        ELSIF x = 6459 THEN
            tanh_f := 2042;
        ELSIF x = 6460 THEN
            tanh_f := 2042;
        ELSIF x = 6461 THEN
            tanh_f := 2042;
        ELSIF x = 6462 THEN
            tanh_f := 2042;
        ELSIF x = 6463 THEN
            tanh_f := 2042;
        ELSIF x = 6464 THEN
            tanh_f := 2042;
        ELSIF x = 6465 THEN
            tanh_f := 2042;
        ELSIF x = 6466 THEN
            tanh_f := 2042;
        ELSIF x = 6467 THEN
            tanh_f := 2042;
        ELSIF x = 6468 THEN
            tanh_f := 2042;
        ELSIF x = 6469 THEN
            tanh_f := 2042;
        ELSIF x = 6470 THEN
            tanh_f := 2042;
        ELSIF x = 6471 THEN
            tanh_f := 2042;
        ELSIF x = 6472 THEN
            tanh_f := 2042;
        ELSIF x = 6473 THEN
            tanh_f := 2042;
        ELSIF x = 6474 THEN
            tanh_f := 2042;
        ELSIF x = 6475 THEN
            tanh_f := 2042;
        ELSIF x = 6476 THEN
            tanh_f := 2042;
        ELSIF x = 6477 THEN
            tanh_f := 2042;
        ELSIF x = 6478 THEN
            tanh_f := 2042;
        ELSIF x = 6479 THEN
            tanh_f := 2042;
        ELSIF x = 6480 THEN
            tanh_f := 2042;
        ELSIF x = 6481 THEN
            tanh_f := 2042;
        ELSIF x = 6482 THEN
            tanh_f := 2042;
        ELSIF x = 6483 THEN
            tanh_f := 2042;
        ELSIF x = 6484 THEN
            tanh_f := 2042;
        ELSIF x = 6485 THEN
            tanh_f := 2042;
        ELSIF x = 6486 THEN
            tanh_f := 2042;
        ELSIF x = 6487 THEN
            tanh_f := 2042;
        ELSIF x = 6488 THEN
            tanh_f := 2042;
        ELSIF x = 6489 THEN
            tanh_f := 2042;
        ELSIF x = 6490 THEN
            tanh_f := 2042;
        ELSIF x = 6491 THEN
            tanh_f := 2042;
        ELSIF x = 6492 THEN
            tanh_f := 2042;
        ELSIF x = 6493 THEN
            tanh_f := 2042;
        ELSIF x = 6494 THEN
            tanh_f := 2042;
        ELSIF x = 6495 THEN
            tanh_f := 2042;
        ELSIF x = 6496 THEN
            tanh_f := 2042;
        ELSIF x = 6497 THEN
            tanh_f := 2042;
        ELSIF x = 6498 THEN
            tanh_f := 2042;
        ELSIF x = 6499 THEN
            tanh_f := 2042;
        ELSIF x = 6500 THEN
            tanh_f := 2042;
        ELSIF x = 6501 THEN
            tanh_f := 2042;
        ELSIF x = 6502 THEN
            tanh_f := 2042;
        ELSIF x = 6503 THEN
            tanh_f := 2042;
        ELSIF x = 6504 THEN
            tanh_f := 2042;
        ELSIF x = 6505 THEN
            tanh_f := 2042;
        ELSIF x = 6506 THEN
            tanh_f := 2042;
        ELSIF x = 6507 THEN
            tanh_f := 2042;
        ELSIF x = 6508 THEN
            tanh_f := 2042;
        ELSIF x = 6509 THEN
            tanh_f := 2042;
        ELSIF x = 6510 THEN
            tanh_f := 2042;
        ELSIF x = 6511 THEN
            tanh_f := 2042;
        ELSIF x = 6512 THEN
            tanh_f := 2042;
        ELSIF x = 6513 THEN
            tanh_f := 2042;
        ELSIF x = 6514 THEN
            tanh_f := 2042;
        ELSIF x = 6515 THEN
            tanh_f := 2042;
        ELSIF x = 6516 THEN
            tanh_f := 2042;
        ELSIF x = 6517 THEN
            tanh_f := 2042;
        ELSIF x = 6518 THEN
            tanh_f := 2042;
        ELSIF x = 6519 THEN
            tanh_f := 2042;
        ELSIF x = 6520 THEN
            tanh_f := 2042;
        ELSIF x = 6521 THEN
            tanh_f := 2042;
        ELSIF x = 6522 THEN
            tanh_f := 2042;
        ELSIF x = 6523 THEN
            tanh_f := 2042;
        ELSIF x = 6524 THEN
            tanh_f := 2042;
        ELSIF x = 6525 THEN
            tanh_f := 2042;
        ELSIF x = 6526 THEN
            tanh_f := 2042;
        ELSIF x = 6527 THEN
            tanh_f := 2042;
        ELSIF x = 6528 THEN
            tanh_f := 2042;
        ELSIF x = 6529 THEN
            tanh_f := 2042;
        ELSIF x = 6530 THEN
            tanh_f := 2042;
        ELSIF x = 6531 THEN
            tanh_f := 2042;
        ELSIF x = 6532 THEN
            tanh_f := 2042;
        ELSIF x = 6533 THEN
            tanh_f := 2042;
        ELSIF x = 6534 THEN
            tanh_f := 2042;
        ELSIF x = 6535 THEN
            tanh_f := 2042;
        ELSIF x = 6536 THEN
            tanh_f := 2042;
        ELSIF x = 6537 THEN
            tanh_f := 2042;
        ELSIF x = 6538 THEN
            tanh_f := 2042;
        ELSIF x = 6539 THEN
            tanh_f := 2042;
        ELSIF x = 6540 THEN
            tanh_f := 2042;
        ELSIF x = 6541 THEN
            tanh_f := 2042;
        ELSIF x = 6542 THEN
            tanh_f := 2042;
        ELSIF x = 6543 THEN
            tanh_f := 2042;
        ELSIF x = 6544 THEN
            tanh_f := 2042;
        ELSIF x = 6545 THEN
            tanh_f := 2042;
        ELSIF x = 6546 THEN
            tanh_f := 2042;
        ELSIF x = 6547 THEN
            tanh_f := 2042;
        ELSIF x = 6548 THEN
            tanh_f := 2042;
        ELSIF x = 6549 THEN
            tanh_f := 2042;
        ELSIF x = 6550 THEN
            tanh_f := 2042;
        ELSIF x = 6551 THEN
            tanh_f := 2042;
        ELSIF x = 6552 THEN
            tanh_f := 2042;
        ELSIF x = 6553 THEN
            tanh_f := 2042;
        ELSIF x = 6554 THEN
            tanh_f := 2042;
        ELSIF x = 6555 THEN
            tanh_f := 2042;
        ELSIF x = 6556 THEN
            tanh_f := 2042;
        ELSIF x = 6557 THEN
            tanh_f := 2042;
        ELSIF x = 6558 THEN
            tanh_f := 2042;
        ELSIF x = 6559 THEN
            tanh_f := 2042;
        ELSIF x = 6560 THEN
            tanh_f := 2042;
        ELSIF x = 6561 THEN
            tanh_f := 2042;
        ELSIF x = 6562 THEN
            tanh_f := 2042;
        ELSIF x = 6563 THEN
            tanh_f := 2042;
        ELSIF x = 6564 THEN
            tanh_f := 2042;
        ELSIF x = 6565 THEN
            tanh_f := 2042;
        ELSIF x = 6566 THEN
            tanh_f := 2042;
        ELSIF x = 6567 THEN
            tanh_f := 2042;
        ELSIF x = 6568 THEN
            tanh_f := 2042;
        ELSIF x = 6569 THEN
            tanh_f := 2042;
        ELSIF x = 6570 THEN
            tanh_f := 2042;
        ELSIF x = 6571 THEN
            tanh_f := 2042;
        ELSIF x = 6572 THEN
            tanh_f := 2042;
        ELSIF x = 6573 THEN
            tanh_f := 2042;
        ELSIF x = 6574 THEN
            tanh_f := 2042;
        ELSIF x = 6575 THEN
            tanh_f := 2042;
        ELSIF x = 6576 THEN
            tanh_f := 2042;
        ELSIF x = 6577 THEN
            tanh_f := 2042;
        ELSIF x = 6578 THEN
            tanh_f := 2042;
        ELSIF x = 6579 THEN
            tanh_f := 2042;
        ELSIF x = 6580 THEN
            tanh_f := 2042;
        ELSIF x = 6581 THEN
            tanh_f := 2042;
        ELSIF x = 6582 THEN
            tanh_f := 2042;
        ELSIF x = 6583 THEN
            tanh_f := 2042;
        ELSIF x = 6584 THEN
            tanh_f := 2042;
        ELSIF x = 6585 THEN
            tanh_f := 2042;
        ELSIF x = 6586 THEN
            tanh_f := 2042;
        ELSIF x = 6587 THEN
            tanh_f := 2042;
        ELSIF x = 6588 THEN
            tanh_f := 2042;
        ELSIF x = 6589 THEN
            tanh_f := 2042;
        ELSIF x = 6590 THEN
            tanh_f := 2042;
        ELSIF x = 6591 THEN
            tanh_f := 2042;
        ELSIF x = 6592 THEN
            tanh_f := 2042;
        ELSIF x = 6593 THEN
            tanh_f := 2042;
        ELSIF x = 6594 THEN
            tanh_f := 2042;
        ELSIF x = 6595 THEN
            tanh_f := 2042;
        ELSIF x = 6596 THEN
            tanh_f := 2042;
        ELSIF x = 6597 THEN
            tanh_f := 2042;
        ELSIF x = 6598 THEN
            tanh_f := 2042;
        ELSIF x = 6599 THEN
            tanh_f := 2042;
        ELSIF x = 6600 THEN
            tanh_f := 2042;
        ELSIF x = 6601 THEN
            tanh_f := 2042;
        ELSIF x = 6602 THEN
            tanh_f := 2042;
        ELSIF x = 6603 THEN
            tanh_f := 2042;
        ELSIF x = 6604 THEN
            tanh_f := 2042;
        ELSIF x = 6605 THEN
            tanh_f := 2042;
        ELSIF x = 6606 THEN
            tanh_f := 2042;
        ELSIF x = 6607 THEN
            tanh_f := 2042;
        ELSIF x = 6608 THEN
            tanh_f := 2042;
        ELSIF x = 6609 THEN
            tanh_f := 2042;
        ELSIF x = 6610 THEN
            tanh_f := 2042;
        ELSIF x = 6611 THEN
            tanh_f := 2042;
        ELSIF x = 6612 THEN
            tanh_f := 2042;
        ELSIF x = 6613 THEN
            tanh_f := 2042;
        ELSIF x = 6614 THEN
            tanh_f := 2042;
        ELSIF x = 6615 THEN
            tanh_f := 2042;
        ELSIF x = 6616 THEN
            tanh_f := 2042;
        ELSIF x = 6617 THEN
            tanh_f := 2042;
        ELSIF x = 6618 THEN
            tanh_f := 2042;
        ELSIF x = 6619 THEN
            tanh_f := 2042;
        ELSIF x = 6620 THEN
            tanh_f := 2042;
        ELSIF x = 6621 THEN
            tanh_f := 2042;
        ELSIF x = 6622 THEN
            tanh_f := 2042;
        ELSIF x = 6623 THEN
            tanh_f := 2042;
        ELSIF x = 6624 THEN
            tanh_f := 2042;
        ELSIF x = 6625 THEN
            tanh_f := 2042;
        ELSIF x = 6626 THEN
            tanh_f := 2042;
        ELSIF x = 6627 THEN
            tanh_f := 2042;
        ELSIF x = 6628 THEN
            tanh_f := 2042;
        ELSIF x = 6629 THEN
            tanh_f := 2042;
        ELSIF x = 6630 THEN
            tanh_f := 2042;
        ELSIF x = 6631 THEN
            tanh_f := 2042;
        ELSIF x = 6632 THEN
            tanh_f := 2042;
        ELSIF x = 6633 THEN
            tanh_f := 2042;
        ELSIF x = 6634 THEN
            tanh_f := 2042;
        ELSIF x = 6635 THEN
            tanh_f := 2042;
        ELSIF x = 6636 THEN
            tanh_f := 2042;
        ELSIF x = 6637 THEN
            tanh_f := 2042;
        ELSIF x = 6638 THEN
            tanh_f := 2042;
        ELSIF x = 6639 THEN
            tanh_f := 2042;
        ELSIF x = 6640 THEN
            tanh_f := 2042;
        ELSIF x = 6641 THEN
            tanh_f := 2042;
        ELSIF x = 6642 THEN
            tanh_f := 2042;
        ELSIF x = 6643 THEN
            tanh_f := 2042;
        ELSIF x = 6644 THEN
            tanh_f := 2042;
        ELSIF x = 6645 THEN
            tanh_f := 2042;
        ELSIF x = 6646 THEN
            tanh_f := 2042;
        ELSIF x = 6647 THEN
            tanh_f := 2042;
        ELSIF x = 6648 THEN
            tanh_f := 2042;
        ELSIF x = 6649 THEN
            tanh_f := 2042;
        ELSIF x = 6650 THEN
            tanh_f := 2042;
        ELSIF x = 6651 THEN
            tanh_f := 2042;
        ELSIF x = 6652 THEN
            tanh_f := 2042;
        ELSIF x = 6653 THEN
            tanh_f := 2042;
        ELSIF x = 6654 THEN
            tanh_f := 2042;
        ELSIF x = 6655 THEN
            tanh_f := 2042;
        ELSIF x = 6656 THEN
            tanh_f := 2042;
        ELSIF x = 6657 THEN
            tanh_f := 2042;
        ELSIF x = 6658 THEN
            tanh_f := 2042;
        ELSIF x = 6659 THEN
            tanh_f := 2042;
        ELSIF x = 6660 THEN
            tanh_f := 2042;
        ELSIF x = 6661 THEN
            tanh_f := 2042;
        ELSIF x = 6662 THEN
            tanh_f := 2042;
        ELSIF x = 6663 THEN
            tanh_f := 2042;
        ELSIF x = 6664 THEN
            tanh_f := 2042;
        ELSIF x = 6665 THEN
            tanh_f := 2042;
        ELSIF x = 6666 THEN
            tanh_f := 2042;
        ELSIF x = 6667 THEN
            tanh_f := 2042;
        ELSIF x = 6668 THEN
            tanh_f := 2042;
        ELSIF x = 6669 THEN
            tanh_f := 2042;
        ELSIF x = 6670 THEN
            tanh_f := 2042;
        ELSIF x = 6671 THEN
            tanh_f := 2042;
        ELSIF x = 6672 THEN
            tanh_f := 2042;
        ELSIF x = 6673 THEN
            tanh_f := 2042;
        ELSIF x = 6674 THEN
            tanh_f := 2042;
        ELSIF x = 6675 THEN
            tanh_f := 2042;
        ELSIF x = 6676 THEN
            tanh_f := 2042;
        ELSIF x = 6677 THEN
            tanh_f := 2042;
        ELSIF x = 6678 THEN
            tanh_f := 2042;
        ELSIF x = 6679 THEN
            tanh_f := 2042;
        ELSIF x = 6680 THEN
            tanh_f := 2042;
        ELSIF x = 6681 THEN
            tanh_f := 2042;
        ELSIF x = 6682 THEN
            tanh_f := 2042;
        ELSIF x = 6683 THEN
            tanh_f := 2042;
        ELSIF x = 6684 THEN
            tanh_f := 2042;
        ELSIF x = 6685 THEN
            tanh_f := 2042;
        ELSIF x = 6686 THEN
            tanh_f := 2042;
        ELSIF x = 6687 THEN
            tanh_f := 2042;
        ELSIF x = 6688 THEN
            tanh_f := 2042;
        ELSIF x = 6689 THEN
            tanh_f := 2042;
        ELSIF x = 6690 THEN
            tanh_f := 2042;
        ELSIF x = 6691 THEN
            tanh_f := 2042;
        ELSIF x = 6692 THEN
            tanh_f := 2042;
        ELSIF x = 6693 THEN
            tanh_f := 2042;
        ELSIF x = 6694 THEN
            tanh_f := 2042;
        ELSIF x = 6695 THEN
            tanh_f := 2042;
        ELSIF x = 6696 THEN
            tanh_f := 2042;
        ELSIF x = 6697 THEN
            tanh_f := 2042;
        ELSIF x = 6698 THEN
            tanh_f := 2042;
        ELSIF x = 6699 THEN
            tanh_f := 2042;
        ELSIF x = 6700 THEN
            tanh_f := 2042;
        ELSIF x = 6701 THEN
            tanh_f := 2042;
        ELSIF x = 6702 THEN
            tanh_f := 2042;
        ELSIF x = 6703 THEN
            tanh_f := 2042;
        ELSIF x = 6704 THEN
            tanh_f := 2042;
        ELSIF x = 6705 THEN
            tanh_f := 2042;
        ELSIF x = 6706 THEN
            tanh_f := 2042;
        ELSIF x = 6707 THEN
            tanh_f := 2042;
        ELSIF x = 6708 THEN
            tanh_f := 2042;
        ELSIF x = 6709 THEN
            tanh_f := 2042;
        ELSIF x = 6710 THEN
            tanh_f := 2042;
        ELSIF x = 6711 THEN
            tanh_f := 2042;
        ELSIF x = 6712 THEN
            tanh_f := 2042;
        ELSIF x = 6713 THEN
            tanh_f := 2042;
        ELSIF x = 6714 THEN
            tanh_f := 2042;
        ELSIF x = 6715 THEN
            tanh_f := 2042;
        ELSIF x = 6716 THEN
            tanh_f := 2042;
        ELSIF x = 6717 THEN
            tanh_f := 2042;
        ELSIF x = 6718 THEN
            tanh_f := 2042;
        ELSIF x = 6719 THEN
            tanh_f := 2042;
        ELSIF x = 6720 THEN
            tanh_f := 2042;
        ELSIF x = 6721 THEN
            tanh_f := 2042;
        ELSIF x = 6722 THEN
            tanh_f := 2042;
        ELSIF x = 6723 THEN
            tanh_f := 2042;
        ELSIF x = 6724 THEN
            tanh_f := 2042;
        ELSIF x = 6725 THEN
            tanh_f := 2042;
        ELSIF x = 6726 THEN
            tanh_f := 2042;
        ELSIF x = 6727 THEN
            tanh_f := 2042;
        ELSIF x = 6728 THEN
            tanh_f := 2042;
        ELSIF x = 6729 THEN
            tanh_f := 2042;
        ELSIF x = 6730 THEN
            tanh_f := 2042;
        ELSIF x = 6731 THEN
            tanh_f := 2042;
        ELSIF x = 6732 THEN
            tanh_f := 2042;
        ELSIF x = 6733 THEN
            tanh_f := 2042;
        ELSIF x = 6734 THEN
            tanh_f := 2042;
        ELSIF x = 6735 THEN
            tanh_f := 2042;
        ELSIF x = 6736 THEN
            tanh_f := 2042;
        ELSIF x = 6737 THEN
            tanh_f := 2042;
        ELSIF x = 6738 THEN
            tanh_f := 2042;
        ELSIF x = 6739 THEN
            tanh_f := 2042;
        ELSIF x = 6740 THEN
            tanh_f := 2042;
        ELSIF x = 6741 THEN
            tanh_f := 2042;
        ELSIF x = 6742 THEN
            tanh_f := 2042;
        ELSIF x = 6743 THEN
            tanh_f := 2042;
        ELSIF x = 6744 THEN
            tanh_f := 2042;
        ELSIF x = 6745 THEN
            tanh_f := 2042;
        ELSIF x = 6746 THEN
            tanh_f := 2042;
        ELSIF x = 6747 THEN
            tanh_f := 2042;
        ELSIF x = 6748 THEN
            tanh_f := 2042;
        ELSIF x = 6749 THEN
            tanh_f := 2042;
        ELSIF x = 6750 THEN
            tanh_f := 2042;
        ELSIF x = 6751 THEN
            tanh_f := 2042;
        ELSIF x = 6752 THEN
            tanh_f := 2042;
        ELSIF x = 6753 THEN
            tanh_f := 2042;
        ELSIF x = 6754 THEN
            tanh_f := 2042;
        ELSIF x = 6755 THEN
            tanh_f := 2042;
        ELSIF x = 6756 THEN
            tanh_f := 2042;
        ELSIF x = 6757 THEN
            tanh_f := 2042;
        ELSIF x = 6758 THEN
            tanh_f := 2042;
        ELSIF x = 6759 THEN
            tanh_f := 2042;
        ELSIF x = 6760 THEN
            tanh_f := 2042;
        ELSIF x = 6761 THEN
            tanh_f := 2042;
        ELSIF x = 6762 THEN
            tanh_f := 2042;
        ELSIF x = 6763 THEN
            tanh_f := 2042;
        ELSIF x = 6764 THEN
            tanh_f := 2042;
        ELSIF x = 6765 THEN
            tanh_f := 2042;
        ELSIF x = 6766 THEN
            tanh_f := 2042;
        ELSIF x = 6767 THEN
            tanh_f := 2042;
        ELSIF x = 6768 THEN
            tanh_f := 2042;
        ELSIF x = 6769 THEN
            tanh_f := 2042;
        ELSIF x = 6770 THEN
            tanh_f := 2042;
        ELSIF x = 6771 THEN
            tanh_f := 2042;
        ELSIF x = 6772 THEN
            tanh_f := 2042;
        ELSIF x = 6773 THEN
            tanh_f := 2042;
        ELSIF x = 6774 THEN
            tanh_f := 2042;
        ELSIF x = 6775 THEN
            tanh_f := 2042;
        ELSIF x = 6776 THEN
            tanh_f := 2042;
        ELSIF x = 6777 THEN
            tanh_f := 2042;
        ELSIF x = 6778 THEN
            tanh_f := 2042;
        ELSIF x = 6779 THEN
            tanh_f := 2042;
        ELSIF x = 6780 THEN
            tanh_f := 2042;
        ELSIF x = 6781 THEN
            tanh_f := 2042;
        ELSIF x = 6782 THEN
            tanh_f := 2042;
        ELSIF x = 6783 THEN
            tanh_f := 2042;
        ELSIF x = 6784 THEN
            tanh_f := 2042;
        ELSIF x = 6785 THEN
            tanh_f := 2042;
        ELSIF x = 6786 THEN
            tanh_f := 2042;
        ELSIF x = 6787 THEN
            tanh_f := 2042;
        ELSIF x = 6788 THEN
            tanh_f := 2042;
        ELSIF x = 6789 THEN
            tanh_f := 2042;
        ELSIF x = 6790 THEN
            tanh_f := 2042;
        ELSIF x = 6791 THEN
            tanh_f := 2042;
        ELSIF x = 6792 THEN
            tanh_f := 2042;
        ELSIF x = 6793 THEN
            tanh_f := 2042;
        ELSIF x = 6794 THEN
            tanh_f := 2042;
        ELSIF x = 6795 THEN
            tanh_f := 2042;
        ELSIF x = 6796 THEN
            tanh_f := 2042;
        ELSIF x = 6797 THEN
            tanh_f := 2042;
        ELSIF x = 6798 THEN
            tanh_f := 2042;
        ELSIF x = 6799 THEN
            tanh_f := 2042;
        ELSIF x = 6800 THEN
            tanh_f := 2042;
        ELSIF x = 6801 THEN
            tanh_f := 2042;
        ELSIF x = 6802 THEN
            tanh_f := 2042;
        ELSIF x = 6803 THEN
            tanh_f := 2042;
        ELSIF x = 6804 THEN
            tanh_f := 2042;
        ELSIF x = 6805 THEN
            tanh_f := 2042;
        ELSIF x = 6806 THEN
            tanh_f := 2042;
        ELSIF x = 6807 THEN
            tanh_f := 2042;
        ELSIF x = 6808 THEN
            tanh_f := 2042;
        ELSIF x = 6809 THEN
            tanh_f := 2042;
        ELSIF x = 6810 THEN
            tanh_f := 2042;
        ELSIF x = 6811 THEN
            tanh_f := 2042;
        ELSIF x = 6812 THEN
            tanh_f := 2042;
        ELSIF x = 6813 THEN
            tanh_f := 2042;
        ELSIF x = 6814 THEN
            tanh_f := 2042;
        ELSIF x = 6815 THEN
            tanh_f := 2042;
        ELSIF x = 6816 THEN
            tanh_f := 2042;
        ELSIF x = 6817 THEN
            tanh_f := 2042;
        ELSIF x = 6818 THEN
            tanh_f := 2042;
        ELSIF x = 6819 THEN
            tanh_f := 2042;
        ELSIF x = 6820 THEN
            tanh_f := 2042;
        ELSIF x = 6821 THEN
            tanh_f := 2042;
        ELSIF x = 6822 THEN
            tanh_f := 2042;
        ELSIF x = 6823 THEN
            tanh_f := 2042;
        ELSIF x = 6824 THEN
            tanh_f := 2042;
        ELSIF x = 6825 THEN
            tanh_f := 2042;
        ELSIF x = 6826 THEN
            tanh_f := 2042;
        ELSIF x = 6827 THEN
            tanh_f := 2042;
        ELSIF x = 6828 THEN
            tanh_f := 2042;
        ELSIF x = 6829 THEN
            tanh_f := 2042;
        ELSIF x = 6830 THEN
            tanh_f := 2042;
        ELSIF x = 6831 THEN
            tanh_f := 2042;
        ELSIF x = 6832 THEN
            tanh_f := 2042;
        ELSIF x = 6833 THEN
            tanh_f := 2042;
        ELSIF x = 6834 THEN
            tanh_f := 2042;
        ELSIF x = 6835 THEN
            tanh_f := 2042;
        ELSIF x = 6836 THEN
            tanh_f := 2042;
        ELSIF x = 6837 THEN
            tanh_f := 2042;
        ELSIF x = 6838 THEN
            tanh_f := 2042;
        ELSIF x = 6839 THEN
            tanh_f := 2042;
        ELSIF x = 6840 THEN
            tanh_f := 2042;
        ELSIF x = 6841 THEN
            tanh_f := 2042;
        ELSIF x = 6842 THEN
            tanh_f := 2042;
        ELSIF x = 6843 THEN
            tanh_f := 2042;
        ELSIF x = 6844 THEN
            tanh_f := 2042;
        ELSIF x = 6845 THEN
            tanh_f := 2042;
        ELSIF x = 6846 THEN
            tanh_f := 2042;
        ELSIF x = 6847 THEN
            tanh_f := 2042;
        ELSIF x = 6848 THEN
            tanh_f := 2042;
        ELSIF x = 6849 THEN
            tanh_f := 2042;
        ELSIF x = 6850 THEN
            tanh_f := 2042;
        ELSIF x = 6851 THEN
            tanh_f := 2042;
        ELSIF x = 6852 THEN
            tanh_f := 2042;
        ELSIF x = 6853 THEN
            tanh_f := 2042;
        ELSIF x = 6854 THEN
            tanh_f := 2042;
        ELSIF x = 6855 THEN
            tanh_f := 2042;
        ELSIF x = 6856 THEN
            tanh_f := 2042;
        ELSIF x = 6857 THEN
            tanh_f := 2042;
        ELSIF x = 6858 THEN
            tanh_f := 2042;
        ELSIF x = 6859 THEN
            tanh_f := 2042;
        ELSIF x = 6860 THEN
            tanh_f := 2042;
        ELSIF x = 6861 THEN
            tanh_f := 2042;
        ELSIF x = 6862 THEN
            tanh_f := 2042;
        ELSIF x = 6863 THEN
            tanh_f := 2042;
        ELSIF x = 6864 THEN
            tanh_f := 2042;
        ELSIF x = 6865 THEN
            tanh_f := 2042;
        ELSIF x = 6866 THEN
            tanh_f := 2042;
        ELSIF x = 6867 THEN
            tanh_f := 2042;
        ELSIF x = 6868 THEN
            tanh_f := 2042;
        ELSIF x = 6869 THEN
            tanh_f := 2042;
        ELSIF x = 6870 THEN
            tanh_f := 2042;
        ELSIF x = 6871 THEN
            tanh_f := 2042;
        ELSIF x = 6872 THEN
            tanh_f := 2042;
        ELSIF x = 6873 THEN
            tanh_f := 2042;
        ELSIF x = 6874 THEN
            tanh_f := 2042;
        ELSIF x = 6875 THEN
            tanh_f := 2042;
        ELSIF x = 6876 THEN
            tanh_f := 2042;
        ELSIF x = 6877 THEN
            tanh_f := 2042;
        ELSIF x = 6878 THEN
            tanh_f := 2042;
        ELSIF x = 6879 THEN
            tanh_f := 2042;
        ELSIF x = 6880 THEN
            tanh_f := 2042;
        ELSIF x = 6881 THEN
            tanh_f := 2042;
        ELSIF x = 6882 THEN
            tanh_f := 2042;
        ELSIF x = 6883 THEN
            tanh_f := 2042;
        ELSIF x = 6884 THEN
            tanh_f := 2042;
        ELSIF x = 6885 THEN
            tanh_f := 2042;
        ELSIF x = 6886 THEN
            tanh_f := 2042;
        ELSIF x = 6887 THEN
            tanh_f := 2042;
        ELSIF x = 6888 THEN
            tanh_f := 2042;
        ELSIF x = 6889 THEN
            tanh_f := 2042;
        ELSIF x = 6890 THEN
            tanh_f := 2042;
        ELSIF x = 6891 THEN
            tanh_f := 2042;
        ELSIF x = 6892 THEN
            tanh_f := 2042;
        ELSIF x = 6893 THEN
            tanh_f := 2042;
        ELSIF x = 6894 THEN
            tanh_f := 2042;
        ELSIF x = 6895 THEN
            tanh_f := 2042;
        ELSIF x = 6896 THEN
            tanh_f := 2042;
        ELSIF x = 6897 THEN
            tanh_f := 2042;
        ELSIF x = 6898 THEN
            tanh_f := 2042;
        ELSIF x = 6899 THEN
            tanh_f := 2042;
        ELSIF x = 6900 THEN
            tanh_f := 2042;
        ELSIF x = 6901 THEN
            tanh_f := 2042;
        ELSIF x = 6902 THEN
            tanh_f := 2042;
        ELSIF x = 6903 THEN
            tanh_f := 2042;
        ELSIF x = 6904 THEN
            tanh_f := 2042;
        ELSIF x = 6905 THEN
            tanh_f := 2042;
        ELSIF x = 6906 THEN
            tanh_f := 2042;
        ELSIF x = 6907 THEN
            tanh_f := 2042;
        ELSIF x = 6908 THEN
            tanh_f := 2042;
        ELSIF x = 6909 THEN
            tanh_f := 2042;
        ELSIF x = 6910 THEN
            tanh_f := 2042;
        ELSIF x = 6911 THEN
            tanh_f := 2042;
        ELSIF x = 6912 THEN
            tanh_f := 2044;
        ELSIF x = 6913 THEN
            tanh_f := 2044;
        ELSIF x = 6914 THEN
            tanh_f := 2044;
        ELSIF x = 6915 THEN
            tanh_f := 2044;
        ELSIF x = 6916 THEN
            tanh_f := 2044;
        ELSIF x = 6917 THEN
            tanh_f := 2044;
        ELSIF x = 6918 THEN
            tanh_f := 2044;
        ELSIF x = 6919 THEN
            tanh_f := 2044;
        ELSIF x = 6920 THEN
            tanh_f := 2044;
        ELSIF x = 6921 THEN
            tanh_f := 2044;
        ELSIF x = 6922 THEN
            tanh_f := 2044;
        ELSIF x = 6923 THEN
            tanh_f := 2044;
        ELSIF x = 6924 THEN
            tanh_f := 2044;
        ELSIF x = 6925 THEN
            tanh_f := 2044;
        ELSIF x = 6926 THEN
            tanh_f := 2044;
        ELSIF x = 6927 THEN
            tanh_f := 2044;
        ELSIF x = 6928 THEN
            tanh_f := 2044;
        ELSIF x = 6929 THEN
            tanh_f := 2044;
        ELSIF x = 6930 THEN
            tanh_f := 2044;
        ELSIF x = 6931 THEN
            tanh_f := 2044;
        ELSIF x = 6932 THEN
            tanh_f := 2044;
        ELSIF x = 6933 THEN
            tanh_f := 2044;
        ELSIF x = 6934 THEN
            tanh_f := 2044;
        ELSIF x = 6935 THEN
            tanh_f := 2044;
        ELSIF x = 6936 THEN
            tanh_f := 2044;
        ELSIF x = 6937 THEN
            tanh_f := 2044;
        ELSIF x = 6938 THEN
            tanh_f := 2044;
        ELSIF x = 6939 THEN
            tanh_f := 2044;
        ELSIF x = 6940 THEN
            tanh_f := 2044;
        ELSIF x = 6941 THEN
            tanh_f := 2044;
        ELSIF x = 6942 THEN
            tanh_f := 2044;
        ELSIF x = 6943 THEN
            tanh_f := 2044;
        ELSIF x = 6944 THEN
            tanh_f := 2044;
        ELSIF x = 6945 THEN
            tanh_f := 2044;
        ELSIF x = 6946 THEN
            tanh_f := 2044;
        ELSIF x = 6947 THEN
            tanh_f := 2044;
        ELSIF x = 6948 THEN
            tanh_f := 2044;
        ELSIF x = 6949 THEN
            tanh_f := 2044;
        ELSIF x = 6950 THEN
            tanh_f := 2044;
        ELSIF x = 6951 THEN
            tanh_f := 2044;
        ELSIF x = 6952 THEN
            tanh_f := 2044;
        ELSIF x = 6953 THEN
            tanh_f := 2044;
        ELSIF x = 6954 THEN
            tanh_f := 2044;
        ELSIF x = 6955 THEN
            tanh_f := 2044;
        ELSIF x = 6956 THEN
            tanh_f := 2044;
        ELSIF x = 6957 THEN
            tanh_f := 2044;
        ELSIF x = 6958 THEN
            tanh_f := 2044;
        ELSIF x = 6959 THEN
            tanh_f := 2044;
        ELSIF x = 6960 THEN
            tanh_f := 2044;
        ELSIF x = 6961 THEN
            tanh_f := 2044;
        ELSIF x = 6962 THEN
            tanh_f := 2044;
        ELSIF x = 6963 THEN
            tanh_f := 2044;
        ELSIF x = 6964 THEN
            tanh_f := 2044;
        ELSIF x = 6965 THEN
            tanh_f := 2044;
        ELSIF x = 6966 THEN
            tanh_f := 2044;
        ELSIF x = 6967 THEN
            tanh_f := 2044;
        ELSIF x = 6968 THEN
            tanh_f := 2044;
        ELSIF x = 6969 THEN
            tanh_f := 2044;
        ELSIF x = 6970 THEN
            tanh_f := 2044;
        ELSIF x = 6971 THEN
            tanh_f := 2044;
        ELSIF x = 6972 THEN
            tanh_f := 2044;
        ELSIF x = 6973 THEN
            tanh_f := 2044;
        ELSIF x = 6974 THEN
            tanh_f := 2044;
        ELSIF x = 6975 THEN
            tanh_f := 2044;
        ELSIF x = 6976 THEN
            tanh_f := 2044;
        ELSIF x = 6977 THEN
            tanh_f := 2044;
        ELSIF x = 6978 THEN
            tanh_f := 2044;
        ELSIF x = 6979 THEN
            tanh_f := 2044;
        ELSIF x = 6980 THEN
            tanh_f := 2044;
        ELSIF x = 6981 THEN
            tanh_f := 2044;
        ELSIF x = 6982 THEN
            tanh_f := 2044;
        ELSIF x = 6983 THEN
            tanh_f := 2044;
        ELSIF x = 6984 THEN
            tanh_f := 2044;
        ELSIF x = 6985 THEN
            tanh_f := 2044;
        ELSIF x = 6986 THEN
            tanh_f := 2044;
        ELSIF x = 6987 THEN
            tanh_f := 2044;
        ELSIF x = 6988 THEN
            tanh_f := 2044;
        ELSIF x = 6989 THEN
            tanh_f := 2044;
        ELSIF x = 6990 THEN
            tanh_f := 2044;
        ELSIF x = 6991 THEN
            tanh_f := 2044;
        ELSIF x = 6992 THEN
            tanh_f := 2044;
        ELSIF x = 6993 THEN
            tanh_f := 2044;
        ELSIF x = 6994 THEN
            tanh_f := 2044;
        ELSIF x = 6995 THEN
            tanh_f := 2044;
        ELSIF x = 6996 THEN
            tanh_f := 2044;
        ELSIF x = 6997 THEN
            tanh_f := 2044;
        ELSIF x = 6998 THEN
            tanh_f := 2044;
        ELSIF x = 6999 THEN
            tanh_f := 2044;
        ELSIF x = 7000 THEN
            tanh_f := 2044;
        ELSIF x = 7001 THEN
            tanh_f := 2044;
        ELSIF x = 7002 THEN
            tanh_f := 2044;
        ELSIF x = 7003 THEN
            tanh_f := 2044;
        ELSIF x = 7004 THEN
            tanh_f := 2044;
        ELSIF x = 7005 THEN
            tanh_f := 2044;
        ELSIF x = 7006 THEN
            tanh_f := 2044;
        ELSIF x = 7007 THEN
            tanh_f := 2044;
        ELSIF x = 7008 THEN
            tanh_f := 2044;
        ELSIF x = 7009 THEN
            tanh_f := 2044;
        ELSIF x = 7010 THEN
            tanh_f := 2044;
        ELSIF x = 7011 THEN
            tanh_f := 2044;
        ELSIF x = 7012 THEN
            tanh_f := 2044;
        ELSIF x = 7013 THEN
            tanh_f := 2044;
        ELSIF x = 7014 THEN
            tanh_f := 2044;
        ELSIF x = 7015 THEN
            tanh_f := 2044;
        ELSIF x = 7016 THEN
            tanh_f := 2044;
        ELSIF x = 7017 THEN
            tanh_f := 2044;
        ELSIF x = 7018 THEN
            tanh_f := 2044;
        ELSIF x = 7019 THEN
            tanh_f := 2044;
        ELSIF x = 7020 THEN
            tanh_f := 2044;
        ELSIF x = 7021 THEN
            tanh_f := 2044;
        ELSIF x = 7022 THEN
            tanh_f := 2044;
        ELSIF x = 7023 THEN
            tanh_f := 2044;
        ELSIF x = 7024 THEN
            tanh_f := 2044;
        ELSIF x = 7025 THEN
            tanh_f := 2044;
        ELSIF x = 7026 THEN
            tanh_f := 2044;
        ELSIF x = 7027 THEN
            tanh_f := 2044;
        ELSIF x = 7028 THEN
            tanh_f := 2044;
        ELSIF x = 7029 THEN
            tanh_f := 2044;
        ELSIF x = 7030 THEN
            tanh_f := 2044;
        ELSIF x = 7031 THEN
            tanh_f := 2044;
        ELSIF x = 7032 THEN
            tanh_f := 2044;
        ELSIF x = 7033 THEN
            tanh_f := 2044;
        ELSIF x = 7034 THEN
            tanh_f := 2044;
        ELSIF x = 7035 THEN
            tanh_f := 2044;
        ELSIF x = 7036 THEN
            tanh_f := 2044;
        ELSIF x = 7037 THEN
            tanh_f := 2044;
        ELSIF x = 7038 THEN
            tanh_f := 2044;
        ELSIF x = 7039 THEN
            tanh_f := 2044;
        ELSIF x = 7040 THEN
            tanh_f := 2044;
        ELSIF x = 7041 THEN
            tanh_f := 2044;
        ELSIF x = 7042 THEN
            tanh_f := 2044;
        ELSIF x = 7043 THEN
            tanh_f := 2044;
        ELSIF x = 7044 THEN
            tanh_f := 2044;
        ELSIF x = 7045 THEN
            tanh_f := 2044;
        ELSIF x = 7046 THEN
            tanh_f := 2044;
        ELSIF x = 7047 THEN
            tanh_f := 2044;
        ELSIF x = 7048 THEN
            tanh_f := 2044;
        ELSIF x = 7049 THEN
            tanh_f := 2044;
        ELSIF x = 7050 THEN
            tanh_f := 2044;
        ELSIF x = 7051 THEN
            tanh_f := 2044;
        ELSIF x = 7052 THEN
            tanh_f := 2044;
        ELSIF x = 7053 THEN
            tanh_f := 2044;
        ELSIF x = 7054 THEN
            tanh_f := 2044;
        ELSIF x = 7055 THEN
            tanh_f := 2044;
        ELSIF x = 7056 THEN
            tanh_f := 2044;
        ELSIF x = 7057 THEN
            tanh_f := 2044;
        ELSIF x = 7058 THEN
            tanh_f := 2044;
        ELSIF x = 7059 THEN
            tanh_f := 2044;
        ELSIF x = 7060 THEN
            tanh_f := 2044;
        ELSIF x = 7061 THEN
            tanh_f := 2044;
        ELSIF x = 7062 THEN
            tanh_f := 2044;
        ELSIF x = 7063 THEN
            tanh_f := 2044;
        ELSIF x = 7064 THEN
            tanh_f := 2044;
        ELSIF x = 7065 THEN
            tanh_f := 2044;
        ELSIF x = 7066 THEN
            tanh_f := 2044;
        ELSIF x = 7067 THEN
            tanh_f := 2044;
        ELSIF x = 7068 THEN
            tanh_f := 2044;
        ELSIF x = 7069 THEN
            tanh_f := 2044;
        ELSIF x = 7070 THEN
            tanh_f := 2044;
        ELSIF x = 7071 THEN
            tanh_f := 2044;
        ELSIF x = 7072 THEN
            tanh_f := 2044;
        ELSIF x = 7073 THEN
            tanh_f := 2044;
        ELSIF x = 7074 THEN
            tanh_f := 2044;
        ELSIF x = 7075 THEN
            tanh_f := 2044;
        ELSIF x = 7076 THEN
            tanh_f := 2044;
        ELSIF x = 7077 THEN
            tanh_f := 2044;
        ELSIF x = 7078 THEN
            tanh_f := 2044;
        ELSIF x = 7079 THEN
            tanh_f := 2044;
        ELSIF x = 7080 THEN
            tanh_f := 2044;
        ELSIF x = 7081 THEN
            tanh_f := 2044;
        ELSIF x = 7082 THEN
            tanh_f := 2044;
        ELSIF x = 7083 THEN
            tanh_f := 2044;
        ELSIF x = 7084 THEN
            tanh_f := 2044;
        ELSIF x = 7085 THEN
            tanh_f := 2044;
        ELSIF x = 7086 THEN
            tanh_f := 2044;
        ELSIF x = 7087 THEN
            tanh_f := 2044;
        ELSIF x = 7088 THEN
            tanh_f := 2044;
        ELSIF x = 7089 THEN
            tanh_f := 2044;
        ELSIF x = 7090 THEN
            tanh_f := 2044;
        ELSIF x = 7091 THEN
            tanh_f := 2044;
        ELSIF x = 7092 THEN
            tanh_f := 2044;
        ELSIF x = 7093 THEN
            tanh_f := 2044;
        ELSIF x = 7094 THEN
            tanh_f := 2044;
        ELSIF x = 7095 THEN
            tanh_f := 2044;
        ELSIF x = 7096 THEN
            tanh_f := 2044;
        ELSIF x = 7097 THEN
            tanh_f := 2044;
        ELSIF x = 7098 THEN
            tanh_f := 2044;
        ELSIF x = 7099 THEN
            tanh_f := 2044;
        ELSIF x = 7100 THEN
            tanh_f := 2044;
        ELSIF x = 7101 THEN
            tanh_f := 2044;
        ELSIF x = 7102 THEN
            tanh_f := 2044;
        ELSIF x = 7103 THEN
            tanh_f := 2044;
        ELSIF x = 7104 THEN
            tanh_f := 2044;
        ELSIF x = 7105 THEN
            tanh_f := 2044;
        ELSIF x = 7106 THEN
            tanh_f := 2044;
        ELSIF x = 7107 THEN
            tanh_f := 2044;
        ELSIF x = 7108 THEN
            tanh_f := 2044;
        ELSIF x = 7109 THEN
            tanh_f := 2044;
        ELSIF x = 7110 THEN
            tanh_f := 2044;
        ELSIF x = 7111 THEN
            tanh_f := 2044;
        ELSIF x = 7112 THEN
            tanh_f := 2044;
        ELSIF x = 7113 THEN
            tanh_f := 2044;
        ELSIF x = 7114 THEN
            tanh_f := 2044;
        ELSIF x = 7115 THEN
            tanh_f := 2044;
        ELSIF x = 7116 THEN
            tanh_f := 2044;
        ELSIF x = 7117 THEN
            tanh_f := 2044;
        ELSIF x = 7118 THEN
            tanh_f := 2044;
        ELSIF x = 7119 THEN
            tanh_f := 2044;
        ELSIF x = 7120 THEN
            tanh_f := 2044;
        ELSIF x = 7121 THEN
            tanh_f := 2044;
        ELSIF x = 7122 THEN
            tanh_f := 2044;
        ELSIF x = 7123 THEN
            tanh_f := 2044;
        ELSIF x = 7124 THEN
            tanh_f := 2044;
        ELSIF x = 7125 THEN
            tanh_f := 2044;
        ELSIF x = 7126 THEN
            tanh_f := 2044;
        ELSIF x = 7127 THEN
            tanh_f := 2044;
        ELSIF x = 7128 THEN
            tanh_f := 2044;
        ELSIF x = 7129 THEN
            tanh_f := 2044;
        ELSIF x = 7130 THEN
            tanh_f := 2044;
        ELSIF x = 7131 THEN
            tanh_f := 2044;
        ELSIF x = 7132 THEN
            tanh_f := 2044;
        ELSIF x = 7133 THEN
            tanh_f := 2044;
        ELSIF x = 7134 THEN
            tanh_f := 2044;
        ELSIF x = 7135 THEN
            tanh_f := 2044;
        ELSIF x = 7136 THEN
            tanh_f := 2044;
        ELSIF x = 7137 THEN
            tanh_f := 2044;
        ELSIF x = 7138 THEN
            tanh_f := 2044;
        ELSIF x = 7139 THEN
            tanh_f := 2044;
        ELSIF x = 7140 THEN
            tanh_f := 2044;
        ELSIF x = 7141 THEN
            tanh_f := 2044;
        ELSIF x = 7142 THEN
            tanh_f := 2044;
        ELSIF x = 7143 THEN
            tanh_f := 2044;
        ELSIF x = 7144 THEN
            tanh_f := 2044;
        ELSIF x = 7145 THEN
            tanh_f := 2044;
        ELSIF x = 7146 THEN
            tanh_f := 2044;
        ELSIF x = 7147 THEN
            tanh_f := 2044;
        ELSIF x = 7148 THEN
            tanh_f := 2044;
        ELSIF x = 7149 THEN
            tanh_f := 2044;
        ELSIF x = 7150 THEN
            tanh_f := 2044;
        ELSIF x = 7151 THEN
            tanh_f := 2044;
        ELSIF x = 7152 THEN
            tanh_f := 2044;
        ELSIF x = 7153 THEN
            tanh_f := 2044;
        ELSIF x = 7154 THEN
            tanh_f := 2044;
        ELSIF x = 7155 THEN
            tanh_f := 2044;
        ELSIF x = 7156 THEN
            tanh_f := 2044;
        ELSIF x = 7157 THEN
            tanh_f := 2044;
        ELSIF x = 7158 THEN
            tanh_f := 2044;
        ELSIF x = 7159 THEN
            tanh_f := 2044;
        ELSIF x = 7160 THEN
            tanh_f := 2044;
        ELSIF x = 7161 THEN
            tanh_f := 2044;
        ELSIF x = 7162 THEN
            tanh_f := 2044;
        ELSIF x = 7163 THEN
            tanh_f := 2044;
        ELSIF x = 7164 THEN
            tanh_f := 2044;
        ELSIF x = 7165 THEN
            tanh_f := 2044;
        ELSIF x = 7166 THEN
            tanh_f := 2044;
        ELSIF x = 7167 THEN
            tanh_f := 2044;
        ELSIF x = 7168 THEN
            tanh_f := 2044;
        ELSIF x = 7169 THEN
            tanh_f := 2044;
        ELSIF x = 7170 THEN
            tanh_f := 2044;
        ELSIF x = 7171 THEN
            tanh_f := 2044;
        ELSIF x = 7172 THEN
            tanh_f := 2044;
        ELSIF x = 7173 THEN
            tanh_f := 2044;
        ELSIF x = 7174 THEN
            tanh_f := 2044;
        ELSIF x = 7175 THEN
            tanh_f := 2044;
        ELSIF x = 7176 THEN
            tanh_f := 2044;
        ELSIF x = 7177 THEN
            tanh_f := 2044;
        ELSIF x = 7178 THEN
            tanh_f := 2044;
        ELSIF x = 7179 THEN
            tanh_f := 2044;
        ELSIF x = 7180 THEN
            tanh_f := 2044;
        ELSIF x = 7181 THEN
            tanh_f := 2044;
        ELSIF x = 7182 THEN
            tanh_f := 2044;
        ELSIF x = 7183 THEN
            tanh_f := 2044;
        ELSIF x = 7184 THEN
            tanh_f := 2044;
        ELSIF x = 7185 THEN
            tanh_f := 2044;
        ELSIF x = 7186 THEN
            tanh_f := 2044;
        ELSIF x = 7187 THEN
            tanh_f := 2044;
        ELSIF x = 7188 THEN
            tanh_f := 2044;
        ELSIF x = 7189 THEN
            tanh_f := 2044;
        ELSIF x = 7190 THEN
            tanh_f := 2044;
        ELSIF x = 7191 THEN
            tanh_f := 2044;
        ELSIF x = 7192 THEN
            tanh_f := 2044;
        ELSIF x = 7193 THEN
            tanh_f := 2044;
        ELSIF x = 7194 THEN
            tanh_f := 2044;
        ELSIF x = 7195 THEN
            tanh_f := 2044;
        ELSIF x = 7196 THEN
            tanh_f := 2044;
        ELSIF x = 7197 THEN
            tanh_f := 2044;
        ELSIF x = 7198 THEN
            tanh_f := 2044;
        ELSIF x = 7199 THEN
            tanh_f := 2044;
        ELSIF x = 7200 THEN
            tanh_f := 2044;
        ELSIF x = 7201 THEN
            tanh_f := 2044;
        ELSIF x = 7202 THEN
            tanh_f := 2044;
        ELSIF x = 7203 THEN
            tanh_f := 2044;
        ELSIF x = 7204 THEN
            tanh_f := 2044;
        ELSIF x = 7205 THEN
            tanh_f := 2044;
        ELSIF x = 7206 THEN
            tanh_f := 2044;
        ELSIF x = 7207 THEN
            tanh_f := 2044;
        ELSIF x = 7208 THEN
            tanh_f := 2044;
        ELSIF x = 7209 THEN
            tanh_f := 2044;
        ELSIF x = 7210 THEN
            tanh_f := 2044;
        ELSIF x = 7211 THEN
            tanh_f := 2044;
        ELSIF x = 7212 THEN
            tanh_f := 2044;
        ELSIF x = 7213 THEN
            tanh_f := 2044;
        ELSIF x = 7214 THEN
            tanh_f := 2044;
        ELSIF x = 7215 THEN
            tanh_f := 2044;
        ELSIF x = 7216 THEN
            tanh_f := 2044;
        ELSIF x = 7217 THEN
            tanh_f := 2044;
        ELSIF x = 7218 THEN
            tanh_f := 2044;
        ELSIF x = 7219 THEN
            tanh_f := 2044;
        ELSIF x = 7220 THEN
            tanh_f := 2044;
        ELSIF x = 7221 THEN
            tanh_f := 2044;
        ELSIF x = 7222 THEN
            tanh_f := 2044;
        ELSIF x = 7223 THEN
            tanh_f := 2044;
        ELSIF x = 7224 THEN
            tanh_f := 2044;
        ELSIF x = 7225 THEN
            tanh_f := 2044;
        ELSIF x = 7226 THEN
            tanh_f := 2044;
        ELSIF x = 7227 THEN
            tanh_f := 2044;
        ELSIF x = 7228 THEN
            tanh_f := 2044;
        ELSIF x = 7229 THEN
            tanh_f := 2044;
        ELSIF x = 7230 THEN
            tanh_f := 2044;
        ELSIF x = 7231 THEN
            tanh_f := 2044;
        ELSIF x = 7232 THEN
            tanh_f := 2044;
        ELSIF x = 7233 THEN
            tanh_f := 2044;
        ELSIF x = 7234 THEN
            tanh_f := 2044;
        ELSIF x = 7235 THEN
            tanh_f := 2044;
        ELSIF x = 7236 THEN
            tanh_f := 2044;
        ELSIF x = 7237 THEN
            tanh_f := 2044;
        ELSIF x = 7238 THEN
            tanh_f := 2044;
        ELSIF x = 7239 THEN
            tanh_f := 2044;
        ELSIF x = 7240 THEN
            tanh_f := 2044;
        ELSIF x = 7241 THEN
            tanh_f := 2044;
        ELSIF x = 7242 THEN
            tanh_f := 2044;
        ELSIF x = 7243 THEN
            tanh_f := 2044;
        ELSIF x = 7244 THEN
            tanh_f := 2044;
        ELSIF x = 7245 THEN
            tanh_f := 2044;
        ELSIF x = 7246 THEN
            tanh_f := 2044;
        ELSIF x = 7247 THEN
            tanh_f := 2044;
        ELSIF x = 7248 THEN
            tanh_f := 2044;
        ELSIF x = 7249 THEN
            tanh_f := 2044;
        ELSIF x = 7250 THEN
            tanh_f := 2044;
        ELSIF x = 7251 THEN
            tanh_f := 2044;
        ELSIF x = 7252 THEN
            tanh_f := 2044;
        ELSIF x = 7253 THEN
            tanh_f := 2044;
        ELSIF x = 7254 THEN
            tanh_f := 2044;
        ELSIF x = 7255 THEN
            tanh_f := 2044;
        ELSIF x = 7256 THEN
            tanh_f := 2044;
        ELSIF x = 7257 THEN
            tanh_f := 2044;
        ELSIF x = 7258 THEN
            tanh_f := 2044;
        ELSIF x = 7259 THEN
            tanh_f := 2044;
        ELSIF x = 7260 THEN
            tanh_f := 2044;
        ELSIF x = 7261 THEN
            tanh_f := 2044;
        ELSIF x = 7262 THEN
            tanh_f := 2044;
        ELSIF x = 7263 THEN
            tanh_f := 2044;
        ELSIF x = 7264 THEN
            tanh_f := 2044;
        ELSIF x = 7265 THEN
            tanh_f := 2044;
        ELSIF x = 7266 THEN
            tanh_f := 2044;
        ELSIF x = 7267 THEN
            tanh_f := 2044;
        ELSIF x = 7268 THEN
            tanh_f := 2044;
        ELSIF x = 7269 THEN
            tanh_f := 2044;
        ELSIF x = 7270 THEN
            tanh_f := 2044;
        ELSIF x = 7271 THEN
            tanh_f := 2044;
        ELSIF x = 7272 THEN
            tanh_f := 2044;
        ELSIF x = 7273 THEN
            tanh_f := 2044;
        ELSIF x = 7274 THEN
            tanh_f := 2044;
        ELSIF x = 7275 THEN
            tanh_f := 2044;
        ELSIF x = 7276 THEN
            tanh_f := 2044;
        ELSIF x = 7277 THEN
            tanh_f := 2044;
        ELSIF x = 7278 THEN
            tanh_f := 2044;
        ELSIF x = 7279 THEN
            tanh_f := 2044;
        ELSIF x = 7280 THEN
            tanh_f := 2044;
        ELSIF x = 7281 THEN
            tanh_f := 2044;
        ELSIF x = 7282 THEN
            tanh_f := 2044;
        ELSIF x = 7283 THEN
            tanh_f := 2044;
        ELSIF x = 7284 THEN
            tanh_f := 2044;
        ELSIF x = 7285 THEN
            tanh_f := 2044;
        ELSIF x = 7286 THEN
            tanh_f := 2044;
        ELSIF x = 7287 THEN
            tanh_f := 2044;
        ELSIF x = 7288 THEN
            tanh_f := 2044;
        ELSIF x = 7289 THEN
            tanh_f := 2044;
        ELSIF x = 7290 THEN
            tanh_f := 2044;
        ELSIF x = 7291 THEN
            tanh_f := 2044;
        ELSIF x = 7292 THEN
            tanh_f := 2044;
        ELSIF x = 7293 THEN
            tanh_f := 2044;
        ELSIF x = 7294 THEN
            tanh_f := 2044;
        ELSIF x = 7295 THEN
            tanh_f := 2044;
        ELSIF x = 7296 THEN
            tanh_f := 2044;
        ELSIF x = 7297 THEN
            tanh_f := 2044;
        ELSIF x = 7298 THEN
            tanh_f := 2044;
        ELSIF x = 7299 THEN
            tanh_f := 2044;
        ELSIF x = 7300 THEN
            tanh_f := 2044;
        ELSIF x = 7301 THEN
            tanh_f := 2044;
        ELSIF x = 7302 THEN
            tanh_f := 2044;
        ELSIF x = 7303 THEN
            tanh_f := 2044;
        ELSIF x = 7304 THEN
            tanh_f := 2044;
        ELSIF x = 7305 THEN
            tanh_f := 2044;
        ELSIF x = 7306 THEN
            tanh_f := 2044;
        ELSIF x = 7307 THEN
            tanh_f := 2044;
        ELSIF x = 7308 THEN
            tanh_f := 2044;
        ELSIF x = 7309 THEN
            tanh_f := 2044;
        ELSIF x = 7310 THEN
            tanh_f := 2044;
        ELSIF x = 7311 THEN
            tanh_f := 2044;
        ELSIF x = 7312 THEN
            tanh_f := 2044;
        ELSIF x = 7313 THEN
            tanh_f := 2044;
        ELSIF x = 7314 THEN
            tanh_f := 2044;
        ELSIF x = 7315 THEN
            tanh_f := 2044;
        ELSIF x = 7316 THEN
            tanh_f := 2044;
        ELSIF x = 7317 THEN
            tanh_f := 2044;
        ELSIF x = 7318 THEN
            tanh_f := 2044;
        ELSIF x = 7319 THEN
            tanh_f := 2044;
        ELSIF x = 7320 THEN
            tanh_f := 2044;
        ELSIF x = 7321 THEN
            tanh_f := 2044;
        ELSIF x = 7322 THEN
            tanh_f := 2044;
        ELSIF x = 7323 THEN
            tanh_f := 2044;
        ELSIF x = 7324 THEN
            tanh_f := 2044;
        ELSIF x = 7325 THEN
            tanh_f := 2044;
        ELSIF x = 7326 THEN
            tanh_f := 2044;
        ELSIF x = 7327 THEN
            tanh_f := 2044;
        ELSIF x = 7328 THEN
            tanh_f := 2044;
        ELSIF x = 7329 THEN
            tanh_f := 2044;
        ELSIF x = 7330 THEN
            tanh_f := 2044;
        ELSIF x = 7331 THEN
            tanh_f := 2044;
        ELSIF x = 7332 THEN
            tanh_f := 2044;
        ELSIF x = 7333 THEN
            tanh_f := 2044;
        ELSIF x = 7334 THEN
            tanh_f := 2044;
        ELSIF x = 7335 THEN
            tanh_f := 2044;
        ELSIF x = 7336 THEN
            tanh_f := 2044;
        ELSIF x = 7337 THEN
            tanh_f := 2044;
        ELSIF x = 7338 THEN
            tanh_f := 2044;
        ELSIF x = 7339 THEN
            tanh_f := 2044;
        ELSIF x = 7340 THEN
            tanh_f := 2044;
        ELSIF x = 7341 THEN
            tanh_f := 2044;
        ELSIF x = 7342 THEN
            tanh_f := 2044;
        ELSIF x = 7343 THEN
            tanh_f := 2044;
        ELSIF x = 7344 THEN
            tanh_f := 2044;
        ELSIF x = 7345 THEN
            tanh_f := 2044;
        ELSIF x = 7346 THEN
            tanh_f := 2044;
        ELSIF x = 7347 THEN
            tanh_f := 2044;
        ELSIF x = 7348 THEN
            tanh_f := 2044;
        ELSIF x = 7349 THEN
            tanh_f := 2044;
        ELSIF x = 7350 THEN
            tanh_f := 2044;
        ELSIF x = 7351 THEN
            tanh_f := 2044;
        ELSIF x = 7352 THEN
            tanh_f := 2044;
        ELSIF x = 7353 THEN
            tanh_f := 2044;
        ELSIF x = 7354 THEN
            tanh_f := 2044;
        ELSIF x = 7355 THEN
            tanh_f := 2044;
        ELSIF x = 7356 THEN
            tanh_f := 2044;
        ELSIF x = 7357 THEN
            tanh_f := 2044;
        ELSIF x = 7358 THEN
            tanh_f := 2044;
        ELSIF x = 7359 THEN
            tanh_f := 2044;
        ELSIF x = 7360 THEN
            tanh_f := 2044;
        ELSIF x = 7361 THEN
            tanh_f := 2044;
        ELSIF x = 7362 THEN
            tanh_f := 2044;
        ELSIF x = 7363 THEN
            tanh_f := 2044;
        ELSIF x = 7364 THEN
            tanh_f := 2044;
        ELSIF x = 7365 THEN
            tanh_f := 2044;
        ELSIF x = 7366 THEN
            tanh_f := 2044;
        ELSIF x = 7367 THEN
            tanh_f := 2044;
        ELSIF x = 7368 THEN
            tanh_f := 2044;
        ELSIF x = 7369 THEN
            tanh_f := 2044;
        ELSIF x = 7370 THEN
            tanh_f := 2044;
        ELSIF x = 7371 THEN
            tanh_f := 2044;
        ELSIF x = 7372 THEN
            tanh_f := 2044;
        ELSIF x = 7373 THEN
            tanh_f := 2044;
        ELSIF x = 7374 THEN
            tanh_f := 2044;
        ELSIF x = 7375 THEN
            tanh_f := 2044;
        ELSIF x = 7376 THEN
            tanh_f := 2044;
        ELSIF x = 7377 THEN
            tanh_f := 2044;
        ELSIF x = 7378 THEN
            tanh_f := 2044;
        ELSIF x = 7379 THEN
            tanh_f := 2044;
        ELSIF x = 7380 THEN
            tanh_f := 2044;
        ELSIF x = 7381 THEN
            tanh_f := 2044;
        ELSIF x = 7382 THEN
            tanh_f := 2044;
        ELSIF x = 7383 THEN
            tanh_f := 2044;
        ELSIF x = 7384 THEN
            tanh_f := 2044;
        ELSIF x = 7385 THEN
            tanh_f := 2044;
        ELSIF x = 7386 THEN
            tanh_f := 2044;
        ELSIF x = 7387 THEN
            tanh_f := 2044;
        ELSIF x = 7388 THEN
            tanh_f := 2044;
        ELSIF x = 7389 THEN
            tanh_f := 2044;
        ELSIF x = 7390 THEN
            tanh_f := 2044;
        ELSIF x = 7391 THEN
            tanh_f := 2044;
        ELSIF x = 7392 THEN
            tanh_f := 2044;
        ELSIF x = 7393 THEN
            tanh_f := 2044;
        ELSIF x = 7394 THEN
            tanh_f := 2044;
        ELSIF x = 7395 THEN
            tanh_f := 2044;
        ELSIF x = 7396 THEN
            tanh_f := 2044;
        ELSIF x = 7397 THEN
            tanh_f := 2044;
        ELSIF x = 7398 THEN
            tanh_f := 2044;
        ELSIF x = 7399 THEN
            tanh_f := 2044;
        ELSIF x = 7400 THEN
            tanh_f := 2044;
        ELSIF x = 7401 THEN
            tanh_f := 2044;
        ELSIF x = 7402 THEN
            tanh_f := 2044;
        ELSIF x = 7403 THEN
            tanh_f := 2044;
        ELSIF x = 7404 THEN
            tanh_f := 2044;
        ELSIF x = 7405 THEN
            tanh_f := 2044;
        ELSIF x = 7406 THEN
            tanh_f := 2044;
        ELSIF x = 7407 THEN
            tanh_f := 2044;
        ELSIF x = 7408 THEN
            tanh_f := 2044;
        ELSIF x = 7409 THEN
            tanh_f := 2044;
        ELSIF x = 7410 THEN
            tanh_f := 2044;
        ELSIF x = 7411 THEN
            tanh_f := 2044;
        ELSIF x = 7412 THEN
            tanh_f := 2044;
        ELSIF x = 7413 THEN
            tanh_f := 2044;
        ELSIF x = 7414 THEN
            tanh_f := 2044;
        ELSIF x = 7415 THEN
            tanh_f := 2044;
        ELSIF x = 7416 THEN
            tanh_f := 2044;
        ELSIF x = 7417 THEN
            tanh_f := 2044;
        ELSIF x = 7418 THEN
            tanh_f := 2044;
        ELSIF x = 7419 THEN
            tanh_f := 2044;
        ELSIF x = 7420 THEN
            tanh_f := 2044;
        ELSIF x = 7421 THEN
            tanh_f := 2044;
        ELSIF x = 7422 THEN
            tanh_f := 2044;
        ELSIF x = 7423 THEN
            tanh_f := 2044;
        ELSIF x = 7424 THEN
            tanh_f := 2046;
        ELSIF x = 7425 THEN
            tanh_f := 2046;
        ELSIF x = 7426 THEN
            tanh_f := 2046;
        ELSIF x = 7427 THEN
            tanh_f := 2046;
        ELSIF x = 7428 THEN
            tanh_f := 2046;
        ELSIF x = 7429 THEN
            tanh_f := 2046;
        ELSIF x = 7430 THEN
            tanh_f := 2046;
        ELSIF x = 7431 THEN
            tanh_f := 2046;
        ELSIF x = 7432 THEN
            tanh_f := 2046;
        ELSIF x = 7433 THEN
            tanh_f := 2046;
        ELSIF x = 7434 THEN
            tanh_f := 2046;
        ELSIF x = 7435 THEN
            tanh_f := 2046;
        ELSIF x = 7436 THEN
            tanh_f := 2046;
        ELSIF x = 7437 THEN
            tanh_f := 2046;
        ELSIF x = 7438 THEN
            tanh_f := 2046;
        ELSIF x = 7439 THEN
            tanh_f := 2046;
        ELSIF x = 7440 THEN
            tanh_f := 2046;
        ELSIF x = 7441 THEN
            tanh_f := 2046;
        ELSIF x = 7442 THEN
            tanh_f := 2046;
        ELSIF x = 7443 THEN
            tanh_f := 2046;
        ELSIF x = 7444 THEN
            tanh_f := 2046;
        ELSIF x = 7445 THEN
            tanh_f := 2046;
        ELSIF x = 7446 THEN
            tanh_f := 2046;
        ELSIF x = 7447 THEN
            tanh_f := 2046;
        ELSIF x = 7448 THEN
            tanh_f := 2046;
        ELSIF x = 7449 THEN
            tanh_f := 2046;
        ELSIF x = 7450 THEN
            tanh_f := 2046;
        ELSIF x = 7451 THEN
            tanh_f := 2046;
        ELSIF x = 7452 THEN
            tanh_f := 2046;
        ELSIF x = 7453 THEN
            tanh_f := 2046;
        ELSIF x = 7454 THEN
            tanh_f := 2046;
        ELSIF x = 7455 THEN
            tanh_f := 2046;
        ELSIF x = 7456 THEN
            tanh_f := 2046;
        ELSIF x = 7457 THEN
            tanh_f := 2046;
        ELSIF x = 7458 THEN
            tanh_f := 2046;
        ELSIF x = 7459 THEN
            tanh_f := 2046;
        ELSIF x = 7460 THEN
            tanh_f := 2046;
        ELSIF x = 7461 THEN
            tanh_f := 2046;
        ELSIF x = 7462 THEN
            tanh_f := 2046;
        ELSIF x = 7463 THEN
            tanh_f := 2046;
        ELSIF x = 7464 THEN
            tanh_f := 2046;
        ELSIF x = 7465 THEN
            tanh_f := 2046;
        ELSIF x = 7466 THEN
            tanh_f := 2046;
        ELSIF x = 7467 THEN
            tanh_f := 2046;
        ELSIF x = 7468 THEN
            tanh_f := 2046;
        ELSIF x = 7469 THEN
            tanh_f := 2046;
        ELSIF x = 7470 THEN
            tanh_f := 2046;
        ELSIF x = 7471 THEN
            tanh_f := 2046;
        ELSIF x = 7472 THEN
            tanh_f := 2046;
        ELSIF x = 7473 THEN
            tanh_f := 2046;
        ELSIF x = 7474 THEN
            tanh_f := 2046;
        ELSIF x = 7475 THEN
            tanh_f := 2046;
        ELSIF x = 7476 THEN
            tanh_f := 2046;
        ELSIF x = 7477 THEN
            tanh_f := 2046;
        ELSIF x = 7478 THEN
            tanh_f := 2046;
        ELSIF x = 7479 THEN
            tanh_f := 2046;
        ELSIF x = 7480 THEN
            tanh_f := 2046;
        ELSIF x = 7481 THEN
            tanh_f := 2046;
        ELSIF x = 7482 THEN
            tanh_f := 2046;
        ELSIF x = 7483 THEN
            tanh_f := 2046;
        ELSIF x = 7484 THEN
            tanh_f := 2046;
        ELSIF x = 7485 THEN
            tanh_f := 2046;
        ELSIF x = 7486 THEN
            tanh_f := 2046;
        ELSIF x = 7487 THEN
            tanh_f := 2046;
        ELSIF x = 7488 THEN
            tanh_f := 2046;
        ELSIF x = 7489 THEN
            tanh_f := 2046;
        ELSIF x = 7490 THEN
            tanh_f := 2046;
        ELSIF x = 7491 THEN
            tanh_f := 2046;
        ELSIF x = 7492 THEN
            tanh_f := 2046;
        ELSIF x = 7493 THEN
            tanh_f := 2046;
        ELSIF x = 7494 THEN
            tanh_f := 2046;
        ELSIF x = 7495 THEN
            tanh_f := 2046;
        ELSIF x = 7496 THEN
            tanh_f := 2046;
        ELSIF x = 7497 THEN
            tanh_f := 2046;
        ELSIF x = 7498 THEN
            tanh_f := 2046;
        ELSIF x = 7499 THEN
            tanh_f := 2046;
        ELSIF x = 7500 THEN
            tanh_f := 2046;
        ELSIF x = 7501 THEN
            tanh_f := 2046;
        ELSIF x = 7502 THEN
            tanh_f := 2046;
        ELSIF x = 7503 THEN
            tanh_f := 2046;
        ELSIF x = 7504 THEN
            tanh_f := 2046;
        ELSIF x = 7505 THEN
            tanh_f := 2046;
        ELSIF x = 7506 THEN
            tanh_f := 2046;
        ELSIF x = 7507 THEN
            tanh_f := 2046;
        ELSIF x = 7508 THEN
            tanh_f := 2046;
        ELSIF x = 7509 THEN
            tanh_f := 2046;
        ELSIF x = 7510 THEN
            tanh_f := 2046;
        ELSIF x = 7511 THEN
            tanh_f := 2046;
        ELSIF x = 7512 THEN
            tanh_f := 2046;
        ELSIF x = 7513 THEN
            tanh_f := 2046;
        ELSIF x = 7514 THEN
            tanh_f := 2046;
        ELSIF x = 7515 THEN
            tanh_f := 2046;
        ELSIF x = 7516 THEN
            tanh_f := 2046;
        ELSIF x = 7517 THEN
            tanh_f := 2046;
        ELSIF x = 7518 THEN
            tanh_f := 2046;
        ELSIF x = 7519 THEN
            tanh_f := 2046;
        ELSIF x = 7520 THEN
            tanh_f := 2046;
        ELSIF x = 7521 THEN
            tanh_f := 2046;
        ELSIF x = 7522 THEN
            tanh_f := 2046;
        ELSIF x = 7523 THEN
            tanh_f := 2046;
        ELSIF x = 7524 THEN
            tanh_f := 2046;
        ELSIF x = 7525 THEN
            tanh_f := 2046;
        ELSIF x = 7526 THEN
            tanh_f := 2046;
        ELSIF x = 7527 THEN
            tanh_f := 2046;
        ELSIF x = 7528 THEN
            tanh_f := 2046;
        ELSIF x = 7529 THEN
            tanh_f := 2046;
        ELSIF x = 7530 THEN
            tanh_f := 2046;
        ELSIF x = 7531 THEN
            tanh_f := 2046;
        ELSIF x = 7532 THEN
            tanh_f := 2046;
        ELSIF x = 7533 THEN
            tanh_f := 2046;
        ELSIF x = 7534 THEN
            tanh_f := 2046;
        ELSIF x = 7535 THEN
            tanh_f := 2046;
        ELSIF x = 7536 THEN
            tanh_f := 2046;
        ELSIF x = 7537 THEN
            tanh_f := 2046;
        ELSIF x = 7538 THEN
            tanh_f := 2046;
        ELSIF x = 7539 THEN
            tanh_f := 2046;
        ELSIF x = 7540 THEN
            tanh_f := 2046;
        ELSIF x = 7541 THEN
            tanh_f := 2046;
        ELSIF x = 7542 THEN
            tanh_f := 2046;
        ELSIF x = 7543 THEN
            tanh_f := 2046;
        ELSIF x = 7544 THEN
            tanh_f := 2046;
        ELSIF x = 7545 THEN
            tanh_f := 2046;
        ELSIF x = 7546 THEN
            tanh_f := 2046;
        ELSIF x = 7547 THEN
            tanh_f := 2046;
        ELSIF x = 7548 THEN
            tanh_f := 2046;
        ELSIF x = 7549 THEN
            tanh_f := 2046;
        ELSIF x = 7550 THEN
            tanh_f := 2046;
        ELSIF x = 7551 THEN
            tanh_f := 2046;
        ELSIF x = 7552 THEN
            tanh_f := 2046;
        ELSIF x = 7553 THEN
            tanh_f := 2046;
        ELSIF x = 7554 THEN
            tanh_f := 2046;
        ELSIF x = 7555 THEN
            tanh_f := 2046;
        ELSIF x = 7556 THEN
            tanh_f := 2046;
        ELSIF x = 7557 THEN
            tanh_f := 2046;
        ELSIF x = 7558 THEN
            tanh_f := 2046;
        ELSIF x = 7559 THEN
            tanh_f := 2046;
        ELSIF x = 7560 THEN
            tanh_f := 2046;
        ELSIF x = 7561 THEN
            tanh_f := 2046;
        ELSIF x = 7562 THEN
            tanh_f := 2046;
        ELSIF x = 7563 THEN
            tanh_f := 2046;
        ELSIF x = 7564 THEN
            tanh_f := 2046;
        ELSIF x = 7565 THEN
            tanh_f := 2046;
        ELSIF x = 7566 THEN
            tanh_f := 2046;
        ELSIF x = 7567 THEN
            tanh_f := 2046;
        ELSIF x = 7568 THEN
            tanh_f := 2046;
        ELSIF x = 7569 THEN
            tanh_f := 2046;
        ELSIF x = 7570 THEN
            tanh_f := 2046;
        ELSIF x = 7571 THEN
            tanh_f := 2046;
        ELSIF x = 7572 THEN
            tanh_f := 2046;
        ELSIF x = 7573 THEN
            tanh_f := 2046;
        ELSIF x = 7574 THEN
            tanh_f := 2046;
        ELSIF x = 7575 THEN
            tanh_f := 2046;
        ELSIF x = 7576 THEN
            tanh_f := 2046;
        ELSIF x = 7577 THEN
            tanh_f := 2046;
        ELSIF x = 7578 THEN
            tanh_f := 2046;
        ELSIF x = 7579 THEN
            tanh_f := 2046;
        ELSIF x = 7580 THEN
            tanh_f := 2046;
        ELSIF x = 7581 THEN
            tanh_f := 2046;
        ELSIF x = 7582 THEN
            tanh_f := 2046;
        ELSIF x = 7583 THEN
            tanh_f := 2046;
        ELSIF x = 7584 THEN
            tanh_f := 2046;
        ELSIF x = 7585 THEN
            tanh_f := 2046;
        ELSIF x = 7586 THEN
            tanh_f := 2046;
        ELSIF x = 7587 THEN
            tanh_f := 2046;
        ELSIF x = 7588 THEN
            tanh_f := 2046;
        ELSIF x = 7589 THEN
            tanh_f := 2046;
        ELSIF x = 7590 THEN
            tanh_f := 2046;
        ELSIF x = 7591 THEN
            tanh_f := 2046;
        ELSIF x = 7592 THEN
            tanh_f := 2046;
        ELSIF x = 7593 THEN
            tanh_f := 2046;
        ELSIF x = 7594 THEN
            tanh_f := 2046;
        ELSIF x = 7595 THEN
            tanh_f := 2046;
        ELSIF x = 7596 THEN
            tanh_f := 2046;
        ELSIF x = 7597 THEN
            tanh_f := 2046;
        ELSIF x = 7598 THEN
            tanh_f := 2046;
        ELSIF x = 7599 THEN
            tanh_f := 2046;
        ELSIF x = 7600 THEN
            tanh_f := 2046;
        ELSIF x = 7601 THEN
            tanh_f := 2046;
        ELSIF x = 7602 THEN
            tanh_f := 2046;
        ELSIF x = 7603 THEN
            tanh_f := 2046;
        ELSIF x = 7604 THEN
            tanh_f := 2046;
        ELSIF x = 7605 THEN
            tanh_f := 2046;
        ELSIF x = 7606 THEN
            tanh_f := 2046;
        ELSIF x = 7607 THEN
            tanh_f := 2046;
        ELSIF x = 7608 THEN
            tanh_f := 2046;
        ELSIF x = 7609 THEN
            tanh_f := 2046;
        ELSIF x = 7610 THEN
            tanh_f := 2046;
        ELSIF x = 7611 THEN
            tanh_f := 2046;
        ELSIF x = 7612 THEN
            tanh_f := 2046;
        ELSIF x = 7613 THEN
            tanh_f := 2046;
        ELSIF x = 7614 THEN
            tanh_f := 2046;
        ELSIF x = 7615 THEN
            tanh_f := 2046;
        ELSIF x = 7616 THEN
            tanh_f := 2046;
        ELSIF x = 7617 THEN
            tanh_f := 2046;
        ELSIF x = 7618 THEN
            tanh_f := 2046;
        ELSIF x = 7619 THEN
            tanh_f := 2046;
        ELSIF x = 7620 THEN
            tanh_f := 2046;
        ELSIF x = 7621 THEN
            tanh_f := 2046;
        ELSIF x = 7622 THEN
            tanh_f := 2046;
        ELSIF x = 7623 THEN
            tanh_f := 2046;
        ELSIF x = 7624 THEN
            tanh_f := 2046;
        ELSIF x = 7625 THEN
            tanh_f := 2046;
        ELSIF x = 7626 THEN
            tanh_f := 2046;
        ELSIF x = 7627 THEN
            tanh_f := 2046;
        ELSIF x = 7628 THEN
            tanh_f := 2046;
        ELSIF x = 7629 THEN
            tanh_f := 2046;
        ELSIF x = 7630 THEN
            tanh_f := 2046;
        ELSIF x = 7631 THEN
            tanh_f := 2046;
        ELSIF x = 7632 THEN
            tanh_f := 2046;
        ELSIF x = 7633 THEN
            tanh_f := 2046;
        ELSIF x = 7634 THEN
            tanh_f := 2046;
        ELSIF x = 7635 THEN
            tanh_f := 2046;
        ELSIF x = 7636 THEN
            tanh_f := 2046;
        ELSIF x = 7637 THEN
            tanh_f := 2046;
        ELSIF x = 7638 THEN
            tanh_f := 2046;
        ELSIF x = 7639 THEN
            tanh_f := 2046;
        ELSIF x = 7640 THEN
            tanh_f := 2046;
        ELSIF x = 7641 THEN
            tanh_f := 2046;
        ELSIF x = 7642 THEN
            tanh_f := 2046;
        ELSIF x = 7643 THEN
            tanh_f := 2046;
        ELSIF x = 7644 THEN
            tanh_f := 2046;
        ELSIF x = 7645 THEN
            tanh_f := 2046;
        ELSIF x = 7646 THEN
            tanh_f := 2046;
        ELSIF x = 7647 THEN
            tanh_f := 2046;
        ELSIF x = 7648 THEN
            tanh_f := 2046;
        ELSIF x = 7649 THEN
            tanh_f := 2046;
        ELSIF x = 7650 THEN
            tanh_f := 2046;
        ELSIF x = 7651 THEN
            tanh_f := 2046;
        ELSIF x = 7652 THEN
            tanh_f := 2046;
        ELSIF x = 7653 THEN
            tanh_f := 2046;
        ELSIF x = 7654 THEN
            tanh_f := 2046;
        ELSIF x = 7655 THEN
            tanh_f := 2046;
        ELSIF x = 7656 THEN
            tanh_f := 2046;
        ELSIF x = 7657 THEN
            tanh_f := 2046;
        ELSIF x = 7658 THEN
            tanh_f := 2046;
        ELSIF x = 7659 THEN
            tanh_f := 2046;
        ELSIF x = 7660 THEN
            tanh_f := 2046;
        ELSIF x = 7661 THEN
            tanh_f := 2046;
        ELSIF x = 7662 THEN
            tanh_f := 2046;
        ELSIF x = 7663 THEN
            tanh_f := 2046;
        ELSIF x = 7664 THEN
            tanh_f := 2046;
        ELSIF x = 7665 THEN
            tanh_f := 2046;
        ELSIF x = 7666 THEN
            tanh_f := 2046;
        ELSIF x = 7667 THEN
            tanh_f := 2046;
        ELSIF x = 7668 THEN
            tanh_f := 2046;
        ELSIF x = 7669 THEN
            tanh_f := 2046;
        ELSIF x = 7670 THEN
            tanh_f := 2046;
        ELSIF x = 7671 THEN
            tanh_f := 2046;
        ELSIF x = 7672 THEN
            tanh_f := 2046;
        ELSIF x = 7673 THEN
            tanh_f := 2046;
        ELSIF x = 7674 THEN
            tanh_f := 2046;
        ELSIF x = 7675 THEN
            tanh_f := 2046;
        ELSIF x = 7676 THEN
            tanh_f := 2046;
        ELSIF x = 7677 THEN
            tanh_f := 2046;
        ELSIF x = 7678 THEN
            tanh_f := 2046;
        ELSIF x = 7679 THEN
            tanh_f := 2046;
        ELSIF x = 7680 THEN
            tanh_f := 2046;
        ELSIF x = 7681 THEN
            tanh_f := 2046;
        ELSIF x = 7682 THEN
            tanh_f := 2046;
        ELSIF x = 7683 THEN
            tanh_f := 2046;
        ELSIF x = 7684 THEN
            tanh_f := 2046;
        ELSIF x = 7685 THEN
            tanh_f := 2046;
        ELSIF x = 7686 THEN
            tanh_f := 2046;
        ELSIF x = 7687 THEN
            tanh_f := 2046;
        ELSIF x = 7688 THEN
            tanh_f := 2046;
        ELSIF x = 7689 THEN
            tanh_f := 2046;
        ELSIF x = 7690 THEN
            tanh_f := 2046;
        ELSIF x = 7691 THEN
            tanh_f := 2046;
        ELSIF x = 7692 THEN
            tanh_f := 2046;
        ELSIF x = 7693 THEN
            tanh_f := 2046;
        ELSIF x = 7694 THEN
            tanh_f := 2046;
        ELSIF x = 7695 THEN
            tanh_f := 2046;
        ELSIF x = 7696 THEN
            tanh_f := 2046;
        ELSIF x = 7697 THEN
            tanh_f := 2046;
        ELSIF x = 7698 THEN
            tanh_f := 2046;
        ELSIF x = 7699 THEN
            tanh_f := 2046;
        ELSIF x = 7700 THEN
            tanh_f := 2046;
        ELSIF x = 7701 THEN
            tanh_f := 2046;
        ELSIF x = 7702 THEN
            tanh_f := 2046;
        ELSIF x = 7703 THEN
            tanh_f := 2046;
        ELSIF x = 7704 THEN
            tanh_f := 2046;
        ELSIF x = 7705 THEN
            tanh_f := 2046;
        ELSIF x = 7706 THEN
            tanh_f := 2046;
        ELSIF x = 7707 THEN
            tanh_f := 2046;
        ELSIF x = 7708 THEN
            tanh_f := 2046;
        ELSIF x = 7709 THEN
            tanh_f := 2046;
        ELSIF x = 7710 THEN
            tanh_f := 2046;
        ELSIF x = 7711 THEN
            tanh_f := 2046;
        ELSIF x = 7712 THEN
            tanh_f := 2046;
        ELSIF x = 7713 THEN
            tanh_f := 2046;
        ELSIF x = 7714 THEN
            tanh_f := 2046;
        ELSIF x = 7715 THEN
            tanh_f := 2046;
        ELSIF x = 7716 THEN
            tanh_f := 2046;
        ELSIF x = 7717 THEN
            tanh_f := 2046;
        ELSIF x = 7718 THEN
            tanh_f := 2046;
        ELSIF x = 7719 THEN
            tanh_f := 2046;
        ELSIF x = 7720 THEN
            tanh_f := 2046;
        ELSIF x = 7721 THEN
            tanh_f := 2046;
        ELSIF x = 7722 THEN
            tanh_f := 2046;
        ELSIF x = 7723 THEN
            tanh_f := 2046;
        ELSIF x = 7724 THEN
            tanh_f := 2046;
        ELSIF x = 7725 THEN
            tanh_f := 2046;
        ELSIF x = 7726 THEN
            tanh_f := 2046;
        ELSIF x = 7727 THEN
            tanh_f := 2046;
        ELSIF x = 7728 THEN
            tanh_f := 2046;
        ELSIF x = 7729 THEN
            tanh_f := 2046;
        ELSIF x = 7730 THEN
            tanh_f := 2046;
        ELSIF x = 7731 THEN
            tanh_f := 2046;
        ELSIF x = 7732 THEN
            tanh_f := 2046;
        ELSIF x = 7733 THEN
            tanh_f := 2046;
        ELSIF x = 7734 THEN
            tanh_f := 2046;
        ELSIF x = 7735 THEN
            tanh_f := 2046;
        ELSIF x = 7736 THEN
            tanh_f := 2046;
        ELSIF x = 7737 THEN
            tanh_f := 2046;
        ELSIF x = 7738 THEN
            tanh_f := 2046;
        ELSIF x = 7739 THEN
            tanh_f := 2046;
        ELSIF x = 7740 THEN
            tanh_f := 2046;
        ELSIF x = 7741 THEN
            tanh_f := 2046;
        ELSIF x = 7742 THEN
            tanh_f := 2046;
        ELSIF x = 7743 THEN
            tanh_f := 2046;
        ELSIF x = 7744 THEN
            tanh_f := 2046;
        ELSIF x = 7745 THEN
            tanh_f := 2046;
        ELSIF x = 7746 THEN
            tanh_f := 2046;
        ELSIF x = 7747 THEN
            tanh_f := 2046;
        ELSIF x = 7748 THEN
            tanh_f := 2046;
        ELSIF x = 7749 THEN
            tanh_f := 2046;
        ELSIF x = 7750 THEN
            tanh_f := 2046;
        ELSIF x = 7751 THEN
            tanh_f := 2046;
        ELSIF x = 7752 THEN
            tanh_f := 2046;
        ELSIF x = 7753 THEN
            tanh_f := 2046;
        ELSIF x = 7754 THEN
            tanh_f := 2046;
        ELSIF x = 7755 THEN
            tanh_f := 2046;
        ELSIF x = 7756 THEN
            tanh_f := 2046;
        ELSIF x = 7757 THEN
            tanh_f := 2046;
        ELSIF x = 7758 THEN
            tanh_f := 2046;
        ELSIF x = 7759 THEN
            tanh_f := 2046;
        ELSIF x = 7760 THEN
            tanh_f := 2046;
        ELSIF x = 7761 THEN
            tanh_f := 2046;
        ELSIF x = 7762 THEN
            tanh_f := 2046;
        ELSIF x = 7763 THEN
            tanh_f := 2046;
        ELSIF x = 7764 THEN
            tanh_f := 2046;
        ELSIF x = 7765 THEN
            tanh_f := 2046;
        ELSIF x = 7766 THEN
            tanh_f := 2046;
        ELSIF x = 7767 THEN
            tanh_f := 2046;
        ELSIF x = 7768 THEN
            tanh_f := 2046;
        ELSIF x = 7769 THEN
            tanh_f := 2046;
        ELSIF x = 7770 THEN
            tanh_f := 2046;
        ELSIF x = 7771 THEN
            tanh_f := 2046;
        ELSIF x = 7772 THEN
            tanh_f := 2046;
        ELSIF x = 7773 THEN
            tanh_f := 2046;
        ELSIF x = 7774 THEN
            tanh_f := 2046;
        ELSIF x = 7775 THEN
            tanh_f := 2046;
        ELSIF x = 7776 THEN
            tanh_f := 2046;
        ELSIF x = 7777 THEN
            tanh_f := 2046;
        ELSIF x = 7778 THEN
            tanh_f := 2046;
        ELSIF x = 7779 THEN
            tanh_f := 2046;
        ELSIF x = 7780 THEN
            tanh_f := 2046;
        ELSIF x = 7781 THEN
            tanh_f := 2046;
        ELSIF x = 7782 THEN
            tanh_f := 2046;
        ELSIF x = 7783 THEN
            tanh_f := 2046;
        ELSIF x = 7784 THEN
            tanh_f := 2046;
        ELSIF x = 7785 THEN
            tanh_f := 2046;
        ELSIF x = 7786 THEN
            tanh_f := 2046;
        ELSIF x = 7787 THEN
            tanh_f := 2046;
        ELSIF x = 7788 THEN
            tanh_f := 2046;
        ELSIF x = 7789 THEN
            tanh_f := 2046;
        ELSIF x = 7790 THEN
            tanh_f := 2046;
        ELSIF x = 7791 THEN
            tanh_f := 2046;
        ELSIF x = 7792 THEN
            tanh_f := 2046;
        ELSIF x = 7793 THEN
            tanh_f := 2046;
        ELSIF x = 7794 THEN
            tanh_f := 2046;
        ELSIF x = 7795 THEN
            tanh_f := 2046;
        ELSIF x = 7796 THEN
            tanh_f := 2046;
        ELSIF x = 7797 THEN
            tanh_f := 2046;
        ELSIF x = 7798 THEN
            tanh_f := 2046;
        ELSIF x = 7799 THEN
            tanh_f := 2046;
        ELSIF x = 7800 THEN
            tanh_f := 2046;
        ELSIF x = 7801 THEN
            tanh_f := 2046;
        ELSIF x = 7802 THEN
            tanh_f := 2046;
        ELSIF x = 7803 THEN
            tanh_f := 2046;
        ELSIF x = 7804 THEN
            tanh_f := 2046;
        ELSIF x = 7805 THEN
            tanh_f := 2046;
        ELSIF x = 7806 THEN
            tanh_f := 2046;
        ELSIF x = 7807 THEN
            tanh_f := 2046;
        ELSIF x = 7808 THEN
            tanh_f := 2046;
        ELSIF x = 7809 THEN
            tanh_f := 2046;
        ELSIF x = 7810 THEN
            tanh_f := 2046;
        ELSIF x = 7811 THEN
            tanh_f := 2046;
        ELSIF x = 7812 THEN
            tanh_f := 2046;
        ELSIF x = 7813 THEN
            tanh_f := 2046;
        ELSIF x = 7814 THEN
            tanh_f := 2046;
        ELSIF x = 7815 THEN
            tanh_f := 2046;
        ELSIF x = 7816 THEN
            tanh_f := 2046;
        ELSIF x = 7817 THEN
            tanh_f := 2046;
        ELSIF x = 7818 THEN
            tanh_f := 2046;
        ELSIF x = 7819 THEN
            tanh_f := 2046;
        ELSIF x = 7820 THEN
            tanh_f := 2046;
        ELSIF x = 7821 THEN
            tanh_f := 2046;
        ELSIF x = 7822 THEN
            tanh_f := 2046;
        ELSIF x = 7823 THEN
            tanh_f := 2046;
        ELSIF x = 7824 THEN
            tanh_f := 2046;
        ELSIF x = 7825 THEN
            tanh_f := 2046;
        ELSIF x = 7826 THEN
            tanh_f := 2046;
        ELSIF x = 7827 THEN
            tanh_f := 2046;
        ELSIF x = 7828 THEN
            tanh_f := 2046;
        ELSIF x = 7829 THEN
            tanh_f := 2046;
        ELSIF x = 7830 THEN
            tanh_f := 2046;
        ELSIF x = 7831 THEN
            tanh_f := 2046;
        ELSIF x = 7832 THEN
            tanh_f := 2046;
        ELSIF x = 7833 THEN
            tanh_f := 2046;
        ELSIF x = 7834 THEN
            tanh_f := 2046;
        ELSIF x = 7835 THEN
            tanh_f := 2046;
        ELSIF x = 7836 THEN
            tanh_f := 2046;
        ELSIF x = 7837 THEN
            tanh_f := 2046;
        ELSIF x = 7838 THEN
            tanh_f := 2046;
        ELSIF x = 7839 THEN
            tanh_f := 2046;
        ELSIF x = 7840 THEN
            tanh_f := 2046;
        ELSIF x = 7841 THEN
            tanh_f := 2046;
        ELSIF x = 7842 THEN
            tanh_f := 2046;
        ELSIF x = 7843 THEN
            tanh_f := 2046;
        ELSIF x = 7844 THEN
            tanh_f := 2046;
        ELSIF x = 7845 THEN
            tanh_f := 2046;
        ELSIF x = 7846 THEN
            tanh_f := 2046;
        ELSIF x = 7847 THEN
            tanh_f := 2046;
        ELSIF x = 7848 THEN
            tanh_f := 2046;
        ELSIF x = 7849 THEN
            tanh_f := 2046;
        ELSIF x = 7850 THEN
            tanh_f := 2046;
        ELSIF x = 7851 THEN
            tanh_f := 2046;
        ELSIF x = 7852 THEN
            tanh_f := 2046;
        ELSIF x = 7853 THEN
            tanh_f := 2046;
        ELSIF x = 7854 THEN
            tanh_f := 2046;
        ELSIF x = 7855 THEN
            tanh_f := 2046;
        ELSIF x = 7856 THEN
            tanh_f := 2046;
        ELSIF x = 7857 THEN
            tanh_f := 2046;
        ELSIF x = 7858 THEN
            tanh_f := 2046;
        ELSIF x = 7859 THEN
            tanh_f := 2046;
        ELSIF x = 7860 THEN
            tanh_f := 2046;
        ELSIF x = 7861 THEN
            tanh_f := 2046;
        ELSIF x = 7862 THEN
            tanh_f := 2046;
        ELSIF x = 7863 THEN
            tanh_f := 2046;
        ELSIF x = 7864 THEN
            tanh_f := 2046;
        ELSIF x = 7865 THEN
            tanh_f := 2046;
        ELSIF x = 7866 THEN
            tanh_f := 2046;
        ELSIF x = 7867 THEN
            tanh_f := 2046;
        ELSIF x = 7868 THEN
            tanh_f := 2046;
        ELSIF x = 7869 THEN
            tanh_f := 2046;
        ELSIF x = 7870 THEN
            tanh_f := 2046;
        ELSIF x = 7871 THEN
            tanh_f := 2046;
        ELSIF x = 7872 THEN
            tanh_f := 2046;
        ELSIF x = 7873 THEN
            tanh_f := 2046;
        ELSIF x = 7874 THEN
            tanh_f := 2046;
        ELSIF x = 7875 THEN
            tanh_f := 2046;
        ELSIF x = 7876 THEN
            tanh_f := 2046;
        ELSIF x = 7877 THEN
            tanh_f := 2046;
        ELSIF x = 7878 THEN
            tanh_f := 2046;
        ELSIF x = 7879 THEN
            tanh_f := 2046;
        ELSIF x = 7880 THEN
            tanh_f := 2046;
        ELSIF x = 7881 THEN
            tanh_f := 2046;
        ELSIF x = 7882 THEN
            tanh_f := 2046;
        ELSIF x = 7883 THEN
            tanh_f := 2046;
        ELSIF x = 7884 THEN
            tanh_f := 2046;
        ELSIF x = 7885 THEN
            tanh_f := 2046;
        ELSIF x = 7886 THEN
            tanh_f := 2046;
        ELSIF x = 7887 THEN
            tanh_f := 2046;
        ELSIF x = 7888 THEN
            tanh_f := 2046;
        ELSIF x = 7889 THEN
            tanh_f := 2046;
        ELSIF x = 7890 THEN
            tanh_f := 2046;
        ELSIF x = 7891 THEN
            tanh_f := 2046;
        ELSIF x = 7892 THEN
            tanh_f := 2046;
        ELSIF x = 7893 THEN
            tanh_f := 2046;
        ELSIF x = 7894 THEN
            tanh_f := 2046;
        ELSIF x = 7895 THEN
            tanh_f := 2046;
        ELSIF x = 7896 THEN
            tanh_f := 2046;
        ELSIF x = 7897 THEN
            tanh_f := 2046;
        ELSIF x = 7898 THEN
            tanh_f := 2046;
        ELSIF x = 7899 THEN
            tanh_f := 2046;
        ELSIF x = 7900 THEN
            tanh_f := 2046;
        ELSIF x = 7901 THEN
            tanh_f := 2046;
        ELSIF x = 7902 THEN
            tanh_f := 2046;
        ELSIF x = 7903 THEN
            tanh_f := 2046;
        ELSIF x = 7904 THEN
            tanh_f := 2046;
        ELSIF x = 7905 THEN
            tanh_f := 2046;
        ELSIF x = 7906 THEN
            tanh_f := 2046;
        ELSIF x = 7907 THEN
            tanh_f := 2046;
        ELSIF x = 7908 THEN
            tanh_f := 2046;
        ELSIF x = 7909 THEN
            tanh_f := 2046;
        ELSIF x = 7910 THEN
            tanh_f := 2046;
        ELSIF x = 7911 THEN
            tanh_f := 2046;
        ELSIF x = 7912 THEN
            tanh_f := 2046;
        ELSIF x = 7913 THEN
            tanh_f := 2046;
        ELSIF x = 7914 THEN
            tanh_f := 2046;
        ELSIF x = 7915 THEN
            tanh_f := 2046;
        ELSIF x = 7916 THEN
            tanh_f := 2046;
        ELSIF x = 7917 THEN
            tanh_f := 2046;
        ELSIF x = 7918 THEN
            tanh_f := 2046;
        ELSIF x = 7919 THEN
            tanh_f := 2046;
        ELSIF x = 7920 THEN
            tanh_f := 2046;
        ELSIF x = 7921 THEN
            tanh_f := 2046;
        ELSIF x = 7922 THEN
            tanh_f := 2046;
        ELSIF x = 7923 THEN
            tanh_f := 2046;
        ELSIF x = 7924 THEN
            tanh_f := 2046;
        ELSIF x = 7925 THEN
            tanh_f := 2046;
        ELSIF x = 7926 THEN
            tanh_f := 2046;
        ELSIF x = 7927 THEN
            tanh_f := 2046;
        ELSIF x = 7928 THEN
            tanh_f := 2046;
        ELSIF x = 7929 THEN
            tanh_f := 2046;
        ELSIF x = 7930 THEN
            tanh_f := 2046;
        ELSIF x = 7931 THEN
            tanh_f := 2046;
        ELSIF x = 7932 THEN
            tanh_f := 2046;
        ELSIF x = 7933 THEN
            tanh_f := 2046;
        ELSIF x = 7934 THEN
            tanh_f := 2046;
        ELSIF x = 7935 THEN
            tanh_f := 2046;
        ELSIF x = 7936 THEN
            tanh_f := 2046;
        ELSIF x = 7937 THEN
            tanh_f := 2046;
        ELSIF x = 7938 THEN
            tanh_f := 2046;
        ELSIF x = 7939 THEN
            tanh_f := 2046;
        ELSIF x = 7940 THEN
            tanh_f := 2046;
        ELSIF x = 7941 THEN
            tanh_f := 2046;
        ELSIF x = 7942 THEN
            tanh_f := 2046;
        ELSIF x = 7943 THEN
            tanh_f := 2046;
        ELSIF x = 7944 THEN
            tanh_f := 2046;
        ELSIF x = 7945 THEN
            tanh_f := 2046;
        ELSIF x = 7946 THEN
            tanh_f := 2046;
        ELSIF x = 7947 THEN
            tanh_f := 2046;
        ELSIF x = 7948 THEN
            tanh_f := 2046;
        ELSIF x = 7949 THEN
            tanh_f := 2046;
        ELSIF x = 7950 THEN
            tanh_f := 2046;
        ELSIF x = 7951 THEN
            tanh_f := 2046;
        ELSIF x = 7952 THEN
            tanh_f := 2046;
        ELSIF x = 7953 THEN
            tanh_f := 2046;
        ELSIF x = 7954 THEN
            tanh_f := 2046;
        ELSIF x = 7955 THEN
            tanh_f := 2046;
        ELSIF x = 7956 THEN
            tanh_f := 2046;
        ELSIF x = 7957 THEN
            tanh_f := 2046;
        ELSIF x = 7958 THEN
            tanh_f := 2046;
        ELSIF x = 7959 THEN
            tanh_f := 2046;
        ELSIF x = 7960 THEN
            tanh_f := 2046;
        ELSIF x = 7961 THEN
            tanh_f := 2046;
        ELSIF x = 7962 THEN
            tanh_f := 2046;
        ELSIF x = 7963 THEN
            tanh_f := 2046;
        ELSIF x = 7964 THEN
            tanh_f := 2046;
        ELSIF x = 7965 THEN
            tanh_f := 2046;
        ELSIF x = 7966 THEN
            tanh_f := 2046;
        ELSIF x = 7967 THEN
            tanh_f := 2046;
        ELSIF x = 7968 THEN
            tanh_f := 2046;
        ELSIF x = 7969 THEN
            tanh_f := 2046;
        ELSIF x = 7970 THEN
            tanh_f := 2046;
        ELSIF x = 7971 THEN
            tanh_f := 2046;
        ELSIF x = 7972 THEN
            tanh_f := 2046;
        ELSIF x = 7973 THEN
            tanh_f := 2046;
        ELSIF x = 7974 THEN
            tanh_f := 2046;
        ELSIF x = 7975 THEN
            tanh_f := 2046;
        ELSIF x = 7976 THEN
            tanh_f := 2046;
        ELSIF x = 7977 THEN
            tanh_f := 2046;
        ELSIF x = 7978 THEN
            tanh_f := 2046;
        ELSIF x = 7979 THEN
            tanh_f := 2046;
        ELSIF x = 7980 THEN
            tanh_f := 2046;
        ELSIF x = 7981 THEN
            tanh_f := 2046;
        ELSIF x = 7982 THEN
            tanh_f := 2046;
        ELSIF x = 7983 THEN
            tanh_f := 2046;
        ELSIF x = 7984 THEN
            tanh_f := 2046;
        ELSIF x = 7985 THEN
            tanh_f := 2046;
        ELSIF x = 7986 THEN
            tanh_f := 2046;
        ELSIF x = 7987 THEN
            tanh_f := 2046;
        ELSIF x = 7988 THEN
            tanh_f := 2046;
        ELSIF x = 7989 THEN
            tanh_f := 2046;
        ELSIF x = 7990 THEN
            tanh_f := 2046;
        ELSIF x = 7991 THEN
            tanh_f := 2046;
        ELSIF x = 7992 THEN
            tanh_f := 2046;
        ELSIF x = 7993 THEN
            tanh_f := 2046;
        ELSIF x = 7994 THEN
            tanh_f := 2046;
        ELSIF x = 7995 THEN
            tanh_f := 2046;
        ELSIF x = 7996 THEN
            tanh_f := 2046;
        ELSIF x = 7997 THEN
            tanh_f := 2046;
        ELSIF x = 7998 THEN
            tanh_f := 2046;
        ELSIF x = 7999 THEN
            tanh_f := 2046;
        ELSIF x = 8000 THEN
            tanh_f := 2046;
        ELSIF x = 8001 THEN
            tanh_f := 2046;
        ELSIF x = 8002 THEN
            tanh_f := 2046;
        ELSIF x = 8003 THEN
            tanh_f := 2046;
        ELSIF x = 8004 THEN
            tanh_f := 2046;
        ELSIF x = 8005 THEN
            tanh_f := 2046;
        ELSIF x = 8006 THEN
            tanh_f := 2046;
        ELSIF x = 8007 THEN
            tanh_f := 2046;
        ELSIF x = 8008 THEN
            tanh_f := 2046;
        ELSIF x = 8009 THEN
            tanh_f := 2046;
        ELSIF x = 8010 THEN
            tanh_f := 2046;
        ELSIF x = 8011 THEN
            tanh_f := 2046;
        ELSIF x = 8012 THEN
            tanh_f := 2046;
        ELSIF x = 8013 THEN
            tanh_f := 2046;
        ELSIF x = 8014 THEN
            tanh_f := 2046;
        ELSIF x = 8015 THEN
            tanh_f := 2046;
        ELSIF x = 8016 THEN
            tanh_f := 2046;
        ELSIF x = 8017 THEN
            tanh_f := 2046;
        ELSIF x = 8018 THEN
            tanh_f := 2046;
        ELSIF x = 8019 THEN
            tanh_f := 2046;
        ELSIF x = 8020 THEN
            tanh_f := 2046;
        ELSIF x = 8021 THEN
            tanh_f := 2046;
        ELSIF x = 8022 THEN
            tanh_f := 2046;
        ELSIF x = 8023 THEN
            tanh_f := 2046;
        ELSIF x = 8024 THEN
            tanh_f := 2046;
        ELSIF x = 8025 THEN
            tanh_f := 2046;
        ELSIF x = 8026 THEN
            tanh_f := 2046;
        ELSIF x = 8027 THEN
            tanh_f := 2046;
        ELSIF x = 8028 THEN
            tanh_f := 2046;
        ELSIF x = 8029 THEN
            tanh_f := 2046;
        ELSIF x = 8030 THEN
            tanh_f := 2046;
        ELSIF x = 8031 THEN
            tanh_f := 2046;
        ELSIF x = 8032 THEN
            tanh_f := 2046;
        ELSIF x = 8033 THEN
            tanh_f := 2046;
        ELSIF x = 8034 THEN
            tanh_f := 2046;
        ELSIF x = 8035 THEN
            tanh_f := 2046;
        ELSIF x = 8036 THEN
            tanh_f := 2046;
        ELSIF x = 8037 THEN
            tanh_f := 2046;
        ELSIF x = 8038 THEN
            tanh_f := 2046;
        ELSIF x = 8039 THEN
            tanh_f := 2046;
        ELSIF x = 8040 THEN
            tanh_f := 2046;
        ELSIF x = 8041 THEN
            tanh_f := 2046;
        ELSIF x = 8042 THEN
            tanh_f := 2046;
        ELSIF x = 8043 THEN
            tanh_f := 2046;
        ELSIF x = 8044 THEN
            tanh_f := 2046;
        ELSIF x = 8045 THEN
            tanh_f := 2046;
        ELSIF x = 8046 THEN
            tanh_f := 2046;
        ELSIF x = 8047 THEN
            tanh_f := 2046;
        ELSIF x = 8048 THEN
            tanh_f := 2046;
        ELSIF x = 8049 THEN
            tanh_f := 2046;
        ELSIF x = 8050 THEN
            tanh_f := 2046;
        ELSIF x = 8051 THEN
            tanh_f := 2046;
        ELSIF x = 8052 THEN
            tanh_f := 2046;
        ELSIF x = 8053 THEN
            tanh_f := 2046;
        ELSIF x = 8054 THEN
            tanh_f := 2046;
        ELSIF x = 8055 THEN
            tanh_f := 2046;
        ELSIF x = 8056 THEN
            tanh_f := 2046;
        ELSIF x = 8057 THEN
            tanh_f := 2046;
        ELSIF x = 8058 THEN
            tanh_f := 2046;
        ELSIF x = 8059 THEN
            tanh_f := 2046;
        ELSIF x = 8060 THEN
            tanh_f := 2046;
        ELSIF x = 8061 THEN
            tanh_f := 2046;
        ELSIF x = 8062 THEN
            tanh_f := 2046;
        ELSIF x = 8063 THEN
            tanh_f := 2046;
        ELSIF x = 8064 THEN
            tanh_f := 2046;
        ELSIF x = 8065 THEN
            tanh_f := 2046;
        ELSIF x = 8066 THEN
            tanh_f := 2046;
        ELSIF x = 8067 THEN
            tanh_f := 2046;
        ELSIF x = 8068 THEN
            tanh_f := 2046;
        ELSIF x = 8069 THEN
            tanh_f := 2046;
        ELSIF x = 8070 THEN
            tanh_f := 2046;
        ELSIF x = 8071 THEN
            tanh_f := 2046;
        ELSIF x = 8072 THEN
            tanh_f := 2046;
        ELSIF x = 8073 THEN
            tanh_f := 2046;
        ELSIF x = 8074 THEN
            tanh_f := 2046;
        ELSIF x = 8075 THEN
            tanh_f := 2046;
        ELSIF x = 8076 THEN
            tanh_f := 2046;
        ELSIF x = 8077 THEN
            tanh_f := 2046;
        ELSIF x = 8078 THEN
            tanh_f := 2046;
        ELSIF x = 8079 THEN
            tanh_f := 2046;
        ELSIF x = 8080 THEN
            tanh_f := 2046;
        ELSIF x = 8081 THEN
            tanh_f := 2046;
        ELSIF x = 8082 THEN
            tanh_f := 2046;
        ELSIF x = 8083 THEN
            tanh_f := 2046;
        ELSIF x = 8084 THEN
            tanh_f := 2046;
        ELSIF x = 8085 THEN
            tanh_f := 2046;
        ELSIF x = 8086 THEN
            tanh_f := 2046;
        ELSIF x = 8087 THEN
            tanh_f := 2046;
        ELSIF x = 8088 THEN
            tanh_f := 2046;
        ELSIF x = 8089 THEN
            tanh_f := 2046;
        ELSIF x = 8090 THEN
            tanh_f := 2046;
        ELSIF x = 8091 THEN
            tanh_f := 2046;
        ELSIF x = 8092 THEN
            tanh_f := 2046;
        ELSIF x = 8093 THEN
            tanh_f := 2046;
        ELSIF x = 8094 THEN
            tanh_f := 2046;
        ELSIF x = 8095 THEN
            tanh_f := 2046;
        ELSIF x = 8096 THEN
            tanh_f := 2046;
        ELSIF x = 8097 THEN
            tanh_f := 2046;
        ELSIF x = 8098 THEN
            tanh_f := 2046;
        ELSIF x = 8099 THEN
            tanh_f := 2046;
        ELSIF x = 8100 THEN
            tanh_f := 2046;
        ELSIF x = 8101 THEN
            tanh_f := 2046;
        ELSIF x = 8102 THEN
            tanh_f := 2046;
        ELSIF x = 8103 THEN
            tanh_f := 2046;
        ELSIF x = 8104 THEN
            tanh_f := 2046;
        ELSIF x = 8105 THEN
            tanh_f := 2046;
        ELSIF x = 8106 THEN
            tanh_f := 2046;
        ELSIF x = 8107 THEN
            tanh_f := 2046;
        ELSIF x = 8108 THEN
            tanh_f := 2046;
        ELSIF x = 8109 THEN
            tanh_f := 2046;
        ELSIF x = 8110 THEN
            tanh_f := 2046;
        ELSIF x = 8111 THEN
            tanh_f := 2046;
        ELSIF x = 8112 THEN
            tanh_f := 2046;
        ELSIF x = 8113 THEN
            tanh_f := 2046;
        ELSIF x = 8114 THEN
            tanh_f := 2046;
        ELSIF x = 8115 THEN
            tanh_f := 2046;
        ELSIF x = 8116 THEN
            tanh_f := 2046;
        ELSIF x = 8117 THEN
            tanh_f := 2046;
        ELSIF x = 8118 THEN
            tanh_f := 2046;
        ELSIF x = 8119 THEN
            tanh_f := 2046;
        ELSIF x = 8120 THEN
            tanh_f := 2046;
        ELSIF x = 8121 THEN
            tanh_f := 2046;
        ELSIF x = 8122 THEN
            tanh_f := 2046;
        ELSIF x = 8123 THEN
            tanh_f := 2046;
        ELSIF x = 8124 THEN
            tanh_f := 2046;
        ELSIF x = 8125 THEN
            tanh_f := 2046;
        ELSIF x = 8126 THEN
            tanh_f := 2046;
        ELSIF x = 8127 THEN
            tanh_f := 2046;
        ELSIF x = 8128 THEN
            tanh_f := 2046;
        ELSIF x = 8129 THEN
            tanh_f := 2046;
        ELSIF x = 8130 THEN
            tanh_f := 2046;
        ELSIF x = 8131 THEN
            tanh_f := 2046;
        ELSIF x = 8132 THEN
            tanh_f := 2046;
        ELSIF x = 8133 THEN
            tanh_f := 2046;
        ELSIF x = 8134 THEN
            tanh_f := 2046;
        ELSIF x = 8135 THEN
            tanh_f := 2046;
        ELSIF x = 8136 THEN
            tanh_f := 2046;
        ELSIF x = 8137 THEN
            tanh_f := 2046;
        ELSIF x = 8138 THEN
            tanh_f := 2046;
        ELSIF x = 8139 THEN
            tanh_f := 2046;
        ELSIF x = 8140 THEN
            tanh_f := 2046;
        ELSIF x = 8141 THEN
            tanh_f := 2046;
        ELSIF x = 8142 THEN
            tanh_f := 2046;
        ELSIF x = 8143 THEN
            tanh_f := 2046;
        ELSIF x = 8144 THEN
            tanh_f := 2046;
        ELSIF x = 8145 THEN
            tanh_f := 2046;
        ELSIF x = 8146 THEN
            tanh_f := 2046;
        ELSIF x = 8147 THEN
            tanh_f := 2046;
        ELSIF x = 8148 THEN
            tanh_f := 2046;
        ELSIF x = 8149 THEN
            tanh_f := 2046;
        ELSIF x = 8150 THEN
            tanh_f := 2046;
        ELSIF x = 8151 THEN
            tanh_f := 2046;
        ELSIF x = 8152 THEN
            tanh_f := 2046;
        ELSIF x = 8153 THEN
            tanh_f := 2046;
        ELSIF x = 8154 THEN
            tanh_f := 2046;
        ELSIF x = 8155 THEN
            tanh_f := 2046;
        ELSIF x = 8156 THEN
            tanh_f := 2046;
        ELSIF x = 8157 THEN
            tanh_f := 2046;
        ELSIF x = 8158 THEN
            tanh_f := 2046;
        ELSIF x = 8159 THEN
            tanh_f := 2046;
        ELSIF x = 8160 THEN
            tanh_f := 2046;
        ELSIF x = 8161 THEN
            tanh_f := 2046;
        ELSIF x = 8162 THEN
            tanh_f := 2046;
        ELSIF x = 8163 THEN
            tanh_f := 2046;
        ELSIF x = 8164 THEN
            tanh_f := 2046;
        ELSIF x = 8165 THEN
            tanh_f := 2046;
        ELSIF x = 8166 THEN
            tanh_f := 2046;
        ELSIF x = 8167 THEN
            tanh_f := 2046;
        ELSIF x = 8168 THEN
            tanh_f := 2046;
        ELSIF x = 8169 THEN
            tanh_f := 2046;
        ELSIF x = 8170 THEN
            tanh_f := 2046;
        ELSIF x = 8171 THEN
            tanh_f := 2046;
        ELSIF x = 8172 THEN
            tanh_f := 2046;
        ELSIF x = 8173 THEN
            tanh_f := 2046;
        ELSIF x = 8174 THEN
            tanh_f := 2046;
        ELSIF x = 8175 THEN
            tanh_f := 2046;
        ELSIF x = 8176 THEN
            tanh_f := 2046;
        ELSIF x = 8177 THEN
            tanh_f := 2046;
        ELSIF x = 8178 THEN
            tanh_f := 2046;
        ELSIF x = 8179 THEN
            tanh_f := 2046;
        ELSIF x = 8180 THEN
            tanh_f := 2046;
        ELSIF x = 8181 THEN
            tanh_f := 2046;
        ELSIF x = 8182 THEN
            tanh_f := 2046;
        ELSIF x = 8183 THEN
            tanh_f := 2046;
        ELSIF x = 8184 THEN
            tanh_f := 2046;
        ELSIF x = 8185 THEN
            tanh_f := 2046;
        ELSIF x = 8186 THEN
            tanh_f := 2046;
        ELSIF x = 8187 THEN
            tanh_f := 2046;
        ELSIF x = 8188 THEN
            tanh_f := 2046;
        ELSIF x = 8189 THEN
            tanh_f := 2046;
        ELSIF x = 8190 THEN
            tanh_f := 2046;
        ELSIF x = 8191 THEN
            tanh_f := 2046;
        ELSIF x = 8192 THEN
            tanh_f := 2046;
        ELSIF x = 8193 THEN
            tanh_f := 2046;
        ELSIF x = 8194 THEN
            tanh_f := 2046;
        ELSIF x = 8195 THEN
            tanh_f := 2046;
        ELSIF x = 8196 THEN
            tanh_f := 2046;
        ELSIF x = 8197 THEN
            tanh_f := 2046;
        ELSIF x = 8198 THEN
            tanh_f := 2046;
        ELSIF x = 8199 THEN
            tanh_f := 2046;
        ELSIF x = 8200 THEN
            tanh_f := 2046;
        ELSIF x = 8201 THEN
            tanh_f := 2046;
        ELSIF x = 8202 THEN
            tanh_f := 2046;
        ELSIF x = 8203 THEN
            tanh_f := 2046;
        ELSIF x = 8204 THEN
            tanh_f := 2046;
        ELSIF x = 8205 THEN
            tanh_f := 2046;
        ELSIF x = 8206 THEN
            tanh_f := 2046;
        ELSIF x = 8207 THEN
            tanh_f := 2046;
        ELSIF x = 8208 THEN
            tanh_f := 2046;
        ELSIF x = 8209 THEN
            tanh_f := 2046;
        ELSIF x = 8210 THEN
            tanh_f := 2046;
        ELSIF x = 8211 THEN
            tanh_f := 2046;
        ELSIF x = 8212 THEN
            tanh_f := 2046;
        ELSIF x = 8213 THEN
            tanh_f := 2046;
        ELSIF x = 8214 THEN
            tanh_f := 2046;
        ELSIF x = 8215 THEN
            tanh_f := 2046;
        ELSIF x = 8216 THEN
            tanh_f := 2046;
        ELSIF x = 8217 THEN
            tanh_f := 2046;
        ELSIF x = 8218 THEN
            tanh_f := 2046;
        ELSIF x = 8219 THEN
            tanh_f := 2046;
        ELSIF x = 8220 THEN
            tanh_f := 2046;
        ELSIF x = 8221 THEN
            tanh_f := 2046;
        ELSIF x = 8222 THEN
            tanh_f := 2046;
        ELSIF x = 8223 THEN
            tanh_f := 2046;
        ELSIF x = 8224 THEN
            tanh_f := 2046;
        ELSIF x = 8225 THEN
            tanh_f := 2046;
        ELSIF x = 8226 THEN
            tanh_f := 2046;
        ELSIF x = 8227 THEN
            tanh_f := 2046;
        ELSIF x = 8228 THEN
            tanh_f := 2046;
        ELSIF x = 8229 THEN
            tanh_f := 2046;
        ELSIF x = 8230 THEN
            tanh_f := 2046;
        ELSIF x = 8231 THEN
            tanh_f := 2046;
        ELSIF x = 8232 THEN
            tanh_f := 2046;
        ELSIF x = 8233 THEN
            tanh_f := 2046;
        ELSIF x = 8234 THEN
            tanh_f := 2046;
        ELSIF x = 8235 THEN
            tanh_f := 2046;
        ELSIF x = 8236 THEN
            tanh_f := 2046;
        ELSIF x = 8237 THEN
            tanh_f := 2046;
        ELSIF x = 8238 THEN
            tanh_f := 2046;
        ELSIF x = 8239 THEN
            tanh_f := 2046;
        ELSIF x = 8240 THEN
            tanh_f := 2046;
        ELSIF x = 8241 THEN
            tanh_f := 2046;
        ELSIF x = 8242 THEN
            tanh_f := 2046;
        ELSIF x = 8243 THEN
            tanh_f := 2046;
        ELSIF x = 8244 THEN
            tanh_f := 2046;
        ELSIF x = 8245 THEN
            tanh_f := 2046;
        ELSIF x = 8246 THEN
            tanh_f := 2046;
        ELSIF x = 8247 THEN
            tanh_f := 2046;
        ELSIF x = 8248 THEN
            tanh_f := 2046;
        ELSIF x = 8249 THEN
            tanh_f := 2046;
        ELSIF x = 8250 THEN
            tanh_f := 2046;
        ELSIF x = 8251 THEN
            tanh_f := 2046;
        ELSIF x = 8252 THEN
            tanh_f := 2046;
        ELSIF x = 8253 THEN
            tanh_f := 2046;
        ELSIF x = 8254 THEN
            tanh_f := 2046;
        ELSIF x = 8255 THEN
            tanh_f := 2046;
        ELSIF x = 8256 THEN
            tanh_f := 2046;
        ELSIF x = 8257 THEN
            tanh_f := 2046;
        ELSIF x = 8258 THEN
            tanh_f := 2046;
        ELSIF x = 8259 THEN
            tanh_f := 2046;
        ELSIF x = 8260 THEN
            tanh_f := 2046;
        ELSIF x = 8261 THEN
            tanh_f := 2046;
        ELSIF x = 8262 THEN
            tanh_f := 2046;
        ELSIF x = 8263 THEN
            tanh_f := 2046;
        ELSIF x = 8264 THEN
            tanh_f := 2046;
        ELSIF x = 8265 THEN
            tanh_f := 2046;
        ELSIF x = 8266 THEN
            tanh_f := 2046;
        ELSIF x = 8267 THEN
            tanh_f := 2046;
        ELSIF x = 8268 THEN
            tanh_f := 2046;
        ELSIF x = 8269 THEN
            tanh_f := 2046;
        ELSIF x = 8270 THEN
            tanh_f := 2046;
        ELSIF x = 8271 THEN
            tanh_f := 2046;
        ELSIF x = 8272 THEN
            tanh_f := 2046;
        ELSIF x = 8273 THEN
            tanh_f := 2046;
        ELSIF x = 8274 THEN
            tanh_f := 2046;
        ELSIF x = 8275 THEN
            tanh_f := 2046;
        ELSIF x = 8276 THEN
            tanh_f := 2046;
        ELSIF x = 8277 THEN
            tanh_f := 2046;
        ELSIF x = 8278 THEN
            tanh_f := 2046;
        ELSIF x = 8279 THEN
            tanh_f := 2046;
        ELSIF x = 8280 THEN
            tanh_f := 2046;
        ELSIF x = 8281 THEN
            tanh_f := 2046;
        ELSIF x = 8282 THEN
            tanh_f := 2046;
        ELSIF x = 8283 THEN
            tanh_f := 2046;
        ELSIF x = 8284 THEN
            tanh_f := 2046;
        ELSIF x = 8285 THEN
            tanh_f := 2046;
        ELSIF x = 8286 THEN
            tanh_f := 2046;
        ELSIF x = 8287 THEN
            tanh_f := 2046;
        ELSIF x = 8288 THEN
            tanh_f := 2046;
        ELSIF x = 8289 THEN
            tanh_f := 2046;
        ELSIF x = 8290 THEN
            tanh_f := 2046;
        ELSIF x = 8291 THEN
            tanh_f := 2046;
        ELSIF x = 8292 THEN
            tanh_f := 2046;
        ELSIF x = 8293 THEN
            tanh_f := 2046;
        ELSIF x = 8294 THEN
            tanh_f := 2046;
        ELSIF x = 8295 THEN
            tanh_f := 2046;
        ELSIF x = 8296 THEN
            tanh_f := 2046;
        ELSIF x = 8297 THEN
            tanh_f := 2046;
        ELSIF x = 8298 THEN
            tanh_f := 2046;
        ELSIF x = 8299 THEN
            tanh_f := 2046;
        ELSIF x = 8300 THEN
            tanh_f := 2046;
        ELSIF x = 8301 THEN
            tanh_f := 2046;
        ELSIF x = 8302 THEN
            tanh_f := 2046;
        ELSIF x = 8303 THEN
            tanh_f := 2046;
        ELSIF x = 8304 THEN
            tanh_f := 2046;
        ELSIF x = 8305 THEN
            tanh_f := 2046;
        ELSIF x = 8306 THEN
            tanh_f := 2046;
        ELSIF x = 8307 THEN
            tanh_f := 2046;
        ELSIF x = 8308 THEN
            tanh_f := 2046;
        ELSIF x = 8309 THEN
            tanh_f := 2046;
        ELSIF x = 8310 THEN
            tanh_f := 2046;
        ELSIF x = 8311 THEN
            tanh_f := 2046;
        ELSIF x = 8312 THEN
            tanh_f := 2046;
        ELSIF x = 8313 THEN
            tanh_f := 2046;
        ELSIF x = 8314 THEN
            tanh_f := 2046;
        ELSIF x = 8315 THEN
            tanh_f := 2046;
        ELSIF x = 8316 THEN
            tanh_f := 2046;
        ELSIF x = 8317 THEN
            tanh_f := 2046;
        ELSIF x = 8318 THEN
            tanh_f := 2046;
        ELSIF x = 8319 THEN
            tanh_f := 2046;
        ELSIF x = 8320 THEN
            tanh_f := 2046;
        ELSIF x = 8321 THEN
            tanh_f := 2046;
        ELSIF x = 8322 THEN
            tanh_f := 2046;
        ELSIF x = 8323 THEN
            tanh_f := 2046;
        ELSIF x = 8324 THEN
            tanh_f := 2046;
        ELSIF x = 8325 THEN
            tanh_f := 2046;
        ELSIF x = 8326 THEN
            tanh_f := 2046;
        ELSIF x = 8327 THEN
            tanh_f := 2046;
        ELSIF x = 8328 THEN
            tanh_f := 2046;
        ELSIF x = 8329 THEN
            tanh_f := 2046;
        ELSIF x = 8330 THEN
            tanh_f := 2046;
        ELSIF x = 8331 THEN
            tanh_f := 2046;
        ELSIF x = 8332 THEN
            tanh_f := 2046;
        ELSIF x = 8333 THEN
            tanh_f := 2046;
        ELSIF x = 8334 THEN
            tanh_f := 2046;
        ELSIF x = 8335 THEN
            tanh_f := 2046;
        ELSIF x = 8336 THEN
            tanh_f := 2046;
        ELSIF x = 8337 THEN
            tanh_f := 2046;
        ELSIF x = 8338 THEN
            tanh_f := 2046;
        ELSIF x = 8339 THEN
            tanh_f := 2046;
        ELSIF x = 8340 THEN
            tanh_f := 2046;
        ELSIF x = 8341 THEN
            tanh_f := 2046;
        ELSIF x = 8342 THEN
            tanh_f := 2046;
        ELSIF x = 8343 THEN
            tanh_f := 2046;
        ELSIF x = 8344 THEN
            tanh_f := 2046;
        ELSIF x = 8345 THEN
            tanh_f := 2046;
        ELSIF x = 8346 THEN
            tanh_f := 2046;
        ELSIF x = 8347 THEN
            tanh_f := 2046;
        ELSIF x = 8348 THEN
            tanh_f := 2046;
        ELSIF x = 8349 THEN
            tanh_f := 2046;
        ELSIF x = 8350 THEN
            tanh_f := 2046;
        ELSIF x = 8351 THEN
            tanh_f := 2046;
        ELSIF x = 8352 THEN
            tanh_f := 2046;
        ELSIF x = 8353 THEN
            tanh_f := 2046;
        ELSIF x = 8354 THEN
            tanh_f := 2046;
        ELSIF x = 8355 THEN
            tanh_f := 2046;
        ELSIF x = 8356 THEN
            tanh_f := 2046;
        ELSIF x = 8357 THEN
            tanh_f := 2046;
        ELSIF x = 8358 THEN
            tanh_f := 2046;
        ELSIF x = 8359 THEN
            tanh_f := 2046;
        ELSIF x = 8360 THEN
            tanh_f := 2046;
        ELSIF x = 8361 THEN
            tanh_f := 2046;
        ELSIF x = 8362 THEN
            tanh_f := 2046;
        ELSIF x = 8363 THEN
            tanh_f := 2046;
        ELSIF x = 8364 THEN
            tanh_f := 2046;
        ELSIF x = 8365 THEN
            tanh_f := 2046;
        ELSIF x = 8366 THEN
            tanh_f := 2046;
        ELSIF x = 8367 THEN
            tanh_f := 2046;
        ELSIF x = 8368 THEN
            tanh_f := 2046;
        ELSIF x = 8369 THEN
            tanh_f := 2046;
        ELSIF x = 8370 THEN
            tanh_f := 2046;
        ELSIF x = 8371 THEN
            tanh_f := 2046;
        ELSIF x = 8372 THEN
            tanh_f := 2046;
        ELSIF x = 8373 THEN
            tanh_f := 2046;
        ELSIF x = 8374 THEN
            tanh_f := 2046;
        ELSIF x = 8375 THEN
            tanh_f := 2046;
        ELSIF x = 8376 THEN
            tanh_f := 2046;
        ELSIF x = 8377 THEN
            tanh_f := 2046;
        ELSIF x = 8378 THEN
            tanh_f := 2046;
        ELSIF x = 8379 THEN
            tanh_f := 2046;
        ELSIF x = 8380 THEN
            tanh_f := 2046;
        ELSIF x = 8381 THEN
            tanh_f := 2046;
        ELSIF x = 8382 THEN
            tanh_f := 2046;
        ELSIF x = 8383 THEN
            tanh_f := 2046;
        ELSIF x = 8384 THEN
            tanh_f := 2046;
        ELSIF x = 8385 THEN
            tanh_f := 2046;
        ELSIF x = 8386 THEN
            tanh_f := 2046;
        ELSIF x = 8387 THEN
            tanh_f := 2046;
        ELSIF x = 8388 THEN
            tanh_f := 2046;
        ELSIF x = 8389 THEN
            tanh_f := 2046;
        ELSIF x = 8390 THEN
            tanh_f := 2046;
        ELSIF x = 8391 THEN
            tanh_f := 2046;
        ELSIF x = 8392 THEN
            tanh_f := 2046;
        ELSIF x = 8393 THEN
            tanh_f := 2046;
        ELSIF x = 8394 THEN
            tanh_f := 2046;
        ELSIF x = 8395 THEN
            tanh_f := 2046;
        ELSIF x = 8396 THEN
            tanh_f := 2046;
        ELSIF x = 8397 THEN
            tanh_f := 2046;
        ELSIF x = 8398 THEN
            tanh_f := 2046;
        ELSIF x = 8399 THEN
            tanh_f := 2046;
        ELSIF x = 8400 THEN
            tanh_f := 2046;
        ELSIF x = 8401 THEN
            tanh_f := 2046;
        ELSIF x = 8402 THEN
            tanh_f := 2046;
        ELSIF x = 8403 THEN
            tanh_f := 2046;
        ELSIF x = 8404 THEN
            tanh_f := 2046;
        ELSIF x = 8405 THEN
            tanh_f := 2046;
        ELSIF x = 8406 THEN
            tanh_f := 2046;
        ELSIF x = 8407 THEN
            tanh_f := 2046;
        ELSIF x = 8408 THEN
            tanh_f := 2046;
        ELSIF x = 8409 THEN
            tanh_f := 2046;
        ELSIF x = 8410 THEN
            tanh_f := 2046;
        ELSIF x = 8411 THEN
            tanh_f := 2046;
        ELSIF x = 8412 THEN
            tanh_f := 2046;
        ELSIF x = 8413 THEN
            tanh_f := 2046;
        ELSIF x = 8414 THEN
            tanh_f := 2046;
        ELSIF x = 8415 THEN
            tanh_f := 2046;
        ELSIF x = 8416 THEN
            tanh_f := 2046;
        ELSIF x = 8417 THEN
            tanh_f := 2046;
        ELSIF x = 8418 THEN
            tanh_f := 2046;
        ELSIF x = 8419 THEN
            tanh_f := 2046;
        ELSIF x = 8420 THEN
            tanh_f := 2046;
        ELSIF x = 8421 THEN
            tanh_f := 2046;
        ELSIF x = 8422 THEN
            tanh_f := 2046;
        ELSIF x = 8423 THEN
            tanh_f := 2046;
        ELSIF x = 8424 THEN
            tanh_f := 2046;
        ELSIF x = 8425 THEN
            tanh_f := 2046;
        ELSIF x = 8426 THEN
            tanh_f := 2046;
        ELSIF x = 8427 THEN
            tanh_f := 2046;
        ELSIF x = 8428 THEN
            tanh_f := 2046;
        ELSIF x = 8429 THEN
            tanh_f := 2046;
        ELSIF x = 8430 THEN
            tanh_f := 2046;
        ELSIF x = 8431 THEN
            tanh_f := 2046;
        ELSIF x = 8432 THEN
            tanh_f := 2046;
        ELSIF x = 8433 THEN
            tanh_f := 2046;
        ELSIF x = 8434 THEN
            tanh_f := 2046;
        ELSIF x = 8435 THEN
            tanh_f := 2046;
        ELSIF x = 8436 THEN
            tanh_f := 2046;
        ELSIF x = 8437 THEN
            tanh_f := 2046;
        ELSIF x = 8438 THEN
            tanh_f := 2046;
        ELSIF x = 8439 THEN
            tanh_f := 2046;
        ELSIF x = 8440 THEN
            tanh_f := 2046;
        ELSIF x = 8441 THEN
            tanh_f := 2046;
        ELSIF x = 8442 THEN
            tanh_f := 2046;
        ELSIF x = 8443 THEN
            tanh_f := 2046;
        ELSIF x = 8444 THEN
            tanh_f := 2046;
        ELSIF x = 8445 THEN
            tanh_f := 2046;
        ELSIF x = 8446 THEN
            tanh_f := 2046;
        ELSIF x = 8447 THEN
            tanh_f := 2046;
        ELSIF x >= 8448 THEN
            tanh_f := 2048;
        END IF;
        RETURN tanh_f;
    END;
END PACKAGE BODY tanh_pkg;